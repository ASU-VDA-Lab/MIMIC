module fake_jpeg_18150_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_18),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_46),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_24),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_38),
.B1(n_44),
.B2(n_34),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_61),
.B1(n_40),
.B2(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_51),
.B(n_54),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_45),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_57),
.A2(n_63),
.B1(n_65),
.B2(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_30),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_25),
.B1(n_20),
.B2(n_23),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_20),
.B1(n_27),
.B2(n_24),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_32),
.B1(n_26),
.B2(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_70),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_59),
.B(n_55),
.C(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_72),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_39),
.B(n_43),
.C(n_40),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_43),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_75),
.B(n_33),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_86),
.B1(n_0),
.B2(n_1),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_0),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_73),
.B1(n_83),
.B2(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_32),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_26),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_96),
.B1(n_78),
.B2(n_70),
.Y(n_124)
);

NOR2xp67_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_88),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_68),
.B1(n_49),
.B2(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_105),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_56),
.B(n_48),
.C(n_62),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_103),
.B1(n_109),
.B2(n_79),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_62),
.B1(n_67),
.B2(n_22),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_120),
.C(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_90),
.B1(n_89),
.B2(n_80),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_115),
.B1(n_124),
.B2(n_125),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_75),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_123),
.Y(n_127)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_74),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_122),
.A2(n_104),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_75),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_87),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_100),
.B(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_102),
.C(n_91),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_102),
.C(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_91),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_124),
.B1(n_120),
.B2(n_111),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_147),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_113),
.B1(n_112),
.B2(n_106),
.Y(n_142)
);

OAI321xp33_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_111),
.A3(n_123),
.B1(n_110),
.B2(n_119),
.C(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_99),
.Y(n_146)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_12),
.B1(n_10),
.B2(n_14),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_129),
.C(n_133),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_150),
.B(n_153),
.Y(n_156)
);

AOI222xp33_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_127),
.B1(n_137),
.B2(n_135),
.C1(n_138),
.C2(n_136),
.Y(n_151)
);

AOI31xp67_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_145),
.A3(n_147),
.B(n_4),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_128),
.C(n_2),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_148),
.Y(n_158)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_159),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_158),
.B(n_1),
.Y(n_164)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_141),
.B1(n_144),
.B2(n_139),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_151),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_1),
.B(n_3),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_164),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_4),
.B(n_5),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_158),
.C(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_166),
.B(n_168),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_165),
.B(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_4),
.C(n_5),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_170),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_7),
.Y(n_173)
);


endmodule