module fake_jpeg_19996_n_285 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_285);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_3),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_18),
.B1(n_29),
.B2(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_33),
.B1(n_36),
.B2(n_26),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_62),
.Y(n_68)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_18),
.B1(n_29),
.B2(n_24),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_24),
.B1(n_36),
.B2(n_23),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_26),
.B(n_23),
.C(n_36),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_69),
.B1(n_78),
.B2(n_80),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_67),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_24),
.B1(n_33),
.B2(n_21),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_74),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_76),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_79),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_30),
.B1(n_19),
.B2(n_21),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_81),
.B(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_34),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_85),
.A2(n_102),
.B1(n_25),
.B2(n_28),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_90),
.Y(n_122)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_17),
.B1(n_22),
.B2(n_19),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_53),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_54),
.B(n_17),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_33),
.B1(n_41),
.B2(n_37),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_95),
.B1(n_103),
.B2(n_25),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_43),
.B1(n_41),
.B2(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_20),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_20),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_32),
.B1(n_22),
.B2(n_30),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_25),
.B1(n_28),
.B2(n_4),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_49),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_20),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_31),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_32),
.B1(n_26),
.B2(n_23),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_56),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_66),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_86),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_70),
.A2(n_25),
.B(n_1),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_127),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_87),
.B1(n_96),
.B2(n_100),
.Y(n_146)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_125),
.B1(n_128),
.B2(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_68),
.A2(n_31),
.B1(n_28),
.B2(n_4),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_68),
.A2(n_97),
.B1(n_65),
.B2(n_98),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_80),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_130),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_88),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_103),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_126),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_101),
.C(n_95),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_95),
.C(n_94),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_91),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_154),
.B1(n_115),
.B2(n_113),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_147),
.A2(n_152),
.B(n_104),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_78),
.B1(n_95),
.B2(n_94),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_151),
.B1(n_145),
.B2(n_143),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_149),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_94),
.B1(n_84),
.B2(n_89),
.Y(n_151)
);

HAxp5_ASAP7_75t_SL g152 ( 
.A(n_114),
.B(n_28),
.CON(n_152),
.SN(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_84),
.B1(n_75),
.B2(n_72),
.Y(n_154)
);

OR2x4_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_129),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_128),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_111),
.B(n_16),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_156),
.B(n_157),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_106),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_158),
.B(n_112),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_167),
.B(n_179),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_171),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_170),
.B1(n_134),
.B2(n_144),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_107),
.B1(n_124),
.B2(n_122),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_172),
.B(n_176),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_107),
.B1(n_115),
.B2(n_108),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_175),
.A2(n_155),
.B1(n_147),
.B2(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_108),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_120),
.B(n_109),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_140),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_183),
.B(n_0),
.Y(n_193)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_120),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_152),
.A2(n_71),
.B(n_3),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_142),
.C(n_143),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_196),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_200),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_192),
.B1(n_204),
.B2(n_174),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_134),
.B1(n_150),
.B2(n_71),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_201),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_166),
.B(n_3),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_150),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_197),
.B(n_185),
.Y(n_217)
);

AO21x2_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_6),
.B(n_7),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_182),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_209),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_15),
.B1(n_16),
.B2(n_10),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_175),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_160),
.B1(n_163),
.B2(n_172),
.Y(n_216)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_218),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_216),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_226),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_179),
.B(n_186),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_201),
.B(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_222),
.B(n_159),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_228),
.B1(n_173),
.B2(n_165),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_225),
.B(n_227),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_177),
.B(n_162),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_163),
.C(n_176),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_191),
.A2(n_162),
.B(n_169),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_201),
.B1(n_207),
.B2(n_188),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_235),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_197),
.C(n_205),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_233),
.C(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_205),
.C(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_203),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_221),
.A2(n_201),
.B(n_203),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_236),
.B(n_244),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_201),
.CI(n_180),
.CON(n_237),
.SN(n_237)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_180),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_237),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_224),
.B1(n_210),
.B2(n_215),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_211),
.B(n_165),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_252),
.C(n_253),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_235),
.C(n_231),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_223),
.C(n_212),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_226),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_241),
.C(n_238),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_237),
.Y(n_260)
);

INVxp33_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_253),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_264),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_258),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_238),
.C(n_240),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_240),
.B(n_255),
.Y(n_266)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_269),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_251),
.B(n_232),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_270),
.B(n_271),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_246),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_239),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_242),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_276),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_246),
.C(n_8),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_269),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_277),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_7),
.C(n_12),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_278),
.A2(n_273),
.B(n_275),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_279),
.C(n_277),
.Y(n_282)
);

AOI211xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_280),
.B(n_13),
.C(n_14),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_12),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_13),
.Y(n_285)
);


endmodule