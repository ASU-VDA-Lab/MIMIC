module fake_jpeg_878_n_256 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_23),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_44),
.B(n_49),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_1),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_18),
.B(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_2),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_3),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_67),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_68),
.B(n_103),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_19),
.B1(n_37),
.B2(n_31),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_73),
.A2(n_33),
.B1(n_5),
.B2(n_6),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_75),
.B(n_33),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_30),
.Y(n_80)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_31),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_20),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_19),
.B1(n_39),
.B2(n_35),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_26),
.C(n_37),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_35),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_4),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_40),
.A2(n_32),
.B1(n_28),
.B2(n_27),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_102),
.B1(n_101),
.B2(n_96),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_45),
.A2(n_32),
.B1(n_28),
.B2(n_27),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_26),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_61),
.B1(n_58),
.B2(n_42),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_41),
.B(n_37),
.Y(n_103)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_107),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_110),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_109),
.B(n_127),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_84),
.C(n_89),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_116),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_112),
.Y(n_138)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_3),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_86),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_17),
.C(n_63),
.Y(n_116)
);

AO22x2_ASAP7_75t_L g117 ( 
.A1(n_75),
.A2(n_33),
.B1(n_5),
.B2(n_6),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_131),
.B(n_74),
.C(n_94),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_125),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_4),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_126),
.Y(n_150)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_14),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_70),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_135),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_70),
.A2(n_10),
.B1(n_13),
.B2(n_104),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_10),
.B(n_13),
.C(n_97),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_86),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_93),
.B1(n_73),
.B2(n_92),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_136),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_71),
.B(n_78),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_142),
.B(n_114),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_90),
.B1(n_94),
.B2(n_96),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_90),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_86),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_159),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_109),
.B1(n_117),
.B2(n_131),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_85),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_158),
.C(n_116),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_101),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_115),
.B(n_74),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_74),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_114),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_108),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_161),
.B(n_162),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_179),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_171),
.B(n_175),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_SL g194 ( 
.A1(n_172),
.A2(n_184),
.B(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_148),
.B(n_117),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_152),
.B(n_130),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_181),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_114),
.C(n_107),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_186),
.C(n_167),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_150),
.B(n_113),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_123),
.C(n_134),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_162),
.B(n_161),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_192),
.B(n_195),
.Y(n_215)
);

AO22x1_ASAP7_75t_SL g189 ( 
.A1(n_164),
.A2(n_154),
.B1(n_163),
.B2(n_152),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_200),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_165),
.A2(n_152),
.B(n_163),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_203),
.B1(n_170),
.B2(n_168),
.Y(n_218)
);

A2O1A1O1Ixp25_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_147),
.B(n_154),
.C(n_142),
.D(n_158),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_196),
.B(n_145),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_180),
.A2(n_157),
.B(n_140),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_155),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_202),
.A2(n_181),
.B1(n_168),
.B2(n_178),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_164),
.B1(n_174),
.B2(n_177),
.Y(n_203)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_186),
.B(n_150),
.CI(n_157),
.CON(n_205),
.SN(n_205)
);

NOR2x1_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_169),
.Y(n_217)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_166),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_209),
.B(n_219),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

AOI221xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_182),
.B1(n_173),
.B2(n_175),
.C(n_171),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_214),
.C(n_217),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_212),
.A2(n_204),
.B1(n_189),
.B2(n_200),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_197),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_218),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_191),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_196),
.C(n_190),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_210),
.B1(n_214),
.B2(n_208),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_207),
.C(n_217),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_190),
.C(n_192),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_225),
.C(n_215),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_203),
.C(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_231),
.B(n_232),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_237),
.B1(n_238),
.B2(n_188),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_224),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_216),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_219),
.B1(n_218),
.B2(n_206),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_206),
.C(n_208),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_227),
.B(n_221),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_236),
.A2(n_228),
.B1(n_230),
.B2(n_205),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_205),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_223),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_247),
.B(n_248),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_212),
.Y(n_247)
);

OAI221xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_195),
.B1(n_189),
.B2(n_199),
.C(n_204),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_249),
.A2(n_138),
.B1(n_131),
.B2(n_112),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_245),
.A2(n_240),
.B(n_244),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_251),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_252),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_245),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_253),
.Y(n_256)
);


endmodule