module fake_jpeg_30095_n_545 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_545);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_545;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx3_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_17),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_53),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_8),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_58),
.Y(n_106)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_8),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_74),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_66),
.Y(n_136)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_70),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_30),
.B(n_8),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_100),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_85),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_22),
.B(n_7),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_86),
.B(n_88),
.Y(n_143)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_30),
.B(n_7),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_31),
.B(n_9),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_94),
.B(n_45),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_46),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_35),
.B1(n_31),
.B2(n_41),
.Y(n_111)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

BUFx4f_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_29),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_20),
.Y(n_122)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_44),
.B1(n_41),
.B2(n_35),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_105),
.A2(n_112),
.B1(n_113),
.B2(n_121),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_111),
.A2(n_141),
.B1(n_25),
.B2(n_1),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_71),
.B1(n_50),
.B2(n_49),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_50),
.B1(n_20),
.B2(n_28),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_91),
.A2(n_50),
.B1(n_20),
.B2(n_28),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_98),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_58),
.B(n_44),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_124),
.B(n_134),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_74),
.B(n_48),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_48),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_146),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_45),
.B1(n_43),
.B2(n_38),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_73),
.A2(n_28),
.B1(n_27),
.B2(n_38),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_145),
.A2(n_151),
.B1(n_164),
.B2(n_121),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_76),
.A2(n_28),
.B1(n_27),
.B2(n_43),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_84),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_62),
.Y(n_163)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_63),
.A2(n_28),
.B1(n_27),
.B2(n_23),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_100),
.B(n_23),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_60),
.Y(n_172)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_125),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_171),
.B(n_173),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_190),
.Y(n_228)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_175),
.Y(n_254)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_176),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_109),
.A2(n_143),
.B(n_106),
.Y(n_177)
);

OR2x2_ASAP7_75t_SL g235 ( 
.A(n_177),
.B(n_185),
.Y(n_235)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_179),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_55),
.B(n_29),
.C(n_25),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_180),
.B(n_187),
.Y(n_278)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_107),
.B(n_25),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_182),
.Y(n_242)
);

XNOR2x1_ASAP7_75t_SL g182 ( 
.A(n_155),
.B(n_79),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_117),
.A2(n_25),
.B(n_29),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_183),
.Y(n_267)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_135),
.A2(n_25),
.B(n_27),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_129),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_25),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_189),
.B(n_193),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_129),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_114),
.A2(n_80),
.B1(n_77),
.B2(n_75),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_192),
.A2(n_207),
.B1(n_211),
.B2(n_223),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_123),
.B(n_52),
.C(n_72),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_194),
.B(n_213),
.C(n_219),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_137),
.B(n_27),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_196),
.B(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_197),
.Y(n_279)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g259 ( 
.A1(n_199),
.A2(n_11),
.B1(n_13),
.B2(n_16),
.Y(n_259)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_142),
.Y(n_200)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_139),
.Y(n_201)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_116),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_202),
.B(n_216),
.Y(n_257)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_204),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_129),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_208),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_126),
.A2(n_70),
.B1(n_1),
.B2(n_2),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_112),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_115),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_218),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_145),
.A2(n_151),
.B1(n_113),
.B2(n_164),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_114),
.Y(n_212)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_212),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_131),
.B(n_10),
.C(n_3),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_126),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_214),
.A2(n_225),
.B1(n_160),
.B2(n_128),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_120),
.Y(n_215)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_215),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_148),
.B(n_127),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_217),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_152),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_153),
.A2(n_18),
.B1(n_5),
.B2(n_6),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_219),
.A2(n_224),
.B1(n_213),
.B2(n_167),
.Y(n_260)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_148),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_227),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_127),
.A2(n_18),
.B(n_5),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_221),
.B(n_9),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_222),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_153),
.A2(n_161),
.B1(n_120),
.B2(n_156),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_136),
.A2(n_12),
.B(n_6),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_133),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_230),
.B(n_259),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_186),
.A2(n_161),
.B1(n_156),
.B2(n_147),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_241),
.A2(n_248),
.B1(n_202),
.B2(n_171),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_244),
.A2(n_250),
.B(n_243),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_199),
.A2(n_147),
.B1(n_162),
.B2(n_110),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_130),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_249),
.B(n_253),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_182),
.A2(n_144),
.B1(n_136),
.B2(n_12),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_169),
.B(n_144),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_260),
.A2(n_270),
.B1(n_277),
.B2(n_265),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_177),
.B(n_13),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_271),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_188),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_175),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_194),
.A2(n_0),
.B1(n_13),
.B2(n_16),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_183),
.B(n_16),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_180),
.B(n_18),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_273),
.B(n_262),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_189),
.B(n_0),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_189),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_242),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_181),
.A2(n_198),
.B1(n_191),
.B2(n_178),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_280),
.A2(n_295),
.B1(n_298),
.B2(n_304),
.Y(n_338)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_283),
.B(n_288),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_261),
.B1(n_260),
.B2(n_267),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_284),
.A2(n_305),
.B1(n_310),
.B2(n_239),
.Y(n_335)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_251),
.Y(n_285)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_258),
.B(n_173),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_286),
.B(n_289),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_235),
.B(n_173),
.C(n_184),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_297),
.C(n_300),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_242),
.B(n_216),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_288),
.B(n_283),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_176),
.Y(n_289)
);

INVx5_ASAP7_75t_SL g290 ( 
.A(n_243),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_290),
.B(n_296),
.Y(n_352)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_232),
.Y(n_294)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_261),
.A2(n_185),
.B1(n_192),
.B2(n_170),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_228),
.B(n_217),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_235),
.A2(n_201),
.B1(n_174),
.B2(n_168),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_242),
.B(n_216),
.C(n_179),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_229),
.B(n_279),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_301),
.B(n_309),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_227),
.C(n_203),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_302),
.B(n_316),
.C(n_297),
.Y(n_364)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_265),
.A2(n_222),
.B1(n_221),
.B2(n_212),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_273),
.A2(n_226),
.B1(n_223),
.B2(n_195),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_271),
.A2(n_264),
.B(n_255),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_306),
.A2(n_319),
.B(n_282),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_274),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_307),
.B(n_308),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_255),
.B(n_230),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_259),
.A2(n_270),
.B1(n_240),
.B2(n_237),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_311),
.A2(n_313),
.B1(n_314),
.B2(n_317),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_231),
.B(n_252),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_312),
.B(n_319),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_259),
.A2(n_230),
.B1(n_237),
.B2(n_257),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_259),
.A2(n_240),
.B1(n_237),
.B2(n_257),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_257),
.B(n_232),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_324),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_252),
.B(n_234),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_266),
.A2(n_272),
.B1(n_233),
.B2(n_269),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_234),
.Y(n_318)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_254),
.B(n_268),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_239),
.Y(n_340)
);

AO21x2_ASAP7_75t_L g322 ( 
.A1(n_233),
.A2(n_262),
.B(n_272),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_323),
.B(n_317),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_266),
.A2(n_254),
.B(n_268),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_263),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_325),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_256),
.B(n_245),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_326),
.B(n_327),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_245),
.B(n_275),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_292),
.B(n_263),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_329),
.B(n_334),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_310),
.A2(n_233),
.B1(n_236),
.B2(n_275),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_330),
.A2(n_335),
.B1(n_355),
.B2(n_356),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_308),
.A2(n_236),
.B(n_246),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g401 ( 
.A1(n_331),
.A2(n_350),
.B(n_362),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_238),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_332),
.A2(n_333),
.B(n_345),
.Y(n_389)
);

AOI21xp33_ASAP7_75t_L g334 ( 
.A1(n_282),
.A2(n_246),
.B(n_238),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_336),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_340),
.B(n_342),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_239),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_336),
.C(n_331),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_326),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_293),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_327),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_354),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_289),
.A2(n_293),
.B1(n_286),
.B2(n_311),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_293),
.A2(n_295),
.B1(n_306),
.B2(n_302),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_357),
.B(n_361),
.Y(n_390)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_294),
.Y(n_358)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_358),
.Y(n_384)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_360),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_300),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_341),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_307),
.B(n_298),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_366),
.Y(n_375)
);

AOI32xp33_ASAP7_75t_L g368 ( 
.A1(n_325),
.A2(n_287),
.A3(n_322),
.B1(n_290),
.B2(n_315),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_368),
.A2(n_360),
.B(n_369),
.Y(n_404)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_285),
.Y(n_369)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_369),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_347),
.A2(n_280),
.B1(n_322),
.B2(n_324),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_370),
.A2(n_378),
.B(n_404),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_316),
.Y(n_371)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_371),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_363),
.B(n_323),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_374),
.B(n_386),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_359),
.A2(n_322),
.B1(n_324),
.B2(n_303),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_376),
.A2(n_379),
.B1(n_381),
.B2(n_387),
.Y(n_405)
);

AOI22x1_ASAP7_75t_SL g377 ( 
.A1(n_368),
.A2(n_322),
.B1(n_290),
.B2(n_299),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_377),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_332),
.A2(n_322),
.B1(n_318),
.B2(n_320),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_359),
.A2(n_299),
.B1(n_333),
.B2(n_338),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_338),
.A2(n_299),
.B1(n_351),
.B2(n_342),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_335),
.A2(n_330),
.B1(n_356),
.B2(n_355),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_382),
.A2(n_396),
.B1(n_371),
.B2(n_370),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_383),
.B(n_387),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_367),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_385),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_363),
.B(n_351),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_353),
.A2(n_365),
.B1(n_367),
.B2(n_364),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_332),
.A2(n_345),
.B1(n_365),
.B2(n_353),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_392),
.A2(n_395),
.B1(n_399),
.B2(n_349),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_394),
.C(n_383),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_345),
.A2(n_350),
.B1(n_344),
.B2(n_357),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_344),
.A2(n_352),
.B1(n_329),
.B2(n_337),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_397),
.Y(n_417)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_346),
.Y(n_398)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_398),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_352),
.A2(n_362),
.B1(n_339),
.B2(n_328),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_401),
.A2(n_372),
.B(n_374),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_358),
.B(n_328),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_402),
.B(n_391),
.Y(n_427)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_339),
.Y(n_403)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_377),
.A2(n_348),
.B1(n_349),
.B2(n_343),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_406),
.A2(n_412),
.B1(n_414),
.B2(n_428),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_375),
.B(n_348),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_407),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_402),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_409),
.B(n_425),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_410),
.A2(n_423),
.B1(n_389),
.B2(n_397),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_377),
.A2(n_343),
.B1(n_380),
.B2(n_382),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_380),
.A2(n_373),
.B1(n_385),
.B2(n_378),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_386),
.B(n_373),
.Y(n_416)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_416),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_419),
.B(n_420),
.Y(n_445)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_400),
.Y(n_422)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_379),
.A2(n_376),
.B1(n_381),
.B2(n_392),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_400),
.Y(n_424)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_424),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_396),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_394),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_433),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_435),
.Y(n_439)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_431),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_388),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_432),
.B(n_421),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_393),
.B(n_395),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_434),
.B(n_390),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_399),
.B(n_371),
.Y(n_435)
);

HAxp5_ASAP7_75t_SL g436 ( 
.A(n_416),
.B(n_401),
.CON(n_436),
.SN(n_436)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_436),
.A2(n_440),
.B(n_420),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_437),
.B(n_405),
.Y(n_475)
);

INVx2_ASAP7_75t_R g438 ( 
.A(n_411),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_438),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_429),
.A2(n_372),
.B(n_404),
.Y(n_440)
);

INVx8_ASAP7_75t_L g442 ( 
.A(n_422),
.Y(n_442)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_442),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_417),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_443),
.B(n_459),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_412),
.A2(n_389),
.B1(n_388),
.B2(n_391),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_448),
.A2(n_455),
.B1(n_461),
.B2(n_415),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_408),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_456),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_390),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_433),
.C(n_434),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_453),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_406),
.A2(n_398),
.B1(n_403),
.B2(n_414),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_424),
.B(n_408),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_411),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_458),
.B(n_418),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_428),
.A2(n_415),
.B1(n_429),
.B2(n_413),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_413),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_464),
.B(n_476),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_484),
.Y(n_491)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_469),
.A2(n_453),
.B1(n_441),
.B2(n_436),
.Y(n_492)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_438),
.Y(n_471)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_471),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_438),
.Y(n_472)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_472),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_419),
.C(n_410),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_445),
.C(n_437),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_475),
.B(n_448),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_405),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_454),
.B(n_432),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_477),
.A2(n_449),
.B1(n_452),
.B2(n_439),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_444),
.A2(n_423),
.B1(n_418),
.B2(n_421),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_478),
.A2(n_441),
.B1(n_444),
.B2(n_442),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_458),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_480),
.Y(n_485)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_447),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_447),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_481),
.B(n_482),
.Y(n_500)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_452),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_439),
.B(n_431),
.Y(n_484)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_488),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_490),
.B(n_496),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_492),
.A2(n_499),
.B1(n_474),
.B2(n_484),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_465),
.B(n_445),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_463),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_451),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_461),
.C(n_440),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_497),
.B(n_491),
.C(n_501),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_455),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_498),
.B(n_479),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_501),
.B(n_495),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_504),
.B(n_508),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_475),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_505),
.B(n_509),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_506),
.B(n_507),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_494),
.A2(n_471),
.B(n_463),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_485),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_510),
.B(n_493),
.Y(n_520)
);

AOI21xp33_ASAP7_75t_L g511 ( 
.A1(n_487),
.A2(n_467),
.B(n_477),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_511),
.A2(n_500),
.B(n_489),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_496),
.B(n_469),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_497),
.C(n_495),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_486),
.B(n_474),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_514),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_492),
.A2(n_470),
.B1(n_482),
.B2(n_481),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_478),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_516),
.A2(n_519),
.B(n_507),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_517),
.B(n_520),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_506),
.A2(n_490),
.B(n_468),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_505),
.B(n_466),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_522),
.A2(n_468),
.B1(n_480),
.B2(n_510),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_525),
.B(n_515),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_526),
.B(n_527),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_518),
.A2(n_503),
.B(n_508),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_528),
.B(n_522),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_529),
.B(n_530),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_483),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_533),
.B(n_534),
.Y(n_536)
);

AOI21xp33_ASAP7_75t_L g534 ( 
.A1(n_531),
.A2(n_523),
.B(n_483),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_457),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_537),
.A2(n_460),
.B(n_457),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_536),
.A2(n_535),
.B(n_517),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_538),
.A2(n_539),
.B(n_443),
.Y(n_540)
);

AOI21x1_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_509),
.B(n_460),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_417),
.C(n_430),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_524),
.B(n_512),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_524),
.Y(n_544)
);

FAx1_ASAP7_75t_SL g545 ( 
.A(n_544),
.B(n_502),
.CI(n_531),
.CON(n_545),
.SN(n_545)
);


endmodule