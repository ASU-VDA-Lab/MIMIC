module fake_jpeg_14060_n_100 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_17),
.B1(n_12),
.B2(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_11),
.B(n_5),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_28),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_22),
.Y(n_49)
);

CKINVDCx6p67_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_48),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_28),
.C(n_26),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_46),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_28),
.C(n_24),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_39),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_19),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_15),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_59),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_41),
.B(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_20),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_13),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_45),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_70),
.B(n_33),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_61),
.B1(n_49),
.B2(n_46),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_63),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_43),
.B1(n_51),
.B2(n_52),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_52),
.B1(n_23),
.B2(n_47),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_54),
.B1(n_31),
.B2(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_5),
.Y(n_73)
);

AOI221xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_70),
.B1(n_39),
.B2(n_23),
.C(n_33),
.Y(n_77)
);

AOI221xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_74),
.B1(n_60),
.B2(n_67),
.C(n_69),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_77),
.B(n_79),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_58),
.B(n_63),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_56),
.C(n_41),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_56),
.B1(n_25),
.B2(n_31),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_18),
.B(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_89),
.B(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_8),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_93),
.A2(n_6),
.B(n_8),
.C(n_18),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_91),
.A2(n_90),
.B(n_7),
.Y(n_94)
);

OAI21x1_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_95),
.B(n_96),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_17),
.C(n_16),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_23),
.B(n_17),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_16),
.Y(n_100)
);


endmodule