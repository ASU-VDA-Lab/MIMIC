module real_jpeg_20177_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_324, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_324;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_0),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_69),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_0),
.A2(n_60),
.B1(n_61),
.B2(n_69),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_69),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_1),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_1),
.A2(n_60),
.B1(n_61),
.B2(n_114),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_114),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_114),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_2),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_2),
.A2(n_30),
.B1(n_60),
.B2(n_61),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_2),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_3),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_82),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_82),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_82),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_4),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_39),
.B1(n_60),
.B2(n_61),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_5),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_280)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_7),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_108),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_7),
.A2(n_60),
.B1(n_61),
.B2(n_108),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_108),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_8),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_8),
.B(n_34),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_8),
.A2(n_57),
.B(n_60),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_117),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_8),
.A2(n_97),
.B1(n_98),
.B2(n_177),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_8),
.B(n_42),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g207 ( 
.A1(n_8),
.A2(n_36),
.B(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_9),
.Y(n_98)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_9),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_10),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_112),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_112),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_112),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_12),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_119),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_119),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_119),
.Y(n_177)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_14),
.A2(n_36),
.A3(n_45),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_22),
.B(n_72),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_52),
.B1(n_53),
.B2(n_71),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_27),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_32),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g116 ( 
.A(n_29),
.B(n_117),
.CON(n_116),
.SN(n_116)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_31),
.A2(n_34),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_31),
.A2(n_34),
.B1(n_81),
.B2(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_32),
.B(n_36),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_33),
.A2(n_35),
.B1(n_116),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_43),
.B(n_46),
.C(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_46),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_35),
.B(n_117),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_47),
.B(n_50),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_47),
.B1(n_50),
.B2(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_42),
.A2(n_47),
.B1(n_64),
.B2(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_42),
.A2(n_47),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_42),
.A2(n_47),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_43),
.A2(n_48),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_43),
.A2(n_48),
.B1(n_113),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_43),
.A2(n_48),
.B1(n_146),
.B2(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_43),
.A2(n_48),
.B1(n_127),
.B2(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_43),
.A2(n_48),
.B1(n_86),
.B2(n_292),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_45),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_44),
.B(n_46),
.Y(n_203)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_45),
.A2(n_58),
.B(n_117),
.C(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_63),
.C(n_65),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_63),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_54),
.A2(n_78),
.B1(n_84),
.B2(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_59),
.B(n_62),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_59),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_59),
.B1(n_102),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_55),
.A2(n_59),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_55),
.A2(n_59),
.B1(n_173),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_55),
.A2(n_59),
.B1(n_193),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_55),
.A2(n_59),
.B1(n_107),
.B2(n_211),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_55),
.A2(n_59),
.B1(n_103),
.B2(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_55),
.A2(n_59),
.B1(n_247),
.B2(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_55),
.A2(n_59),
.B1(n_62),
.B2(n_280),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

CKINVDCx9p33_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_59),
.B(n_117),
.Y(n_178)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_61),
.B(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_66),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_68),
.B1(n_70),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_67),
.A2(n_70),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_67),
.A2(n_70),
.B1(n_125),
.B2(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_67),
.A2(n_70),
.B1(n_254),
.B2(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_79),
.C(n_83),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_310),
.Y(n_314)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_79),
.C(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_79),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_79),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_83),
.B(n_314),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_84),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI321xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_303),
.A3(n_315),
.B1(n_321),
.B2(n_322),
.C(n_324),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_284),
.B(n_302),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_260),
.B(n_283),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_152),
.B(n_236),
.C(n_259),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_137),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_93),
.B(n_137),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_120),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_95),
.B(n_104),
.C(n_120),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_101),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_96),
.B(n_101),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_97),
.A2(n_99),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_97),
.A2(n_133),
.B1(n_136),
.B2(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_97),
.A2(n_134),
.B1(n_162),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_97),
.A2(n_98),
.B1(n_165),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_97),
.A2(n_134),
.B1(n_151),
.B2(n_195),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_97),
.A2(n_100),
.B1(n_136),
.B2(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_97),
.A2(n_134),
.B(n_245),
.Y(n_278)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_98),
.B(n_117),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_115),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_129),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_128),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_122),
.B(n_128),
.C(n_129),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_126),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_132),
.Y(n_141)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_142),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_138),
.B(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_149),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_144),
.B(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_148),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_235),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_230),
.B(n_234),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_216),
.B(n_229),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_197),
.B(n_215),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_185),
.B(n_196),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_174),
.B(n_184),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_166),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_166),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_170),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_179),
.B(n_183),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_187),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_199),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_205),
.B1(n_213),
.B2(n_214),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_200),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_202),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_217),
.B(n_218),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_226),
.C(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_225),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_237),
.B(n_238),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_258),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_239),
.Y(n_258)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_248),
.B2(n_249),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_249),
.C(n_258),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_252),
.C(n_257),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_257),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_255),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_262),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_282),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_275),
.B2(n_276),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_276),
.C(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_268),
.C(n_272),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_270),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_274),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_281),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_277),
.A2(n_278),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_279),
.Y(n_295)
);

AOI21xp33_ASAP7_75t_L g312 ( 
.A1(n_278),
.A2(n_295),
.B(n_298),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_279),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_286),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_300),
.B2(n_301),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_294),
.C(n_301),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B(n_293),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_305),
.C(n_311),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_293),
.A2(n_305),
.B1(n_306),
.B2(n_320),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_293),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_300),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_313),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_313),
.Y(n_322)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_307),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_311),
.A2(n_312),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);


endmodule