module fake_jpeg_28879_n_184 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_184);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_5),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_2),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_17),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_8),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_0),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_3),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_3),
.B(n_4),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_58),
.Y(n_86)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_4),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_76),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_66),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_64),
.C(n_73),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_67),
.B1(n_58),
.B2(n_66),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_67),
.B1(n_73),
.B2(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_53),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_61),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_56),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_104),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_60),
.B(n_63),
.C(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_108),
.B(n_9),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_84),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_71),
.C(n_77),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_85),
.B1(n_56),
.B2(n_59),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_114),
.B1(n_117),
.B2(n_25),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_6),
.Y(n_135)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_54),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_116),
.B(n_120),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_56),
.B1(n_75),
.B2(n_85),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_121),
.Y(n_123)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_77),
.Y(n_120)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_128),
.Y(n_155)
);

AOI22x1_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_97),
.B1(n_77),
.B2(n_71),
.Y(n_127)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_133),
.B1(n_41),
.B2(n_19),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_5),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_143),
.B(n_18),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_59),
.B(n_26),
.C(n_28),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_135),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_103),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_7),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_8),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_31),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_141),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_145)
);

CKINVDCx12_ASAP7_75t_R g144 ( 
.A(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_48),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_150),
.B1(n_131),
.B2(n_50),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_13),
.B(n_14),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_157),
.B(n_49),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_125),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_156),
.B1(n_160),
.B2(n_45),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_150)
);

AOI221xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_152),
.B1(n_158),
.B2(n_133),
.C(n_124),
.Y(n_163)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_20),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_24),
.B1(n_29),
.B2(n_32),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_33),
.B(n_34),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_36),
.B(n_44),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_52),
.B1(n_46),
.B2(n_47),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_164),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_166),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_138),
.B1(n_131),
.B2(n_142),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_167),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_126),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_150),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_126),
.C(n_142),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_169),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_177),
.B(n_176),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_176),
.B(n_148),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_179),
.A2(n_168),
.B(n_148),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_173),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_154),
.A3(n_171),
.B1(n_174),
.B2(n_161),
.C1(n_146),
.C2(n_147),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_165),
.C(n_159),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_149),
.Y(n_184)
);


endmodule