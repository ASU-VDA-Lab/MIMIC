module fake_jpeg_6333_n_40 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_40);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_40;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_32;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx6p67_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_13),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_6),
.B(n_2),
.Y(n_28)
);

NOR3xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_29),
.C(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_5),
.B1(n_14),
.B2(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_18),
.B1(n_19),
.B2(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_26),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_33),
.C(n_20),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_35),
.B(n_25),
.Y(n_40)
);


endmodule