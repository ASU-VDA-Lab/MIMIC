module fake_aes_812_n_1582 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1582);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1582;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_822;
wire n_706;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1533;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1563;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1557;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1435;
wire n_1179;
wire n_1539;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_799;
wire n_423;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1577;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_1425;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_386;
wire n_659;
wire n_432;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_1576;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_1570;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_351;
wire n_401;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_1275;
wire n_955;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_1531;
wire n_371;
wire n_1548;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g347 ( .A(n_298), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_64), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_320), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_31), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_275), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_80), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_206), .Y(n_353) );
CKINVDCx16_ASAP7_75t_R g354 ( .A(n_323), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_0), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_70), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_132), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_216), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_172), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_337), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_133), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_54), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_283), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_292), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_1), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_8), .Y(n_366) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_144), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_77), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_46), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_91), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_72), .Y(n_371) );
BUFx2_ASAP7_75t_SL g372 ( .A(n_231), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_0), .Y(n_373) );
CKINVDCx16_ASAP7_75t_R g374 ( .A(n_197), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_300), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_280), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_73), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_173), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_88), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_170), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_249), .Y(n_381) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_35), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_72), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_154), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_279), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_171), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_281), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_14), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_316), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_126), .Y(n_390) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_252), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_256), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_335), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_165), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_204), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_45), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_14), .Y(n_397) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_339), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_274), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_47), .Y(n_400) );
INVxp67_ASAP7_75t_SL g401 ( .A(n_56), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_71), .Y(n_402) );
BUFx2_ASAP7_75t_L g403 ( .A(n_73), .Y(n_403) );
INVxp33_ASAP7_75t_L g404 ( .A(n_53), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_248), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_345), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_40), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_130), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_291), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_321), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_134), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_82), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_38), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_267), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_213), .Y(n_415) );
NOR2xp67_ASAP7_75t_L g416 ( .A(n_302), .B(n_217), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_129), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_293), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_89), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_166), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_294), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_228), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_297), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_43), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_24), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_247), .Y(n_426) );
CKINVDCx16_ASAP7_75t_R g427 ( .A(n_329), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_104), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_303), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_315), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_226), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_295), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_306), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_342), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_54), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_187), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_30), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_200), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_121), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_142), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_289), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_108), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_331), .Y(n_443) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_70), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_177), .B(n_64), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_15), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_29), .Y(n_447) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_181), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_34), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_307), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_287), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_112), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_153), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_199), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_227), .Y(n_455) );
INVxp33_ASAP7_75t_L g456 ( .A(n_138), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_179), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_101), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_273), .Y(n_459) );
INVxp33_ASAP7_75t_SL g460 ( .A(n_41), .Y(n_460) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_84), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_251), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_93), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_325), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_86), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_254), .Y(n_466) );
INVxp67_ASAP7_75t_SL g467 ( .A(n_4), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_241), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_93), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_240), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_145), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_109), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_67), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_301), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_86), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_74), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_313), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_147), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_229), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_195), .Y(n_480) );
INVxp67_ASAP7_75t_SL g481 ( .A(n_218), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_186), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_115), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_221), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_158), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_6), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_131), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_30), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_90), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_150), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_45), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_97), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_31), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_122), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_272), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_76), .Y(n_496) );
INVxp33_ASAP7_75t_SL g497 ( .A(n_243), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_258), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_103), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_66), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_222), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_76), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_224), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_232), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_96), .Y(n_505) );
BUFx3_ASAP7_75t_L g506 ( .A(n_189), .Y(n_506) );
CKINVDCx14_ASAP7_75t_R g507 ( .A(n_46), .Y(n_507) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_47), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_12), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_263), .Y(n_510) );
CKINVDCx14_ASAP7_75t_R g511 ( .A(n_136), .Y(n_511) );
BUFx3_ASAP7_75t_L g512 ( .A(n_152), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_209), .Y(n_513) );
INVxp67_ASAP7_75t_SL g514 ( .A(n_161), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_290), .Y(n_515) );
INVxp33_ASAP7_75t_SL g516 ( .A(n_29), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_262), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_123), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_97), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_105), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_149), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_43), .B(n_244), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_349), .B(n_1), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_359), .B(n_2), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_457), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_488), .Y(n_526) );
INVx4_ASAP7_75t_L g527 ( .A(n_380), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_457), .Y(n_528) );
INVx3_ASAP7_75t_L g529 ( .A(n_371), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_488), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_371), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_404), .B(n_2), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_377), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_377), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_347), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_353), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_354), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_457), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_457), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_360), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_408), .B(n_455), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_380), .B(n_3), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_476), .Y(n_543) );
NOR2x1_ASAP7_75t_L g544 ( .A(n_361), .B(n_3), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_468), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_404), .B(n_4), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_507), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_468), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_484), .B(n_5), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_364), .Y(n_550) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_468), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_433), .B(n_7), .Y(n_552) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_468), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_374), .Y(n_554) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_433), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_507), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_510), .B(n_8), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_375), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_363), .Y(n_559) );
BUFx3_ASAP7_75t_L g560 ( .A(n_436), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_376), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_458), .B(n_9), .Y(n_562) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_436), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_528), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_543), .B(n_496), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_559), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_556), .B(n_403), .Y(n_567) );
OR2x6_ASAP7_75t_SL g568 ( .A(n_537), .B(n_350), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_542), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_528), .Y(n_570) );
INVx4_ASAP7_75t_L g571 ( .A(n_542), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_556), .B(n_509), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_528), .Y(n_573) );
INVx5_ASAP7_75t_L g574 ( .A(n_555), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_559), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_542), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_541), .B(n_456), .Y(n_577) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_528), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_559), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_529), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_535), .B(n_456), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_554), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_535), .B(n_394), .Y(n_583) );
AND2x6_ASAP7_75t_L g584 ( .A(n_542), .B(n_451), .Y(n_584) );
AO21x2_ASAP7_75t_L g585 ( .A1(n_532), .A2(n_381), .B(n_378), .Y(n_585) );
INVx3_ASAP7_75t_L g586 ( .A(n_552), .Y(n_586) );
OR2x6_ASAP7_75t_L g587 ( .A(n_547), .B(n_372), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_529), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_529), .Y(n_589) );
NOR2xp33_ASAP7_75t_SL g590 ( .A(n_552), .B(n_427), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g591 ( .A(n_552), .B(n_445), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_528), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_532), .B(n_546), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_552), .B(n_348), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_536), .B(n_414), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_536), .B(n_511), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_540), .B(n_350), .Y(n_597) );
AND2x6_ASAP7_75t_L g598 ( .A(n_544), .B(n_451), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_540), .B(n_365), .Y(n_599) );
INVx5_ASAP7_75t_L g600 ( .A(n_555), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_546), .A2(n_352), .B1(n_362), .B2(n_356), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_529), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_524), .Y(n_603) );
INVx3_ASAP7_75t_L g604 ( .A(n_527), .Y(n_604) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_528), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_524), .B(n_365), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_550), .B(n_366), .Y(n_607) );
AO21x2_ASAP7_75t_L g608 ( .A1(n_549), .A2(n_385), .B(n_384), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_525), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_549), .B(n_369), .Y(n_610) );
INVx4_ASAP7_75t_L g611 ( .A(n_527), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_587), .A2(n_430), .B1(n_472), .B2(n_426), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_593), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_584), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_593), .B(n_550), .Y(n_615) );
BUFx4f_ASAP7_75t_L g616 ( .A(n_591), .Y(n_616) );
AND3x2_ASAP7_75t_SL g617 ( .A(n_568), .B(n_373), .C(n_368), .Y(n_617) );
NOR3xp33_ASAP7_75t_SL g618 ( .A(n_582), .B(n_547), .C(n_379), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_596), .B(n_562), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_596), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_580), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_565), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_581), .B(n_558), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_569), .A2(n_561), .B(n_558), .Y(n_624) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_584), .Y(n_625) );
INVx3_ASAP7_75t_L g626 ( .A(n_571), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_581), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_603), .B(n_561), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_577), .B(n_523), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_588), .Y(n_630) );
BUFx8_ASAP7_75t_L g631 ( .A(n_565), .Y(n_631) );
OAI22xp5_ASAP7_75t_SL g632 ( .A1(n_587), .A2(n_373), .B1(n_397), .B2(n_368), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_571), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_608), .B(n_527), .Y(n_634) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_584), .Y(n_635) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_571), .B(n_544), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_588), .Y(n_637) );
NAND3xp33_ASAP7_75t_SL g638 ( .A(n_590), .B(n_430), .C(n_426), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_566), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_610), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_566), .Y(n_641) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_584), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_575), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_610), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_607), .B(n_557), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_606), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_590), .A2(n_516), .B1(n_460), .B2(n_487), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_584), .A2(n_516), .B1(n_460), .B2(n_560), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_567), .B(n_497), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_575), .Y(n_650) );
AND2x6_ASAP7_75t_L g651 ( .A(n_569), .B(n_506), .Y(n_651) );
NOR2x1p5_ASAP7_75t_L g652 ( .A(n_567), .B(n_369), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_579), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_589), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_608), .B(n_560), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_572), .B(n_497), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_572), .A2(n_487), .B1(n_472), .B2(n_383), .Y(n_657) );
NAND2x1p5_ASAP7_75t_L g658 ( .A(n_571), .B(n_370), .Y(n_658) );
AO22x1_ASAP7_75t_L g659 ( .A1(n_584), .A2(n_383), .B1(n_400), .B2(n_379), .Y(n_659) );
NAND2x1p5_ASAP7_75t_L g660 ( .A(n_607), .B(n_396), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_585), .B(n_531), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_587), .A2(n_400), .B1(n_449), .B2(n_437), .Y(n_662) );
BUFx2_ASAP7_75t_L g663 ( .A(n_568), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_585), .B(n_531), .Y(n_664) );
INVx2_ASAP7_75t_SL g665 ( .A(n_591), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_579), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_589), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_585), .B(n_533), .Y(n_668) );
NOR2x1_ASAP7_75t_R g669 ( .A(n_594), .B(n_437), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_569), .B(n_533), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_594), .B(n_357), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_602), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_591), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_584), .Y(n_674) );
BUFx3_ASAP7_75t_L g675 ( .A(n_598), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_569), .B(n_534), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_597), .B(n_449), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_602), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_599), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_576), .B(n_534), .Y(n_680) );
INVx5_ASAP7_75t_L g681 ( .A(n_611), .Y(n_681) );
INVxp67_ASAP7_75t_L g682 ( .A(n_583), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_607), .B(n_526), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_607), .B(n_357), .Y(n_684) );
BUFx2_ASAP7_75t_L g685 ( .A(n_587), .Y(n_685) );
BUFx4f_ASAP7_75t_SL g686 ( .A(n_598), .Y(n_686) );
AO22x1_ASAP7_75t_L g687 ( .A1(n_598), .A2(n_500), .B1(n_463), .B2(n_358), .Y(n_687) );
AND2x4_ASAP7_75t_L g688 ( .A(n_594), .B(n_526), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_587), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_594), .B(n_417), .Y(n_690) );
BUFx2_ASAP7_75t_L g691 ( .A(n_598), .Y(n_691) );
INVxp67_ASAP7_75t_L g692 ( .A(n_595), .Y(n_692) );
AND2x4_ASAP7_75t_L g693 ( .A(n_576), .B(n_530), .Y(n_693) );
AND2x6_ASAP7_75t_SL g694 ( .A(n_601), .B(n_402), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_576), .Y(n_695) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_576), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_586), .A2(n_511), .B1(n_412), .B2(n_413), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_586), .B(n_358), .Y(n_698) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_586), .Y(n_699) );
INVxp67_ASAP7_75t_L g700 ( .A(n_598), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_586), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_598), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_604), .Y(n_703) );
BUFx2_ASAP7_75t_L g704 ( .A(n_611), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_631), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_613), .A2(n_397), .B1(n_425), .B2(n_424), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_696), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_660), .Y(n_708) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_644), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_615), .B(n_463), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_660), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_696), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_688), .Y(n_713) );
BUFx2_ASAP7_75t_SL g714 ( .A(n_665), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g715 ( .A1(n_624), .A2(n_604), .B(n_419), .C(n_435), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_624), .A2(n_604), .B(n_446), .C(n_465), .Y(n_716) );
INVx2_ASAP7_75t_SL g717 ( .A(n_616), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_634), .A2(n_611), .B(n_391), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_644), .A2(n_425), .B1(n_447), .B2(n_424), .Y(n_719) );
AND2x4_ASAP7_75t_L g720 ( .A(n_640), .B(n_382), .Y(n_720) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_614), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_646), .A2(n_627), .B1(n_689), .B2(n_685), .Y(n_722) );
AOI222xp33_ASAP7_75t_L g723 ( .A1(n_632), .A2(n_447), .B1(n_355), .B2(n_461), .C1(n_444), .C2(n_401), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_616), .B(n_405), .Y(n_724) );
CKINVDCx8_ASAP7_75t_R g725 ( .A(n_694), .Y(n_725) );
INVx3_ASAP7_75t_L g726 ( .A(n_626), .Y(n_726) );
BUFx2_ASAP7_75t_L g727 ( .A(n_631), .Y(n_727) );
INVx1_ASAP7_75t_SL g728 ( .A(n_646), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_620), .A2(n_469), .B1(n_473), .B2(n_407), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_688), .Y(n_730) );
NOR2x1_ASAP7_75t_R g731 ( .A(n_663), .B(n_500), .Y(n_731) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_634), .A2(n_398), .B(n_367), .Y(n_732) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_614), .Y(n_733) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_614), .Y(n_734) );
INVx8_ASAP7_75t_L g735 ( .A(n_625), .Y(n_735) );
INVx3_ASAP7_75t_L g736 ( .A(n_626), .Y(n_736) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_625), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_657), .B(n_467), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_623), .A2(n_475), .B1(n_489), .B2(n_486), .Y(n_739) );
INVx4_ASAP7_75t_L g740 ( .A(n_625), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_679), .A2(n_481), .B1(n_514), .B2(n_448), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_693), .Y(n_742) );
BUFx3_ASAP7_75t_L g743 ( .A(n_622), .Y(n_743) );
CKINVDCx5p33_ASAP7_75t_R g744 ( .A(n_612), .Y(n_744) );
BUFx2_ASAP7_75t_L g745 ( .A(n_669), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_673), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g747 ( .A(n_635), .B(n_405), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_656), .A2(n_492), .B1(n_499), .B2(n_493), .C(n_491), .Y(n_748) );
HAxp5_ASAP7_75t_L g749 ( .A(n_652), .B(n_388), .CON(n_749), .SN(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_679), .B(n_505), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_649), .B(n_682), .Y(n_751) );
AND2x4_ASAP7_75t_L g752 ( .A(n_619), .B(n_502), .Y(n_752) );
O2A1O1Ixp5_ASAP7_75t_L g753 ( .A1(n_655), .A2(n_522), .B(n_363), .C(n_454), .Y(n_753) );
AND2x2_ASAP7_75t_SL g754 ( .A(n_647), .B(n_519), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_628), .B(n_409), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_692), .B(n_418), .Y(n_756) );
O2A1O1Ixp33_ASAP7_75t_L g757 ( .A1(n_628), .A2(n_530), .B(n_387), .C(n_390), .Y(n_757) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_658), .Y(n_758) );
AND2x4_ASAP7_75t_SL g759 ( .A(n_635), .B(n_508), .Y(n_759) );
INVx1_ASAP7_75t_SL g760 ( .A(n_635), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_629), .A2(n_386), .B1(n_393), .B2(n_392), .Y(n_761) );
INVx3_ASAP7_75t_L g762 ( .A(n_633), .Y(n_762) );
BUFx6f_ASAP7_75t_L g763 ( .A(n_642), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_623), .B(n_409), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_693), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_683), .B(n_442), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_683), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_642), .B(n_442), .Y(n_768) );
BUFx2_ASAP7_75t_L g769 ( .A(n_659), .Y(n_769) );
AND2x4_ASAP7_75t_L g770 ( .A(n_619), .B(n_395), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_677), .A2(n_399), .B1(n_410), .B2(n_406), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_645), .B(n_671), .Y(n_772) );
INVx6_ASAP7_75t_L g773 ( .A(n_681), .Y(n_773) );
NAND2xp5_ASAP7_75t_SL g774 ( .A(n_642), .B(n_452), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_612), .B(n_452), .Y(n_775) );
BUFx2_ASAP7_75t_L g776 ( .A(n_658), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_645), .B(n_471), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_684), .B(n_471), .Y(n_778) );
BUFx2_ASAP7_75t_L g779 ( .A(n_687), .Y(n_779) );
AND2x4_ASAP7_75t_L g780 ( .A(n_675), .B(n_415), .Y(n_780) );
INVxp67_ASAP7_75t_L g781 ( .A(n_638), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_648), .A2(n_508), .B1(n_563), .B2(n_555), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_699), .Y(n_783) );
INVxp67_ASAP7_75t_L g784 ( .A(n_662), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_691), .A2(n_690), .B1(n_674), .B2(n_686), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_655), .A2(n_609), .B(n_422), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_670), .A2(n_428), .B(n_421), .Y(n_787) );
AND2x4_ASAP7_75t_L g788 ( .A(n_702), .B(n_429), .Y(n_788) );
INVxp67_ASAP7_75t_L g789 ( .A(n_698), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_700), .B(n_479), .Y(n_790) );
BUFx4f_ASAP7_75t_L g791 ( .A(n_651), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_670), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_618), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_661), .A2(n_431), .B1(n_438), .B2(n_434), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_676), .Y(n_795) );
INVx3_ASAP7_75t_L g796 ( .A(n_633), .Y(n_796) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_639), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_676), .A2(n_440), .B(n_439), .Y(n_798) );
INVx2_ASAP7_75t_SL g799 ( .A(n_636), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_695), .Y(n_800) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_641), .Y(n_801) );
BUFx6f_ASAP7_75t_SL g802 ( .A(n_617), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_701), .A2(n_508), .B1(n_563), .B2(n_555), .Y(n_803) );
INVx1_ASAP7_75t_SL g804 ( .A(n_704), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_697), .B(n_490), .Y(n_805) );
BUFx6f_ASAP7_75t_L g806 ( .A(n_681), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_680), .Y(n_807) );
BUFx2_ASAP7_75t_L g808 ( .A(n_651), .Y(n_808) );
NAND2x1p5_ASAP7_75t_L g809 ( .A(n_681), .B(n_508), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_643), .B(n_490), .Y(n_810) );
BUFx2_ASAP7_75t_L g811 ( .A(n_651), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_680), .Y(n_812) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_681), .Y(n_813) );
INVx5_ASAP7_75t_L g814 ( .A(n_651), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_650), .B(n_498), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_636), .B(n_498), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_661), .A2(n_443), .B(n_441), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_621), .Y(n_818) );
BUFx6f_ASAP7_75t_L g819 ( .A(n_653), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_664), .A2(n_453), .B(n_450), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_667), .Y(n_821) );
INVx3_ASAP7_75t_L g822 ( .A(n_630), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_668), .A2(n_462), .B1(n_464), .B2(n_459), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_668), .A2(n_470), .B1(n_474), .B2(n_466), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_703), .A2(n_478), .B(n_477), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_666), .B(n_501), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_637), .B(n_501), .Y(n_827) );
BUFx3_ASAP7_75t_L g828 ( .A(n_654), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_672), .Y(n_829) );
BUFx2_ASAP7_75t_L g830 ( .A(n_678), .Y(n_830) );
BUFx6f_ASAP7_75t_L g831 ( .A(n_614), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_613), .Y(n_832) );
INVx3_ASAP7_75t_L g833 ( .A(n_626), .Y(n_833) );
NAND3xp33_ASAP7_75t_L g834 ( .A(n_629), .B(n_563), .C(n_555), .Y(n_834) );
INVx4_ASAP7_75t_L g835 ( .A(n_616), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_615), .A2(n_482), .B1(n_483), .B2(n_480), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_696), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_644), .B(n_503), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_644), .B(n_503), .Y(n_839) );
CKINVDCx11_ASAP7_75t_R g840 ( .A(n_622), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_696), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_615), .B(n_518), .Y(n_842) );
AOI221xp5_ASAP7_75t_L g843 ( .A1(n_613), .A2(n_518), .B1(n_495), .B2(n_515), .C(n_513), .Y(n_843) );
OR2x6_ASAP7_75t_L g844 ( .A(n_612), .B(n_416), .Y(n_844) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_613), .Y(n_845) );
BUFx3_ASAP7_75t_L g846 ( .A(n_613), .Y(n_846) );
INVx1_ASAP7_75t_SL g847 ( .A(n_728), .Y(n_847) );
INVx6_ASAP7_75t_L g848 ( .A(n_835), .Y(n_848) );
AO21x2_ASAP7_75t_L g849 ( .A1(n_834), .A2(n_517), .B(n_494), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_792), .B(n_520), .Y(n_850) );
AND2x4_ASAP7_75t_L g851 ( .A(n_835), .B(n_521), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_751), .A2(n_563), .B1(n_512), .B2(n_506), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_845), .Y(n_853) );
OA21x2_ASAP7_75t_L g854 ( .A1(n_834), .A2(n_485), .B(n_411), .Y(n_854) );
BUFx6f_ASAP7_75t_L g855 ( .A(n_806), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_705), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_728), .B(n_9), .Y(n_857) );
AND2x4_ASAP7_75t_L g858 ( .A(n_708), .B(n_512), .Y(n_858) );
AND2x4_ASAP7_75t_L g859 ( .A(n_711), .B(n_485), .Y(n_859) );
NAND2x1p5_ASAP7_75t_L g860 ( .A(n_776), .B(n_389), .Y(n_860) );
CKINVDCx6p67_ASAP7_75t_R g861 ( .A(n_840), .Y(n_861) );
O2A1O1Ixp33_ASAP7_75t_SL g862 ( .A1(n_715), .A2(n_525), .B(n_539), .C(n_538), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_846), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_709), .B(n_838), .Y(n_864) );
AO21x2_ASAP7_75t_L g865 ( .A1(n_786), .A2(n_538), .B(n_525), .Y(n_865) );
INVx3_ASAP7_75t_L g866 ( .A(n_806), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_819), .Y(n_867) );
OR2x2_ASAP7_75t_L g868 ( .A(n_719), .B(n_10), .Y(n_868) );
OAI22xp33_ASAP7_75t_L g869 ( .A1(n_744), .A2(n_563), .B1(n_504), .B2(n_420), .Y(n_869) );
BUFx4f_ASAP7_75t_SL g870 ( .A(n_727), .Y(n_870) );
BUFx2_ASAP7_75t_L g871 ( .A(n_743), .Y(n_871) );
INVx2_ASAP7_75t_SL g872 ( .A(n_717), .Y(n_872) );
BUFx2_ASAP7_75t_L g873 ( .A(n_746), .Y(n_873) );
OAI21x1_ASAP7_75t_L g874 ( .A1(n_809), .A2(n_570), .B(n_564), .Y(n_874) );
OAI21xp5_ASAP7_75t_L g875 ( .A1(n_753), .A2(n_592), .B(n_573), .Y(n_875) );
OAI21xp5_ASAP7_75t_L g876 ( .A1(n_817), .A2(n_592), .B(n_573), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_832), .Y(n_877) );
AO21x2_ASAP7_75t_L g878 ( .A1(n_820), .A2(n_539), .B(n_538), .Y(n_878) );
AO31x2_ASAP7_75t_L g879 ( .A1(n_794), .A2(n_545), .A3(n_548), .B(n_539), .Y(n_879) );
O2A1O1Ixp33_ASAP7_75t_SL g880 ( .A1(n_716), .A2(n_548), .B(n_545), .C(n_107), .Y(n_880) );
OAI21x1_ASAP7_75t_L g881 ( .A1(n_718), .A2(n_600), .B(n_574), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_797), .Y(n_882) );
OAI21x1_ASAP7_75t_SL g883 ( .A1(n_799), .A2(n_10), .B(n_11), .Y(n_883) );
AO21x2_ASAP7_75t_L g884 ( .A1(n_823), .A2(n_553), .B(n_551), .Y(n_884) );
AOI21x1_ASAP7_75t_L g885 ( .A1(n_794), .A2(n_600), .B(n_574), .Y(n_885) );
OAI21x1_ASAP7_75t_L g886 ( .A1(n_822), .A2(n_600), .B(n_574), .Y(n_886) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_758), .Y(n_887) );
AOI21xp33_ASAP7_75t_L g888 ( .A1(n_757), .A2(n_600), .B(n_574), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_754), .A2(n_423), .B1(n_432), .B2(n_351), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_801), .Y(n_890) );
OAI21x1_ASAP7_75t_L g891 ( .A1(n_822), .A2(n_600), .B(n_574), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_830), .Y(n_892) );
AO21x2_ASAP7_75t_L g893 ( .A1(n_823), .A2(n_553), .B(n_551), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_795), .B(n_574), .Y(n_894) );
AO32x2_ASAP7_75t_L g895 ( .A1(n_824), .A2(n_551), .A3(n_553), .B1(n_600), .B2(n_15), .Y(n_895) );
AOI22xp33_ASAP7_75t_SL g896 ( .A1(n_844), .A2(n_13), .B1(n_11), .B2(n_12), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_807), .A2(n_553), .B1(n_551), .B2(n_578), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_802), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_821), .Y(n_899) );
BUFx3_ASAP7_75t_L g900 ( .A(n_745), .Y(n_900) );
OAI21xp5_ASAP7_75t_L g901 ( .A1(n_812), .A2(n_553), .B(n_551), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_839), .B(n_13), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g903 ( .A1(n_775), .A2(n_553), .B1(n_551), .B2(n_578), .Y(n_903) );
AO21x2_ASAP7_75t_L g904 ( .A1(n_824), .A2(n_605), .B(n_578), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_784), .B(n_16), .Y(n_905) );
AO21x2_ASAP7_75t_L g906 ( .A1(n_787), .A2(n_605), .B(n_578), .Y(n_906) );
OAI21x1_ASAP7_75t_L g907 ( .A1(n_798), .A2(n_110), .B(n_106), .Y(n_907) );
OAI21x1_ASAP7_75t_L g908 ( .A1(n_825), .A2(n_113), .B(n_111), .Y(n_908) );
BUFx3_ASAP7_75t_L g909 ( .A(n_806), .Y(n_909) );
OAI21xp5_ASAP7_75t_L g910 ( .A1(n_732), .A2(n_16), .B(n_17), .Y(n_910) );
OAI21x1_ASAP7_75t_L g911 ( .A1(n_707), .A2(n_116), .B(n_114), .Y(n_911) );
NAND2x1p5_ASAP7_75t_L g912 ( .A(n_814), .B(n_17), .Y(n_912) );
NAND2xp5_ASAP7_75t_SL g913 ( .A(n_819), .B(n_605), .Y(n_913) );
OAI21x1_ASAP7_75t_L g914 ( .A1(n_712), .A2(n_118), .B(n_117), .Y(n_914) );
BUFx2_ASAP7_75t_L g915 ( .A(n_719), .Y(n_915) );
INVxp67_ASAP7_75t_L g916 ( .A(n_714), .Y(n_916) );
AO21x1_ASAP7_75t_L g917 ( .A1(n_788), .A2(n_120), .B(n_119), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_767), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_772), .B(n_18), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_772), .B(n_18), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_829), .Y(n_921) );
OAI21x1_ASAP7_75t_L g922 ( .A1(n_783), .A2(n_125), .B(n_124), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g923 ( .A(n_802), .Y(n_923) );
OAI21x1_ASAP7_75t_L g924 ( .A1(n_837), .A2(n_128), .B(n_127), .Y(n_924) );
AND2x4_ASAP7_75t_L g925 ( .A(n_713), .B(n_19), .Y(n_925) );
OAI21x1_ASAP7_75t_L g926 ( .A1(n_841), .A2(n_137), .B(n_135), .Y(n_926) );
CKINVDCx14_ASAP7_75t_R g927 ( .A(n_793), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_730), .Y(n_928) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_813), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_752), .Y(n_930) );
INVx2_ASAP7_75t_SL g931 ( .A(n_773), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_748), .B(n_19), .Y(n_932) );
AOI21xp5_ASAP7_75t_L g933 ( .A1(n_842), .A2(n_605), .B(n_578), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_723), .B(n_20), .Y(n_934) );
AOI21xp5_ASAP7_75t_L g935 ( .A1(n_818), .A2(n_605), .B(n_578), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g936 ( .A1(n_755), .A2(n_605), .B(n_140), .Y(n_936) );
OAI21x1_ASAP7_75t_L g937 ( .A1(n_800), .A2(n_141), .B(n_139), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_844), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_938) );
AOI21x1_ASAP7_75t_L g939 ( .A1(n_788), .A2(n_146), .B(n_143), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_771), .B(n_21), .Y(n_940) );
OAI21xp5_ASAP7_75t_L g941 ( .A1(n_771), .A2(n_22), .B(n_23), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_752), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_742), .Y(n_943) );
BUFx6f_ASAP7_75t_L g944 ( .A(n_813), .Y(n_944) );
OAI21x1_ASAP7_75t_L g945 ( .A1(n_803), .A2(n_151), .B(n_148), .Y(n_945) );
OAI21x1_ASAP7_75t_L g946 ( .A1(n_782), .A2(n_768), .B(n_747), .Y(n_946) );
A2O1A1Ixp33_ASAP7_75t_L g947 ( .A1(n_761), .A2(n_23), .B(n_24), .C(n_25), .Y(n_947) );
BUFx12f_ASAP7_75t_L g948 ( .A(n_844), .Y(n_948) );
OAI21x1_ASAP7_75t_L g949 ( .A1(n_774), .A2(n_156), .B(n_155), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_819), .Y(n_950) );
NAND3xp33_ASAP7_75t_L g951 ( .A(n_756), .B(n_25), .C(n_26), .Y(n_951) );
HB1xp67_ASAP7_75t_L g952 ( .A(n_813), .Y(n_952) );
INVx4_ASAP7_75t_L g953 ( .A(n_735), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_723), .B(n_26), .Y(n_954) );
CKINVDCx16_ASAP7_75t_R g955 ( .A(n_779), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_765), .Y(n_956) );
AND2x4_ASAP7_75t_L g957 ( .A(n_789), .B(n_27), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_722), .B(n_27), .Y(n_958) );
AND2x4_ASAP7_75t_L g959 ( .A(n_814), .B(n_28), .Y(n_959) );
OAI21x1_ASAP7_75t_L g960 ( .A1(n_726), .A2(n_159), .B(n_157), .Y(n_960) );
INVx3_ASAP7_75t_L g961 ( .A(n_773), .Y(n_961) );
BUFx8_ASAP7_75t_L g962 ( .A(n_769), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_828), .Y(n_963) );
A2O1A1Ixp33_ASAP7_75t_L g964 ( .A1(n_761), .A2(n_28), .B(n_32), .C(n_33), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_764), .B(n_32), .Y(n_965) );
OA21x2_ASAP7_75t_L g966 ( .A1(n_836), .A2(n_162), .B(n_160), .Y(n_966) );
INVx2_ASAP7_75t_L g967 ( .A(n_726), .Y(n_967) );
INVx2_ASAP7_75t_SL g968 ( .A(n_720), .Y(n_968) );
A2O1A1Ixp33_ASAP7_75t_L g969 ( .A1(n_781), .A2(n_33), .B(n_34), .C(n_35), .Y(n_969) );
AOI22xp5_ASAP7_75t_L g970 ( .A1(n_804), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_804), .Y(n_971) );
OA21x2_ASAP7_75t_L g972 ( .A1(n_836), .A2(n_164), .B(n_163), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_720), .B(n_36), .Y(n_973) );
A2O1A1Ixp33_ASAP7_75t_L g974 ( .A1(n_827), .A2(n_37), .B(n_39), .C(n_40), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_710), .B(n_39), .Y(n_975) );
OA21x2_ASAP7_75t_L g976 ( .A1(n_810), .A2(n_168), .B(n_167), .Y(n_976) );
INVx2_ASAP7_75t_L g977 ( .A(n_736), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_770), .Y(n_978) );
OAI21x1_ASAP7_75t_L g979 ( .A1(n_736), .A2(n_174), .B(n_169), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_791), .A2(n_41), .B1(n_42), .B2(n_44), .Y(n_980) );
AOI21x1_ASAP7_75t_L g981 ( .A1(n_808), .A2(n_176), .B(n_175), .Y(n_981) );
AO21x2_ASAP7_75t_L g982 ( .A1(n_739), .A2(n_180), .B(n_178), .Y(n_982) );
OA21x2_ASAP7_75t_L g983 ( .A1(n_815), .A2(n_183), .B(n_182), .Y(n_983) );
OAI222xp33_ASAP7_75t_L g984 ( .A1(n_725), .A2(n_42), .B1(n_44), .B2(n_48), .C1(n_49), .C2(n_50), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_706), .B(n_48), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_826), .B(n_49), .Y(n_986) );
AO31x2_ASAP7_75t_L g987 ( .A1(n_739), .A2(n_50), .A3(n_51), .B(n_52), .Y(n_987) );
OAI221xp5_ASAP7_75t_L g988 ( .A1(n_843), .A2(n_51), .B1(n_52), .B2(n_53), .C(n_55), .Y(n_988) );
BUFx3_ASAP7_75t_L g989 ( .A(n_735), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_770), .B(n_55), .Y(n_990) );
INVx2_ASAP7_75t_L g991 ( .A(n_762), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_766), .Y(n_992) );
OA21x2_ASAP7_75t_L g993 ( .A1(n_778), .A2(n_185), .B(n_184), .Y(n_993) );
OAI21x1_ASAP7_75t_SL g994 ( .A1(n_740), .A2(n_56), .B(n_57), .Y(n_994) );
A2O1A1Ixp33_ASAP7_75t_L g995 ( .A1(n_741), .A2(n_791), .B(n_790), .C(n_750), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_814), .A2(n_57), .B1(n_58), .B2(n_59), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g997 ( .A1(n_816), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_997) );
INVx4_ASAP7_75t_L g998 ( .A(n_735), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_729), .Y(n_999) );
OAI21x1_ASAP7_75t_SL g1000 ( .A1(n_740), .A2(n_60), .B(n_61), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_729), .Y(n_1001) );
AOI21xp5_ASAP7_75t_L g1002 ( .A1(n_805), .A2(n_190), .B(n_188), .Y(n_1002) );
OAI211xp5_ASAP7_75t_SL g1003 ( .A1(n_738), .A2(n_61), .B(n_62), .C(n_63), .Y(n_1003) );
OA21x2_ASAP7_75t_L g1004 ( .A1(n_780), .A2(n_235), .B(n_344), .Y(n_1004) );
AO21x2_ASAP7_75t_L g1005 ( .A1(n_741), .A2(n_234), .B(n_343), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_749), .B(n_62), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_777), .B(n_63), .Y(n_1007) );
NAND2x1p5_ASAP7_75t_L g1008 ( .A(n_721), .B(n_65), .Y(n_1008) );
CKINVDCx20_ASAP7_75t_R g1009 ( .A(n_724), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_780), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_811), .Y(n_1011) );
NAND2x1p5_ASAP7_75t_L g1012 ( .A(n_721), .B(n_65), .Y(n_1012) );
OAI22xp5_ASAP7_75t_SL g1013 ( .A1(n_731), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1014 ( .A(n_971), .Y(n_1014) );
OR2x2_ASAP7_75t_L g1015 ( .A(n_915), .B(n_731), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_861), .Y(n_1016) );
AOI21xp5_ASAP7_75t_L g1017 ( .A1(n_933), .A2(n_760), .B(n_759), .Y(n_1017) );
AND2x4_ASAP7_75t_L g1018 ( .A(n_916), .B(n_762), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_999), .B(n_796), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_899), .Y(n_1020) );
INVx3_ASAP7_75t_L g1021 ( .A(n_953), .Y(n_1021) );
AND2x4_ASAP7_75t_L g1022 ( .A(n_916), .B(n_796), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_850), .A2(n_785), .B1(n_760), .B2(n_831), .Y(n_1023) );
AOI222xp33_ASAP7_75t_L g1024 ( .A1(n_934), .A2(n_833), .B1(n_831), .B2(n_763), .C1(n_737), .C2(n_734), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_954), .A2(n_1001), .B1(n_948), .B2(n_957), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_957), .A2(n_833), .B1(n_831), .B2(n_763), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_877), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_853), .Y(n_1028) );
AOI222xp33_ASAP7_75t_L g1029 ( .A1(n_1013), .A2(n_763), .B1(n_737), .B2(n_734), .C1(n_733), .C2(n_721), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_847), .B(n_68), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_850), .A2(n_734), .B1(n_733), .B2(n_737), .Y(n_1031) );
AOI31xp33_ASAP7_75t_L g1032 ( .A1(n_860), .A2(n_69), .A3(n_71), .B(n_74), .Y(n_1032) );
OR2x6_ASAP7_75t_L g1033 ( .A(n_860), .B(n_733), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_921), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_919), .A2(n_69), .B1(n_75), .B2(n_77), .Y(n_1035) );
AOI221xp5_ASAP7_75t_L g1036 ( .A1(n_992), .A2(n_75), .B1(n_78), .B2(n_79), .C(n_80), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_864), .B(n_78), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_847), .B(n_79), .Y(n_1038) );
AOI222xp33_ASAP7_75t_L g1039 ( .A1(n_985), .A2(n_81), .B1(n_82), .B2(n_83), .C1(n_84), .C2(n_85), .Y(n_1039) );
OAI321xp33_ASAP7_75t_L g1040 ( .A1(n_980), .A2(n_81), .A3(n_83), .B1(n_85), .B2(n_87), .C(n_88), .Y(n_1040) );
OAI211xp5_ASAP7_75t_L g1041 ( .A1(n_896), .A2(n_87), .B(n_89), .C(n_90), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_919), .A2(n_91), .B1(n_92), .B2(n_94), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_940), .A2(n_92), .B1(n_94), .B2(n_95), .Y(n_1043) );
OAI21xp5_ASAP7_75t_SL g1044 ( .A1(n_984), .A2(n_95), .B(n_96), .Y(n_1044) );
OR2x2_ASAP7_75t_L g1045 ( .A(n_887), .B(n_98), .Y(n_1045) );
AOI21xp5_ASAP7_75t_L g1046 ( .A1(n_995), .A2(n_259), .B(n_341), .Y(n_1046) );
A2O1A1Ixp33_ASAP7_75t_L g1047 ( .A1(n_941), .A2(n_98), .B(n_99), .C(n_100), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_988), .A2(n_99), .B1(n_100), .B2(n_101), .Y(n_1048) );
OAI22xp33_ASAP7_75t_L g1049 ( .A1(n_868), .A2(n_102), .B1(n_103), .B2(n_191), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_971), .B(n_102), .Y(n_1050) );
OAI21xp33_ASAP7_75t_SL g1051 ( .A1(n_941), .A2(n_192), .B(n_193), .Y(n_1051) );
AOI21xp33_ASAP7_75t_L g1052 ( .A1(n_975), .A2(n_346), .B(n_194), .Y(n_1052) );
AOI21xp33_ASAP7_75t_L g1053 ( .A1(n_975), .A2(n_340), .B(n_198), .Y(n_1053) );
CKINVDCx5p33_ASAP7_75t_R g1054 ( .A(n_856), .Y(n_1054) );
BUFx6f_ASAP7_75t_L g1055 ( .A(n_855), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_932), .B(n_338), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_1006), .A2(n_196), .B1(n_201), .B2(n_202), .Y(n_1057) );
INVxp67_ASAP7_75t_SL g1058 ( .A(n_925), .Y(n_1058) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_887), .Y(n_1059) );
AOI22xp33_ASAP7_75t_SL g1060 ( .A1(n_955), .A2(n_203), .B1(n_205), .B2(n_207), .Y(n_1060) );
OAI221xp5_ASAP7_75t_L g1061 ( .A1(n_905), .A2(n_208), .B1(n_210), .B2(n_211), .C(n_212), .Y(n_1061) );
AOI211xp5_ASAP7_75t_L g1062 ( .A1(n_980), .A2(n_214), .B(n_215), .C(n_219), .Y(n_1062) );
INVx3_ASAP7_75t_L g1063 ( .A(n_953), .Y(n_1063) );
NAND4xp25_ASAP7_75t_L g1064 ( .A(n_896), .B(n_220), .C(n_223), .D(n_225), .Y(n_1064) );
AND2x4_ASAP7_75t_L g1065 ( .A(n_998), .B(n_230), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_882), .Y(n_1066) );
OAI221xp5_ASAP7_75t_L g1067 ( .A1(n_905), .A2(n_233), .B1(n_236), .B2(n_237), .C(n_238), .Y(n_1067) );
HB1xp67_ASAP7_75t_L g1068 ( .A(n_873), .Y(n_1068) );
OAI221xp5_ASAP7_75t_SL g1069 ( .A1(n_938), .A2(n_239), .B1(n_242), .B2(n_245), .C(n_246), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_892), .B(n_250), .Y(n_1070) );
INVx11_ASAP7_75t_L g1071 ( .A(n_962), .Y(n_1071) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_890), .B(n_253), .Y(n_1072) );
INVx3_ASAP7_75t_L g1073 ( .A(n_998), .Y(n_1073) );
OR2x2_ASAP7_75t_L g1074 ( .A(n_990), .B(n_255), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_932), .B(n_336), .Y(n_1075) );
AOI21xp5_ASAP7_75t_L g1076 ( .A1(n_935), .A2(n_257), .B(n_260), .Y(n_1076) );
OAI222xp33_ASAP7_75t_L g1077 ( .A1(n_988), .A2(n_261), .B1(n_264), .B2(n_265), .C1(n_266), .C2(n_268), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1078 ( .A(n_990), .B(n_269), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_902), .A2(n_270), .B1(n_271), .B2(n_276), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_940), .A2(n_277), .B1(n_278), .B2(n_282), .Y(n_1080) );
OAI221xp5_ASAP7_75t_L g1081 ( .A1(n_968), .A2(n_978), .B1(n_930), .B2(n_942), .C(n_938), .Y(n_1081) );
OAI22xp33_ASAP7_75t_L g1082 ( .A1(n_870), .A2(n_284), .B1(n_285), .B2(n_286), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_925), .Y(n_1083) );
AOI21xp5_ASAP7_75t_L g1084 ( .A1(n_935), .A2(n_288), .B(n_296), .Y(n_1084) );
CKINVDCx5p33_ASAP7_75t_R g1085 ( .A(n_898), .Y(n_1085) );
AOI21xp5_ASAP7_75t_L g1086 ( .A1(n_913), .A2(n_299), .B(n_304), .Y(n_1086) );
AO31x2_ASAP7_75t_L g1087 ( .A1(n_917), .A2(n_305), .A3(n_308), .B(n_309), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_943), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_986), .A2(n_310), .B1(n_311), .B2(n_312), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_973), .B(n_334), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_958), .A2(n_314), .B1(n_317), .B2(n_318), .Y(n_1091) );
A2O1A1Ixp33_ASAP7_75t_L g1092 ( .A1(n_910), .A2(n_319), .B(n_322), .C(n_324), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_958), .A2(n_326), .B1(n_327), .B2(n_328), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_857), .B(n_333), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1007), .B(n_330), .Y(n_1095) );
INVx2_ASAP7_75t_L g1096 ( .A(n_918), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_956), .Y(n_1097) );
OAI21xp33_ASAP7_75t_L g1098 ( .A1(n_1003), .A2(n_332), .B(n_910), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_928), .Y(n_1099) );
A2O1A1Ixp33_ASAP7_75t_L g1100 ( .A1(n_965), .A2(n_951), .B(n_947), .C(n_974), .Y(n_1100) );
INVx3_ASAP7_75t_L g1101 ( .A(n_855), .Y(n_1101) );
AOI22xp33_ASAP7_75t_SL g1102 ( .A1(n_962), .A2(n_870), .B1(n_996), .B2(n_959), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_920), .Y(n_1103) );
AO31x2_ASAP7_75t_L g1104 ( .A1(n_897), .A2(n_936), .A3(n_1002), .B(n_947), .Y(n_1104) );
INVx3_ASAP7_75t_L g1105 ( .A(n_855), .Y(n_1105) );
A2O1A1Ixp33_ASAP7_75t_L g1106 ( .A1(n_965), .A2(n_1003), .B(n_969), .C(n_964), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_863), .B(n_1010), .Y(n_1107) );
AOI22xp33_ASAP7_75t_SL g1108 ( .A1(n_996), .A2(n_959), .B1(n_912), .B2(n_883), .Y(n_1108) );
NAND3xp33_ASAP7_75t_L g1109 ( .A(n_903), .B(n_1002), .C(n_997), .Y(n_1109) );
AOI21xp5_ASAP7_75t_L g1110 ( .A1(n_913), .A2(n_875), .B(n_936), .Y(n_1110) );
AND2x4_ASAP7_75t_L g1111 ( .A(n_909), .B(n_989), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_859), .B(n_858), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_920), .B(n_963), .Y(n_1113) );
BUFx8_ASAP7_75t_SL g1114 ( .A(n_871), .Y(n_1114) );
OAI22xp33_ASAP7_75t_L g1115 ( .A1(n_889), .A2(n_970), .B1(n_912), .B2(n_848), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_851), .A2(n_859), .B1(n_858), .B2(n_1009), .Y(n_1116) );
OAI22xp33_ASAP7_75t_L g1117 ( .A1(n_848), .A2(n_900), .B1(n_1012), .B2(n_1008), .Y(n_1117) );
AOI221xp5_ASAP7_75t_SL g1118 ( .A1(n_869), .A2(n_984), .B1(n_852), .B2(n_901), .C(n_897), .Y(n_1118) );
NOR2xp33_ASAP7_75t_L g1119 ( .A(n_851), .B(n_872), .Y(n_1119) );
OAI22xp5_ASAP7_75t_L g1120 ( .A1(n_869), .A2(n_852), .B1(n_1012), .B2(n_1008), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_1011), .A2(n_848), .B1(n_931), .B2(n_961), .Y(n_1121) );
INVx3_ASAP7_75t_L g1122 ( .A(n_944), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_929), .B(n_952), .Y(n_1123) );
OAI22xp33_ASAP7_75t_L g1124 ( .A1(n_894), .A2(n_923), .B1(n_1011), .B2(n_966), .Y(n_1124) );
AOI22xp5_ASAP7_75t_L g1125 ( .A1(n_894), .A2(n_982), .B1(n_966), .B2(n_972), .Y(n_1125) );
AOI22xp33_ASAP7_75t_SL g1126 ( .A1(n_994), .A2(n_1000), .B1(n_972), .B2(n_982), .Y(n_1126) );
AOI221xp5_ASAP7_75t_L g1127 ( .A1(n_862), .A2(n_927), .B1(n_888), .B2(n_880), .C(n_961), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_929), .B(n_952), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_987), .Y(n_1129) );
AOI221xp5_ASAP7_75t_L g1130 ( .A1(n_862), .A2(n_888), .B1(n_880), .B2(n_967), .C(n_991), .Y(n_1130) );
OAI21xp5_ASAP7_75t_L g1131 ( .A1(n_946), .A2(n_881), .B(n_885), .Y(n_1131) );
OAI221xp5_ASAP7_75t_L g1132 ( .A1(n_875), .A2(n_977), .B1(n_876), .B2(n_866), .C(n_854), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_987), .B(n_866), .Y(n_1133) );
INVxp67_ASAP7_75t_L g1134 ( .A(n_944), .Y(n_1134) );
NAND4xp25_ASAP7_75t_L g1135 ( .A(n_876), .B(n_987), .C(n_867), .D(n_950), .Y(n_1135) );
INVx1_ASAP7_75t_SL g1136 ( .A(n_944), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_895), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_1004), .A2(n_854), .B1(n_993), .B2(n_976), .Y(n_1138) );
OAI22xp5_ASAP7_75t_L g1139 ( .A1(n_1004), .A2(n_993), .B1(n_976), .B2(n_983), .Y(n_1139) );
AO22x1_ASAP7_75t_L g1140 ( .A1(n_895), .A2(n_1005), .B1(n_939), .B2(n_893), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_983), .A2(n_981), .B1(n_895), .B2(n_904), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_904), .B(n_878), .Y(n_1142) );
BUFx2_ASAP7_75t_L g1143 ( .A(n_886), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_895), .B(n_879), .Y(n_1144) );
NOR2xp33_ASAP7_75t_L g1145 ( .A(n_849), .B(n_878), .Y(n_1145) );
AOI22xp33_ASAP7_75t_SL g1146 ( .A1(n_1005), .A2(n_893), .B1(n_884), .B2(n_979), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_879), .Y(n_1147) );
AO21x2_ASAP7_75t_L g1148 ( .A1(n_884), .A2(n_849), .B(n_906), .Y(n_1148) );
OAI22xp33_ASAP7_75t_L g1149 ( .A1(n_960), .A2(n_879), .B1(n_907), .B2(n_908), .Y(n_1149) );
BUFx2_ASAP7_75t_L g1150 ( .A(n_891), .Y(n_1150) );
INVx3_ASAP7_75t_L g1151 ( .A(n_874), .Y(n_1151) );
OAI22xp33_ASAP7_75t_L g1152 ( .A1(n_945), .A2(n_949), .B1(n_937), .B2(n_911), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_865), .Y(n_1153) );
OAI321xp33_ASAP7_75t_L g1154 ( .A1(n_914), .A2(n_980), .A3(n_1003), .B1(n_941), .B2(n_996), .C(n_1013), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_922), .B(n_924), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_926), .A2(n_844), .B1(n_754), .B2(n_632), .Y(n_1156) );
INVx2_ASAP7_75t_L g1157 ( .A(n_899), .Y(n_1157) );
OAI22xp5_ASAP7_75t_L g1158 ( .A1(n_915), .A2(n_612), .B1(n_744), .B2(n_728), .Y(n_1158) );
OAI221xp5_ASAP7_75t_L g1159 ( .A1(n_999), .A2(n_751), .B1(n_644), .B2(n_646), .C(n_725), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_877), .Y(n_1160) );
AOI21xp33_ASAP7_75t_L g1161 ( .A1(n_975), .A2(n_751), .B(n_757), .Y(n_1161) );
AND2x4_ASAP7_75t_L g1162 ( .A(n_916), .B(n_835), .Y(n_1162) );
NAND3xp33_ASAP7_75t_L g1163 ( .A(n_951), .B(n_753), .C(n_974), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_877), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_877), .Y(n_1165) );
OAI211xp5_ASAP7_75t_SL g1166 ( .A1(n_930), .A2(n_618), .B(n_723), .C(n_725), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1019), .Y(n_1167) );
INVx2_ASAP7_75t_SL g1168 ( .A(n_1021), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1103), .B(n_1020), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1129), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_1102), .A2(n_1159), .B1(n_1025), .B2(n_1166), .Y(n_1171) );
AOI22xp5_ASAP7_75t_L g1172 ( .A1(n_1044), .A2(n_1158), .B1(n_1048), .B2(n_1039), .Y(n_1172) );
INVx4_ASAP7_75t_L g1173 ( .A(n_1055), .Y(n_1173) );
BUFx2_ASAP7_75t_L g1174 ( .A(n_1143), .Y(n_1174) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1153), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1137), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1147), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1133), .Y(n_1178) );
INVx3_ASAP7_75t_L g1179 ( .A(n_1055), .Y(n_1179) );
NOR2xp33_ASAP7_75t_L g1180 ( .A(n_1015), .B(n_1112), .Y(n_1180) );
INVx2_ASAP7_75t_L g1181 ( .A(n_1148), .Y(n_1181) );
AND2x4_ASAP7_75t_L g1182 ( .A(n_1101), .B(n_1105), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_1161), .A2(n_1156), .B1(n_1098), .B2(n_1081), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1027), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1160), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1164), .B(n_1165), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1157), .B(n_1034), .Y(n_1187) );
NOR2x1_ASAP7_75t_L g1188 ( .A(n_1135), .B(n_1117), .Y(n_1188) );
BUFx3_ASAP7_75t_L g1189 ( .A(n_1021), .Y(n_1189) );
OR2x2_ASAP7_75t_L g1190 ( .A(n_1014), .B(n_1058), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1123), .B(n_1096), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1088), .B(n_1097), .Y(n_1192) );
HB1xp67_ASAP7_75t_L g1193 ( .A(n_1059), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g1194 ( .A1(n_1098), .A2(n_1108), .B1(n_1115), .B2(n_1048), .Y(n_1194) );
BUFx3_ASAP7_75t_L g1195 ( .A(n_1063), .Y(n_1195) );
NAND2xp5_ASAP7_75t_SL g1196 ( .A(n_1029), .B(n_1062), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1099), .B(n_1028), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1144), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1142), .Y(n_1199) );
OR2x6_ASAP7_75t_L g1200 ( .A(n_1120), .B(n_1033), .Y(n_1200) );
INVx2_ASAP7_75t_L g1201 ( .A(n_1055), .Y(n_1201) );
HB1xp67_ASAP7_75t_L g1202 ( .A(n_1068), .Y(n_1202) );
OAI211xp5_ASAP7_75t_L g1203 ( .A1(n_1035), .A2(n_1042), .B(n_1116), .C(n_1041), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1066), .B(n_1050), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1037), .B(n_1083), .Y(n_1205) );
INVx2_ASAP7_75t_L g1206 ( .A(n_1151), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1113), .B(n_1106), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1132), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1119), .B(n_1107), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1128), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1145), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1212 ( .A(n_1045), .B(n_1033), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1150), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1047), .B(n_1033), .Y(n_1214) );
BUFx2_ASAP7_75t_L g1215 ( .A(n_1131), .Y(n_1215) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_1064), .A2(n_1049), .B1(n_1024), .B2(n_1163), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1101), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1094), .B(n_1100), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1105), .Y(n_1219) );
INVx2_ASAP7_75t_SL g1220 ( .A(n_1063), .Y(n_1220) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_1134), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1122), .Y(n_1222) );
BUFx2_ASAP7_75t_L g1223 ( .A(n_1051), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1065), .B(n_1030), .Y(n_1224) );
OAI31xp33_ASAP7_75t_SL g1225 ( .A1(n_1124), .A2(n_1082), .A3(n_1043), .B(n_1065), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1122), .Y(n_1226) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1155), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1140), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1087), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1104), .Y(n_1230) );
NOR2xp67_ASAP7_75t_L g1231 ( .A(n_1051), .B(n_1154), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1062), .B(n_1070), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1162), .B(n_1073), .Y(n_1233) );
OR2x2_ASAP7_75t_L g1234 ( .A(n_1072), .B(n_1038), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1136), .B(n_1118), .Y(n_1235) );
INVx3_ASAP7_75t_L g1236 ( .A(n_1073), .Y(n_1236) );
AND2x4_ASAP7_75t_L g1237 ( .A(n_1104), .B(n_1125), .Y(n_1237) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1087), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1087), .Y(n_1239) );
BUFx3_ASAP7_75t_L g1240 ( .A(n_1162), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1141), .Y(n_1241) );
HB1xp67_ASAP7_75t_L g1242 ( .A(n_1111), .Y(n_1242) );
INVx2_ASAP7_75t_L g1243 ( .A(n_1104), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1074), .B(n_1078), .Y(n_1244) );
AND2x4_ASAP7_75t_L g1245 ( .A(n_1125), .B(n_1110), .Y(n_1245) );
NAND2x1p5_ASAP7_75t_L g1246 ( .A(n_1111), .B(n_1018), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1121), .B(n_1018), .Y(n_1247) );
INVxp67_ASAP7_75t_SL g1248 ( .A(n_1026), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1022), .B(n_1036), .Y(n_1249) );
BUFx2_ASAP7_75t_L g1250 ( .A(n_1031), .Y(n_1250) );
INVx1_ASAP7_75t_SL g1251 ( .A(n_1114), .Y(n_1251) );
BUFx3_ASAP7_75t_L g1252 ( .A(n_1022), .Y(n_1252) );
INVxp67_ASAP7_75t_L g1253 ( .A(n_1032), .Y(n_1253) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1138), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1056), .B(n_1075), .Y(n_1255) );
INVxp67_ASAP7_75t_L g1256 ( .A(n_1054), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1126), .B(n_1090), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1092), .B(n_1095), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1149), .Y(n_1259) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1139), .Y(n_1260) );
AND2x4_ASAP7_75t_SL g1261 ( .A(n_1057), .B(n_1079), .Y(n_1261) );
BUFx6f_ASAP7_75t_L g1262 ( .A(n_1109), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1023), .B(n_1127), .Y(n_1263) );
BUFx3_ASAP7_75t_L g1264 ( .A(n_1061), .Y(n_1264) );
AOI21xp5_ASAP7_75t_SL g1265 ( .A1(n_1080), .A2(n_1067), .B(n_1130), .Y(n_1265) );
INVx3_ASAP7_75t_L g1266 ( .A(n_1071), .Y(n_1266) );
BUFx2_ASAP7_75t_L g1267 ( .A(n_1152), .Y(n_1267) );
INVx2_ASAP7_75t_SL g1268 ( .A(n_1085), .Y(n_1268) );
HB1xp67_ASAP7_75t_L g1269 ( .A(n_1077), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1060), .B(n_1093), .Y(n_1270) );
INVx3_ASAP7_75t_L g1271 ( .A(n_1017), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1091), .B(n_1146), .Y(n_1272) );
INVx1_ASAP7_75t_SL g1273 ( .A(n_1016), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1089), .B(n_1052), .Y(n_1274) );
INVx3_ASAP7_75t_L g1275 ( .A(n_1069), .Y(n_1275) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1040), .Y(n_1276) );
AND2x4_ASAP7_75t_L g1277 ( .A(n_1046), .B(n_1086), .Y(n_1277) );
AND2x4_ASAP7_75t_L g1278 ( .A(n_1076), .B(n_1084), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1191), .B(n_1053), .Y(n_1279) );
AO21x2_ASAP7_75t_L g1280 ( .A1(n_1231), .A2(n_1229), .B(n_1239), .Y(n_1280) );
OR2x2_ASAP7_75t_L g1281 ( .A(n_1191), .B(n_1193), .Y(n_1281) );
INVx2_ASAP7_75t_L g1282 ( .A(n_1177), .Y(n_1282) );
OAI211xp5_ASAP7_75t_L g1283 ( .A1(n_1171), .A2(n_1253), .B(n_1172), .C(n_1225), .Y(n_1283) );
AOI221xp5_ASAP7_75t_L g1284 ( .A1(n_1207), .A2(n_1172), .B1(n_1211), .B2(n_1183), .C(n_1209), .Y(n_1284) );
HB1xp67_ASAP7_75t_L g1285 ( .A(n_1174), .Y(n_1285) );
AND3x2_ASAP7_75t_L g1286 ( .A(n_1269), .B(n_1223), .C(n_1232), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1197), .Y(n_1287) );
AND2x4_ASAP7_75t_L g1288 ( .A(n_1178), .B(n_1198), .Y(n_1288) );
OAI22xp33_ASAP7_75t_L g1289 ( .A1(n_1275), .A2(n_1223), .B1(n_1249), .B2(n_1196), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1197), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1204), .B(n_1180), .Y(n_1291) );
INVx2_ASAP7_75t_SL g1292 ( .A(n_1189), .Y(n_1292) );
AOI22xp5_ASAP7_75t_L g1293 ( .A1(n_1203), .A2(n_1224), .B1(n_1232), .B2(n_1244), .Y(n_1293) );
INVx2_ASAP7_75t_SL g1294 ( .A(n_1266), .Y(n_1294) );
BUFx3_ASAP7_75t_L g1295 ( .A(n_1240), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1192), .Y(n_1296) );
AOI21xp5_ASAP7_75t_L g1297 ( .A1(n_1265), .A2(n_1231), .B(n_1277), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1204), .B(n_1187), .Y(n_1298) );
INVx5_ASAP7_75t_L g1299 ( .A(n_1266), .Y(n_1299) );
AOI22xp33_ASAP7_75t_SL g1300 ( .A1(n_1275), .A2(n_1224), .B1(n_1214), .B2(n_1244), .Y(n_1300) );
INVxp67_ASAP7_75t_SL g1301 ( .A(n_1199), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1192), .B(n_1187), .Y(n_1302) );
AND2x4_ASAP7_75t_L g1303 ( .A(n_1178), .B(n_1198), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1205), .B(n_1169), .Y(n_1304) );
AOI21xp5_ASAP7_75t_L g1305 ( .A1(n_1265), .A2(n_1277), .B(n_1239), .Y(n_1305) );
HB1xp67_ASAP7_75t_L g1306 ( .A(n_1174), .Y(n_1306) );
NOR2x1_ASAP7_75t_SL g1307 ( .A(n_1200), .B(n_1189), .Y(n_1307) );
AND2x4_ASAP7_75t_L g1308 ( .A(n_1211), .B(n_1200), .Y(n_1308) );
OR2x2_ASAP7_75t_SL g1309 ( .A(n_1202), .B(n_1242), .Y(n_1309) );
AOI22xp5_ASAP7_75t_L g1310 ( .A1(n_1275), .A2(n_1194), .B1(n_1207), .B2(n_1270), .Y(n_1310) );
INVx2_ASAP7_75t_SL g1311 ( .A(n_1266), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1169), .B(n_1210), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1210), .B(n_1184), .Y(n_1313) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1175), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1184), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_1275), .A2(n_1276), .B1(n_1218), .B2(n_1216), .Y(n_1316) );
INVx2_ASAP7_75t_L g1317 ( .A(n_1175), .Y(n_1317) );
INVx4_ASAP7_75t_L g1318 ( .A(n_1189), .Y(n_1318) );
HB1xp67_ASAP7_75t_L g1319 ( .A(n_1199), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1185), .Y(n_1320) );
OR2x2_ASAP7_75t_L g1321 ( .A(n_1190), .B(n_1185), .Y(n_1321) );
INVx2_ASAP7_75t_L g1322 ( .A(n_1170), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1205), .B(n_1240), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1240), .B(n_1221), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1221), .B(n_1246), .Y(n_1325) );
AND2x4_ASAP7_75t_SL g1326 ( .A(n_1266), .B(n_1236), .Y(n_1326) );
INVx1_ASAP7_75t_SL g1327 ( .A(n_1251), .Y(n_1327) );
OAI221xp5_ASAP7_75t_L g1328 ( .A1(n_1234), .A2(n_1212), .B1(n_1233), .B2(n_1276), .C(n_1247), .Y(n_1328) );
AND2x4_ASAP7_75t_L g1329 ( .A(n_1200), .B(n_1170), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1186), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1190), .Y(n_1331) );
INVx2_ASAP7_75t_L g1332 ( .A(n_1181), .Y(n_1332) );
HB1xp67_ASAP7_75t_L g1333 ( .A(n_1213), .Y(n_1333) );
INVx4_ASAP7_75t_L g1334 ( .A(n_1195), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1167), .Y(n_1335) );
INVx3_ASAP7_75t_L g1336 ( .A(n_1195), .Y(n_1336) );
HB1xp67_ASAP7_75t_L g1337 ( .A(n_1213), .Y(n_1337) );
INVx2_ASAP7_75t_SL g1338 ( .A(n_1268), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1167), .B(n_1218), .Y(n_1339) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1176), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1246), .B(n_1195), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1234), .B(n_1212), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1176), .Y(n_1343) );
OAI222xp33_ASAP7_75t_L g1344 ( .A1(n_1200), .A2(n_1188), .B1(n_1214), .B2(n_1220), .C1(n_1168), .C2(n_1263), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1168), .B(n_1220), .Y(n_1345) );
NOR2xp33_ASAP7_75t_L g1346 ( .A(n_1252), .B(n_1256), .Y(n_1346) );
OR2x2_ASAP7_75t_L g1347 ( .A(n_1252), .B(n_1246), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1252), .B(n_1236), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1217), .Y(n_1349) );
AOI211xp5_ASAP7_75t_SL g1350 ( .A1(n_1270), .A2(n_1257), .B(n_1236), .C(n_1248), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1236), .B(n_1235), .Y(n_1351) );
OR2x2_ASAP7_75t_L g1352 ( .A(n_1217), .B(n_1226), .Y(n_1352) );
AOI221x1_ASAP7_75t_L g1353 ( .A1(n_1229), .A2(n_1276), .B1(n_1228), .B2(n_1219), .C(n_1222), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1235), .B(n_1255), .Y(n_1354) );
NAND3xp33_ASAP7_75t_L g1355 ( .A(n_1262), .B(n_1228), .C(n_1257), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1219), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1268), .B(n_1226), .Y(n_1357) );
INVx4_ASAP7_75t_L g1358 ( .A(n_1173), .Y(n_1358) );
OAI221xp5_ASAP7_75t_L g1359 ( .A1(n_1264), .A2(n_1188), .B1(n_1208), .B2(n_1255), .C(n_1200), .Y(n_1359) );
AOI31xp33_ASAP7_75t_L g1360 ( .A1(n_1273), .A2(n_1272), .A3(n_1274), .B(n_1258), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1222), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1362 ( .A(n_1208), .B(n_1182), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1182), .B(n_1237), .Y(n_1363) );
AND2x4_ASAP7_75t_L g1364 ( .A(n_1237), .B(n_1259), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1182), .Y(n_1365) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1182), .Y(n_1366) );
AND2x4_ASAP7_75t_L g1367 ( .A(n_1237), .B(n_1259), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1322), .Y(n_1368) );
AND2x4_ASAP7_75t_SL g1369 ( .A(n_1318), .B(n_1173), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1322), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1287), .B(n_1241), .Y(n_1371) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1354), .B(n_1241), .Y(n_1372) );
NAND5xp2_ASAP7_75t_SL g1373 ( .A(n_1283), .B(n_1272), .C(n_1274), .D(n_1258), .E(n_1261), .Y(n_1373) );
BUFx2_ASAP7_75t_L g1374 ( .A(n_1318), .Y(n_1374) );
NAND3xp33_ASAP7_75t_L g1375 ( .A(n_1316), .B(n_1262), .C(n_1243), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1288), .B(n_1237), .Y(n_1376) );
INVx1_ASAP7_75t_SL g1377 ( .A(n_1327), .Y(n_1377) );
HB1xp67_ASAP7_75t_L g1378 ( .A(n_1285), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1290), .B(n_1230), .Y(n_1379) );
NAND3xp33_ASAP7_75t_L g1380 ( .A(n_1316), .B(n_1262), .C(n_1243), .Y(n_1380) );
OR2x2_ASAP7_75t_L g1381 ( .A(n_1319), .B(n_1230), .Y(n_1381) );
HB1xp67_ASAP7_75t_L g1382 ( .A(n_1285), .Y(n_1382) );
INVx1_ASAP7_75t_SL g1383 ( .A(n_1298), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1288), .B(n_1230), .Y(n_1384) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1340), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1288), .B(n_1245), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1387 ( .A(n_1296), .B(n_1262), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1303), .B(n_1245), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1343), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1303), .B(n_1245), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1303), .B(n_1245), .Y(n_1391) );
BUFx2_ASAP7_75t_L g1392 ( .A(n_1318), .Y(n_1392) );
INVx3_ASAP7_75t_L g1393 ( .A(n_1334), .Y(n_1393) );
NOR2xp33_ASAP7_75t_L g1394 ( .A(n_1338), .B(n_1173), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1364), .B(n_1267), .Y(n_1395) );
INVx1_ASAP7_75t_SL g1396 ( .A(n_1281), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1304), .B(n_1262), .Y(n_1397) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1314), .Y(n_1398) );
HB1xp67_ASAP7_75t_L g1399 ( .A(n_1306), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1364), .B(n_1267), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1364), .B(n_1215), .Y(n_1401) );
BUFx3_ASAP7_75t_L g1402 ( .A(n_1299), .Y(n_1402) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1317), .Y(n_1403) );
AND2x4_ASAP7_75t_L g1404 ( .A(n_1329), .B(n_1271), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1405 ( .A(n_1331), .B(n_1201), .Y(n_1405) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1317), .Y(n_1406) );
NOR2xp33_ASAP7_75t_L g1407 ( .A(n_1291), .B(n_1173), .Y(n_1407) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1282), .Y(n_1408) );
INVxp67_ASAP7_75t_L g1409 ( .A(n_1346), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1367), .B(n_1215), .Y(n_1410) );
BUFx3_ASAP7_75t_L g1411 ( .A(n_1299), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_1367), .B(n_1351), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1315), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1367), .B(n_1260), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1320), .Y(n_1415) );
OR2x2_ASAP7_75t_L g1416 ( .A(n_1319), .B(n_1301), .Y(n_1416) );
OR2x2_ASAP7_75t_L g1417 ( .A(n_1301), .B(n_1227), .Y(n_1417) );
HB1xp67_ASAP7_75t_L g1418 ( .A(n_1306), .Y(n_1418) );
OR2x2_ASAP7_75t_L g1419 ( .A(n_1342), .B(n_1227), .Y(n_1419) );
OR2x2_ASAP7_75t_L g1420 ( .A(n_1321), .B(n_1227), .Y(n_1420) );
OR2x2_ASAP7_75t_L g1421 ( .A(n_1302), .B(n_1260), .Y(n_1421) );
NOR2xp67_ASAP7_75t_L g1422 ( .A(n_1334), .B(n_1238), .Y(n_1422) );
INVx2_ASAP7_75t_L g1423 ( .A(n_1332), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1363), .B(n_1254), .Y(n_1424) );
INVx2_ASAP7_75t_L g1425 ( .A(n_1332), .Y(n_1425) );
OR2x2_ASAP7_75t_L g1426 ( .A(n_1339), .B(n_1254), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1308), .B(n_1254), .Y(n_1427) );
OR2x2_ASAP7_75t_L g1428 ( .A(n_1333), .B(n_1206), .Y(n_1428) );
INVx2_ASAP7_75t_SL g1429 ( .A(n_1334), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1430 ( .A(n_1330), .B(n_1201), .Y(n_1430) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1383), .B(n_1284), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_1424), .B(n_1308), .Y(n_1432) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1385), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1396), .B(n_1335), .Y(n_1434) );
HB1xp67_ASAP7_75t_L g1435 ( .A(n_1416), .Y(n_1435) );
NOR2xp33_ASAP7_75t_L g1436 ( .A(n_1409), .B(n_1360), .Y(n_1436) );
NOR2xp33_ASAP7_75t_L g1437 ( .A(n_1377), .B(n_1310), .Y(n_1437) );
NAND2xp5_ASAP7_75t_L g1438 ( .A(n_1372), .B(n_1293), .Y(n_1438) );
AOI21xp33_ASAP7_75t_L g1439 ( .A1(n_1394), .A2(n_1289), .B(n_1359), .Y(n_1439) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1385), .Y(n_1440) );
NAND2xp5_ASAP7_75t_L g1441 ( .A(n_1372), .B(n_1312), .Y(n_1441) );
BUFx2_ASAP7_75t_L g1442 ( .A(n_1374), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1424), .B(n_1414), .Y(n_1443) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_1397), .B(n_1309), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1389), .Y(n_1445) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1413), .Y(n_1446) );
AND2x4_ASAP7_75t_L g1447 ( .A(n_1404), .B(n_1329), .Y(n_1447) );
OR2x2_ASAP7_75t_L g1448 ( .A(n_1421), .B(n_1333), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1413), .Y(n_1449) );
OR2x6_ASAP7_75t_L g1450 ( .A(n_1374), .B(n_1392), .Y(n_1450) );
HB1xp67_ASAP7_75t_L g1451 ( .A(n_1416), .Y(n_1451) );
INVx2_ASAP7_75t_L g1452 ( .A(n_1423), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1414), .B(n_1308), .Y(n_1453) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1415), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_1421), .B(n_1313), .Y(n_1455) );
INVx2_ASAP7_75t_L g1456 ( .A(n_1423), .Y(n_1456) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1415), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1412), .B(n_1329), .Y(n_1458) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1378), .Y(n_1459) );
NOR2x1_ASAP7_75t_L g1460 ( .A(n_1402), .B(n_1358), .Y(n_1460) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1382), .Y(n_1461) );
NAND2x1_ASAP7_75t_L g1462 ( .A(n_1392), .B(n_1358), .Y(n_1462) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1425), .Y(n_1463) );
NOR3xp33_ASAP7_75t_SL g1464 ( .A(n_1380), .B(n_1289), .C(n_1344), .Y(n_1464) );
AND2x4_ASAP7_75t_L g1465 ( .A(n_1404), .B(n_1307), .Y(n_1465) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1399), .Y(n_1466) );
OR2x2_ASAP7_75t_L g1467 ( .A(n_1420), .B(n_1337), .Y(n_1467) );
OR2x2_ASAP7_75t_L g1468 ( .A(n_1420), .B(n_1337), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1412), .B(n_1323), .Y(n_1469) );
OAI21xp5_ASAP7_75t_L g1470 ( .A1(n_1429), .A2(n_1350), .B(n_1297), .Y(n_1470) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1418), .Y(n_1471) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1368), .Y(n_1472) );
INVxp67_ASAP7_75t_L g1473 ( .A(n_1407), .Y(n_1473) );
AND2x4_ASAP7_75t_L g1474 ( .A(n_1404), .B(n_1355), .Y(n_1474) );
OR2x2_ASAP7_75t_L g1475 ( .A(n_1419), .B(n_1362), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1386), .B(n_1280), .Y(n_1476) );
INVx1_ASAP7_75t_SL g1477 ( .A(n_1369), .Y(n_1477) );
HB1xp67_ASAP7_75t_L g1478 ( .A(n_1428), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1368), .Y(n_1479) );
O2A1O1Ixp33_ASAP7_75t_L g1480 ( .A1(n_1437), .A2(n_1373), .B(n_1346), .C(n_1311), .Y(n_1480) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1478), .Y(n_1481) );
AND2x4_ASAP7_75t_L g1482 ( .A(n_1450), .B(n_1404), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1443), .B(n_1427), .Y(n_1483) );
INVx2_ASAP7_75t_L g1484 ( .A(n_1452), .Y(n_1484) );
NAND2xp5_ASAP7_75t_L g1485 ( .A(n_1435), .B(n_1426), .Y(n_1485) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1478), .Y(n_1486) );
NOR2xp33_ASAP7_75t_SL g1487 ( .A(n_1477), .B(n_1373), .Y(n_1487) );
INVx2_ASAP7_75t_L g1488 ( .A(n_1452), .Y(n_1488) );
INVx1_ASAP7_75t_SL g1489 ( .A(n_1442), .Y(n_1489) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1435), .Y(n_1490) );
OAI21xp5_ASAP7_75t_L g1491 ( .A1(n_1464), .A2(n_1300), .B(n_1429), .Y(n_1491) );
AOI211xp5_ASAP7_75t_L g1492 ( .A1(n_1439), .A2(n_1328), .B(n_1380), .C(n_1375), .Y(n_1492) );
CKINVDCx16_ASAP7_75t_R g1493 ( .A(n_1450), .Y(n_1493) );
AOI22xp5_ASAP7_75t_L g1494 ( .A1(n_1436), .A2(n_1300), .B1(n_1286), .B2(n_1401), .Y(n_1494) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1451), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g1496 ( .A(n_1451), .B(n_1426), .Y(n_1496) );
OAI31xp33_ASAP7_75t_L g1497 ( .A1(n_1436), .A2(n_1369), .A3(n_1393), .B(n_1326), .Y(n_1497) );
NAND2xp5_ASAP7_75t_L g1498 ( .A(n_1438), .B(n_1371), .Y(n_1498) );
AOI22xp33_ASAP7_75t_L g1499 ( .A1(n_1437), .A2(n_1395), .B1(n_1400), .B2(n_1401), .Y(n_1499) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_1443), .B(n_1427), .Y(n_1500) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1448), .B(n_1419), .Y(n_1501) );
INVx1_ASAP7_75t_SL g1502 ( .A(n_1469), .Y(n_1502) );
AOI21xp5_ASAP7_75t_L g1503 ( .A1(n_1462), .A2(n_1422), .B(n_1393), .Y(n_1503) );
AOI221xp5_ASAP7_75t_L g1504 ( .A1(n_1431), .A2(n_1357), .B1(n_1430), .B2(n_1400), .C(n_1395), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1476), .B(n_1410), .Y(n_1505) );
AOI21xp5_ASAP7_75t_L g1506 ( .A1(n_1470), .A2(n_1422), .B(n_1393), .Y(n_1506) );
OR2x2_ASAP7_75t_L g1507 ( .A(n_1467), .B(n_1381), .Y(n_1507) );
AOI22xp33_ASAP7_75t_SL g1508 ( .A1(n_1465), .A2(n_1402), .B1(n_1411), .B2(n_1376), .Y(n_1508) );
AOI22xp5_ASAP7_75t_L g1509 ( .A1(n_1473), .A2(n_1286), .B1(n_1410), .B2(n_1386), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1476), .B(n_1388), .Y(n_1510) );
INVx2_ASAP7_75t_L g1511 ( .A(n_1456), .Y(n_1511) );
AOI21xp5_ASAP7_75t_L g1512 ( .A1(n_1450), .A2(n_1292), .B(n_1358), .Y(n_1512) );
BUFx2_ASAP7_75t_L g1513 ( .A(n_1460), .Y(n_1513) );
NAND2xp5_ASAP7_75t_L g1514 ( .A(n_1490), .B(n_1459), .Y(n_1514) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1485), .Y(n_1515) );
NAND2xp5_ASAP7_75t_L g1516 ( .A(n_1490), .B(n_1461), .Y(n_1516) );
NOR2xp33_ASAP7_75t_L g1517 ( .A(n_1498), .B(n_1444), .Y(n_1517) );
HB1xp67_ASAP7_75t_L g1518 ( .A(n_1495), .Y(n_1518) );
NAND2xp5_ASAP7_75t_L g1519 ( .A(n_1495), .B(n_1466), .Y(n_1519) );
NAND2xp5_ASAP7_75t_L g1520 ( .A(n_1481), .B(n_1471), .Y(n_1520) );
AOI222xp33_ASAP7_75t_L g1521 ( .A1(n_1491), .A2(n_1441), .B1(n_1455), .B2(n_1434), .C1(n_1474), .C2(n_1440), .Y(n_1521) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1496), .Y(n_1522) );
INVx2_ASAP7_75t_L g1523 ( .A(n_1484), .Y(n_1523) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1507), .Y(n_1524) );
INVx2_ASAP7_75t_L g1525 ( .A(n_1484), .Y(n_1525) );
O2A1O1Ixp33_ASAP7_75t_L g1526 ( .A1(n_1487), .A2(n_1464), .B(n_1294), .C(n_1345), .Y(n_1526) );
XNOR2x1_ASAP7_75t_L g1527 ( .A(n_1502), .B(n_1475), .Y(n_1527) );
AOI322xp5_ASAP7_75t_L g1528 ( .A1(n_1493), .A2(n_1458), .A3(n_1432), .B1(n_1453), .B2(n_1376), .C1(n_1388), .C2(n_1390), .Y(n_1528) );
AOI221xp5_ASAP7_75t_L g1529 ( .A1(n_1504), .A2(n_1432), .B1(n_1449), .B2(n_1433), .C(n_1445), .Y(n_1529) );
OR2x2_ASAP7_75t_L g1530 ( .A(n_1507), .B(n_1468), .Y(n_1530) );
NAND2xp5_ASAP7_75t_SL g1531 ( .A(n_1513), .B(n_1465), .Y(n_1531) );
AOI22xp5_ASAP7_75t_L g1532 ( .A1(n_1494), .A2(n_1447), .B1(n_1453), .B2(n_1458), .Y(n_1532) );
NOR2x1_ASAP7_75t_L g1533 ( .A(n_1513), .B(n_1411), .Y(n_1533) );
OR2x2_ASAP7_75t_L g1534 ( .A(n_1501), .B(n_1417), .Y(n_1534) );
AOI21xp33_ASAP7_75t_L g1535 ( .A1(n_1480), .A2(n_1405), .B(n_1474), .Y(n_1535) );
O2A1O1Ixp5_ASAP7_75t_L g1536 ( .A1(n_1503), .A2(n_1465), .B(n_1474), .C(n_1446), .Y(n_1536) );
AOI211xp5_ASAP7_75t_L g1537 ( .A1(n_1526), .A2(n_1497), .B(n_1506), .C(n_1512), .Y(n_1537) );
NAND2xp5_ASAP7_75t_L g1538 ( .A(n_1529), .B(n_1492), .Y(n_1538) );
A2O1A1Ixp33_ASAP7_75t_L g1539 ( .A1(n_1536), .A2(n_1508), .B(n_1482), .C(n_1509), .Y(n_1539) );
AOI322xp5_ASAP7_75t_L g1540 ( .A1(n_1532), .A2(n_1499), .A3(n_1505), .B1(n_1483), .B2(n_1500), .C1(n_1510), .C2(n_1489), .Y(n_1540) );
AOI22xp5_ASAP7_75t_L g1541 ( .A1(n_1521), .A2(n_1482), .B1(n_1486), .B2(n_1510), .Y(n_1541) );
NOR2xp67_ASAP7_75t_L g1542 ( .A(n_1531), .B(n_1482), .Y(n_1542) );
INVx2_ASAP7_75t_SL g1543 ( .A(n_1527), .Y(n_1543) );
AOI22xp5_ASAP7_75t_L g1544 ( .A1(n_1517), .A2(n_1486), .B1(n_1505), .B2(n_1447), .Y(n_1544) );
INVx2_ASAP7_75t_L g1545 ( .A(n_1523), .Y(n_1545) );
AOI211xp5_ASAP7_75t_L g1546 ( .A1(n_1526), .A2(n_1341), .B(n_1325), .C(n_1347), .Y(n_1546) );
AOI221xp5_ASAP7_75t_L g1547 ( .A1(n_1517), .A2(n_1500), .B1(n_1483), .B2(n_1457), .C(n_1454), .Y(n_1547) );
AOI22xp33_ASAP7_75t_L g1548 ( .A1(n_1535), .A2(n_1447), .B1(n_1390), .B2(n_1391), .Y(n_1548) );
OA21x2_ASAP7_75t_L g1549 ( .A1(n_1536), .A2(n_1353), .B(n_1511), .Y(n_1549) );
INVx2_ASAP7_75t_L g1550 ( .A(n_1525), .Y(n_1550) );
OAI22xp33_ASAP7_75t_L g1551 ( .A1(n_1533), .A2(n_1299), .B1(n_1292), .B2(n_1295), .Y(n_1551) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1514), .Y(n_1552) );
AOI22xp5_ASAP7_75t_L g1553 ( .A1(n_1543), .A2(n_1522), .B1(n_1515), .B2(n_1524), .Y(n_1553) );
INVx1_ASAP7_75t_SL g1554 ( .A(n_1552), .Y(n_1554) );
NAND4xp25_ASAP7_75t_L g1555 ( .A(n_1539), .B(n_1528), .C(n_1305), .D(n_1279), .Y(n_1555) );
OAI222xp33_ASAP7_75t_L g1556 ( .A1(n_1541), .A2(n_1530), .B1(n_1534), .B2(n_1520), .C1(n_1519), .C2(n_1516), .Y(n_1556) );
AOI221xp5_ASAP7_75t_L g1557 ( .A1(n_1538), .A2(n_1547), .B1(n_1548), .B2(n_1537), .C(n_1546), .Y(n_1557) );
AOI22xp5_ASAP7_75t_L g1558 ( .A1(n_1537), .A2(n_1518), .B1(n_1391), .B2(n_1384), .Y(n_1558) );
AND2x2_ASAP7_75t_L g1559 ( .A(n_1542), .B(n_1518), .Y(n_1559) );
AOI321xp33_ASAP7_75t_L g1560 ( .A1(n_1546), .A2(n_1324), .A3(n_1387), .B1(n_1366), .B2(n_1365), .C(n_1384), .Y(n_1560) );
INVx1_ASAP7_75t_SL g1561 ( .A(n_1545), .Y(n_1561) );
AOI222xp33_ASAP7_75t_L g1562 ( .A1(n_1551), .A2(n_1511), .B1(n_1488), .B2(n_1479), .C1(n_1472), .C2(n_1299), .Y(n_1562) );
AOI221xp5_ASAP7_75t_L g1563 ( .A1(n_1544), .A2(n_1488), .B1(n_1379), .B2(n_1349), .C(n_1356), .Y(n_1563) );
AND2x4_ASAP7_75t_L g1564 ( .A(n_1554), .B(n_1550), .Y(n_1564) );
OR5x1_ASAP7_75t_L g1565 ( .A(n_1555), .B(n_1540), .C(n_1549), .D(n_1326), .E(n_1295), .Y(n_1565) );
OAI311xp33_ASAP7_75t_L g1566 ( .A1(n_1557), .A2(n_1549), .A3(n_1352), .B1(n_1336), .C1(n_1428), .Y(n_1566) );
AND2x4_ASAP7_75t_L g1567 ( .A(n_1553), .B(n_1463), .Y(n_1567) );
HB1xp67_ASAP7_75t_L g1568 ( .A(n_1561), .Y(n_1568) );
AOI22xp5_ASAP7_75t_L g1569 ( .A1(n_1558), .A2(n_1261), .B1(n_1348), .B2(n_1264), .Y(n_1569) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1563), .B(n_1456), .Y(n_1570) );
OR4x2_ASAP7_75t_L g1571 ( .A(n_1565), .B(n_1556), .C(n_1560), .D(n_1559), .Y(n_1571) );
AND4x1_ASAP7_75t_L g1572 ( .A(n_1569), .B(n_1562), .C(n_1560), .D(n_1361), .Y(n_1572) );
OA22x2_ASAP7_75t_L g1573 ( .A1(n_1568), .A2(n_1261), .B1(n_1336), .B2(n_1370), .Y(n_1573) );
NOR3xp33_ASAP7_75t_L g1574 ( .A(n_1564), .B(n_1179), .C(n_1264), .Y(n_1574) );
OAI22x1_ASAP7_75t_L g1575 ( .A1(n_1572), .A2(n_1567), .B1(n_1566), .B2(n_1570), .Y(n_1575) );
OR2x6_ASAP7_75t_L g1576 ( .A(n_1573), .B(n_1567), .Y(n_1576) );
OAI22xp5_ASAP7_75t_SL g1577 ( .A1(n_1575), .A2(n_1571), .B1(n_1576), .B2(n_1574), .Y(n_1577) );
OAI22xp5_ASAP7_75t_SL g1578 ( .A1(n_1576), .A2(n_1250), .B1(n_1278), .B2(n_1277), .Y(n_1578) );
OAI22xp5_ASAP7_75t_L g1579 ( .A1(n_1577), .A2(n_1398), .B1(n_1403), .B2(n_1406), .Y(n_1579) );
OAI222xp33_ASAP7_75t_L g1580 ( .A1(n_1579), .A2(n_1578), .B1(n_1278), .B2(n_1179), .C1(n_1277), .C2(n_1271), .Y(n_1580) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1580), .Y(n_1581) );
OAI22xp33_ASAP7_75t_L g1582 ( .A1(n_1581), .A2(n_1398), .B1(n_1406), .B2(n_1408), .Y(n_1582) );
endmodule