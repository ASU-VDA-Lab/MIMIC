module real_jpeg_11771_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_276, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_276;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx2_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_6),
.A2(n_32),
.B1(n_34),
.B2(n_58),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_58),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_6),
.A2(n_58),
.B1(n_64),
.B2(n_67),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_7),
.A2(n_32),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_7),
.A2(n_42),
.B1(n_64),
.B2(n_67),
.Y(n_209)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_63),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_10),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_102),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_10),
.A2(n_64),
.B1(n_67),
.B2(n_102),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_10),
.A2(n_32),
.B1(n_34),
.B2(n_102),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_12),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_12),
.A2(n_64),
.B1(n_67),
.B2(n_83),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_12),
.A2(n_32),
.B1(n_34),
.B2(n_83),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_13),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_13),
.B(n_64),
.C(n_79),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_13),
.B(n_35),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_68),
.B(n_156),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_13),
.A2(n_31),
.B(n_34),
.C(n_183),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_13),
.A2(n_32),
.B1(n_34),
.B2(n_141),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_13),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_13),
.B(n_45),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_14),
.A2(n_49),
.B1(n_64),
.B2(n_67),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_49),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_14),
.A2(n_32),
.B1(n_34),
.B2(n_49),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_64),
.B1(n_67),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_15),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_72),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_16),
.A2(n_32),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_16),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_16),
.A2(n_39),
.B1(n_64),
.B2(n_67),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_129),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_106),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_21),
.B(n_106),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_86),
.C(n_94),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_22),
.A2(n_23),
.B1(n_86),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_59),
.B2(n_85),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_26),
.B(n_43),
.C(n_85),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_27),
.A2(n_40),
.B1(n_41),
.B2(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_27),
.A2(n_188),
.B(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_27),
.A2(n_40),
.B1(n_202),
.B2(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_27),
.A2(n_189),
.B(n_229),
.Y(n_249)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_28),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_29)
);

AO22x1_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_30),
.A2(n_36),
.B(n_141),
.Y(n_183)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_34),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g238 ( 
.A(n_32),
.B(n_52),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI32xp33_ASAP7_75t_L g237 ( 
.A1(n_34),
.A2(n_46),
.A3(n_53),
.B1(n_226),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_35),
.B(n_105),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_36),
.A2(n_37),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_37),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_38),
.A2(n_40),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_40),
.A2(n_104),
.B(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_50),
.B(n_55),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_44),
.A2(n_50),
.B1(n_51),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_46),
.B1(n_52),
.B2(n_53),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_46),
.A2(n_50),
.B(n_141),
.C(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_51),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_51),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_51),
.A2(n_101),
.B(n_123),
.Y(n_250)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_56),
.B(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_74),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_60),
.A2(n_74),
.B1(n_75),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_60),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_68),
.B1(n_71),
.B2(n_73),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_69),
.B1(n_70),
.B2(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_67),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_67),
.B(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_68),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_68),
.A2(n_73),
.B1(n_185),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_68),
.A2(n_73),
.B1(n_209),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_70),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_69),
.A2(n_70),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_69),
.B(n_157),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_70),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_70),
.B(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_73),
.A2(n_162),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_73),
.B(n_141),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_73),
.A2(n_170),
.B(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_82),
.B2(n_84),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_77),
.B1(n_84),
.B2(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_82),
.B1(n_84),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_77),
.B(n_143),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_77),
.A2(n_84),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_92),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_81),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_81),
.B(n_141),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_81),
.A2(n_153),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_84),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_86),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_93),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_88),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_93),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_90),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_94),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.C(n_103),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_95),
.B(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_96),
.B(n_98),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_97),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_99),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_100),
.B(n_103),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_128),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_116),
.B2(n_117),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B(n_115),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_113),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_140),
.B(n_142),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_111),
.A2(n_142),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_126),
.B2(n_127),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_269),
.B(n_274),
.Y(n_130)
);

OAI321xp33_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_243),
.A3(n_262),
.B1(n_267),
.B2(n_268),
.C(n_276),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_218),
.B(n_242),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_196),
.B(n_217),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_178),
.B(n_195),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_158),
.B(n_177),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_146),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_139),
.B1(n_144),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_151),
.C(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_155),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_166),
.B(n_176),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_164),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_171),
.B(n_175),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_168),
.B(n_169),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_180),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_186),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_190),
.C(n_194),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_184),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_186)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_192),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_197),
.B(n_198),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_210),
.B2(n_211),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_213),
.C(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_204),
.C(n_208),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_219),
.B(n_220),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_233),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_234),
.C(n_235),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_227),
.B2(n_232),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_228),
.C(n_230),
.Y(n_254)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_227),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_255),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_255),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_253),
.C(n_254),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_245),
.A2(n_246),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_252),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_251),
.C(n_252),
.Y(n_261)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_253),
.B(n_254),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_261),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_259),
.C(n_261),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_263),
.B(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_273),
.Y(n_274)
);


endmodule