module fake_netlist_6_979_n_772 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_772);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_772;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_544;
wire n_468;
wire n_372;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_30),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_15),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_145),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_85),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_64),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_116),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_32),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_25),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_96),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_4),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_128),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_44),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_69),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_100),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_2),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_4),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_87),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_99),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_131),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_20),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_136),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_31),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_36),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_46),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_140),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_26),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_66),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_76),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_79),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_52),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_55),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_34),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_39),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_57),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_86),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_113),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_141),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_7),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_21),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_15),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_139),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_1),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_16),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_0),
.Y(n_199)
);

BUFx8_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_149),
.B(n_0),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_150),
.B(n_1),
.Y(n_208)
);

BUFx8_ASAP7_75t_SL g209 ( 
.A(n_193),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_23),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_148),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_24),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_165),
.B(n_2),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_168),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_146),
.Y(n_223)
);

BUFx8_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

BUFx8_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_152),
.B(n_27),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_153),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_151),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_147),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_147),
.B(n_3),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_154),
.B(n_3),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_220),
.B1(n_208),
.B2(n_199),
.Y(n_239)
);

AO22x2_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_167),
.B1(n_6),
.B2(n_7),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_217),
.B(n_192),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_236),
.A2(n_162),
.B1(n_172),
.B2(n_196),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_196),
.B1(n_191),
.B2(n_190),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

AO22x2_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_186),
.B1(n_183),
.B2(n_182),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_156),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_211),
.A2(n_181),
.B1(n_180),
.B2(n_179),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_211),
.A2(n_169),
.B1(n_175),
.B2(n_174),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_217),
.B(n_157),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_209),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_211),
.A2(n_166),
.B1(n_173),
.B2(n_171),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_158),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_178),
.B1(n_170),
.B2(n_164),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_234),
.A2(n_204),
.B1(n_206),
.B2(n_237),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_161),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_234),
.A2(n_163),
.B1(n_8),
.B2(n_9),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_214),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_265)
);

AO22x2_ASAP7_75t_L g266 ( 
.A1(n_232),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_202),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_268)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_28),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_203),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_223),
.B(n_29),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_223),
.B(n_237),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_202),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_275)
);

AO22x2_ASAP7_75t_L g276 ( 
.A1(n_202),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_213),
.Y(n_277)
);

AO22x2_ASAP7_75t_L g278 ( 
.A1(n_212),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_212),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_279)
);

AO22x2_ASAP7_75t_L g280 ( 
.A1(n_212),
.A2(n_22),
.B1(n_33),
.B2(n_35),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_223),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_213),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_237),
.B(n_40),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_215),
.B(n_41),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_215),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_255),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_245),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_248),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_227),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_227),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_233),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_241),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_269),
.B(n_209),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_260),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_230),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_243),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_247),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_239),
.B(n_230),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_269),
.B(n_200),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_257),
.B(n_233),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_276),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_273),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_280),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_269),
.B(n_231),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_274),
.B(n_231),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_250),
.B(n_231),
.Y(n_322)
);

NAND2xp33_ASAP7_75t_R g323 ( 
.A(n_240),
.B(n_47),
.Y(n_323)
);

NAND2x1p5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_210),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_281),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_285),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_252),
.B(n_233),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_249),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_266),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_240),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_252),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_253),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_253),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_256),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_256),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_250),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_244),
.B(n_200),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_242),
.B(n_222),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_254),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_264),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_268),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_264),
.B(n_48),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_258),
.Y(n_347)
);

NAND2xp33_ASAP7_75t_SL g348 ( 
.A(n_265),
.B(n_222),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_233),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_219),
.Y(n_350)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_320),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_320),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_287),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_289),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_322),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_287),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_233),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_305),
.B(n_219),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_299),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_305),
.B(n_219),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_337),
.B(n_275),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_292),
.B(n_219),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_292),
.B(n_219),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_322),
.Y(n_364)
);

AND2x6_ASAP7_75t_L g365 ( 
.A(n_326),
.B(n_320),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_300),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_312),
.B(n_226),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_289),
.B(n_226),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_303),
.Y(n_370)
);

INVx8_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_304),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_306),
.Y(n_373)
);

AND2x2_ASAP7_75t_SL g374 ( 
.A(n_307),
.B(n_226),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_226),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_311),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_288),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_342),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_290),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_310),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_291),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_318),
.B(n_226),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_319),
.B(n_228),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_228),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_298),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_310),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_308),
.B(n_228),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_327),
.B(n_228),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_338),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_343),
.B(n_228),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_332),
.B(n_330),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_316),
.A2(n_218),
.B(n_221),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_347),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_317),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_293),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_347),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_339),
.A2(n_218),
.B(n_221),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_347),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_R g407 ( 
.A(n_286),
.B(n_49),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_345),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_309),
.B(n_218),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_309),
.B(n_218),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_294),
.Y(n_413)
);

INVxp33_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_294),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_331),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_369),
.B(n_325),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_354),
.B(n_392),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_351),
.B(n_329),
.Y(n_420)
);

BUFx8_ASAP7_75t_SL g421 ( 
.A(n_408),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_355),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_351),
.B(n_333),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_351),
.B(n_344),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_416),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_399),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_358),
.B(n_295),
.Y(n_428)
);

CKINVDCx6p67_ASAP7_75t_R g429 ( 
.A(n_415),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_364),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_406),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_353),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_358),
.B(n_341),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_360),
.B(n_346),
.Y(n_435)
);

NAND2x1p5_ASAP7_75t_L g436 ( 
.A(n_351),
.B(n_205),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_387),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_360),
.B(n_336),
.Y(n_439)
);

NAND2x1p5_ASAP7_75t_L g440 ( 
.A(n_352),
.B(n_205),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_369),
.B(n_336),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_375),
.B(n_224),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_301),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_375),
.B(n_224),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_387),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_387),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_406),
.B(n_323),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_406),
.B(n_210),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_352),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_400),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_356),
.Y(n_451)
);

OR2x6_ASAP7_75t_L g452 ( 
.A(n_371),
.B(n_265),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_50),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_350),
.B(n_224),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_352),
.B(n_301),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_350),
.B(n_225),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_387),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_387),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_400),
.B(n_403),
.Y(n_459)
);

BUFx12f_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_416),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_403),
.B(n_225),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_405),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_408),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_415),
.B(n_286),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_356),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_371),
.B(n_296),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_371),
.B(n_296),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_406),
.B(n_323),
.Y(n_470)
);

NAND2x1p5_ASAP7_75t_L g471 ( 
.A(n_352),
.B(n_406),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_384),
.B(n_225),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_418),
.B(n_405),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_432),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_447),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_447),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_438),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_439),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_447),
.A2(n_371),
.B1(n_405),
.B2(n_378),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_438),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_438),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_425),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_445),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_439),
.Y(n_485)
);

INVx6_ASAP7_75t_L g486 ( 
.A(n_445),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_432),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_425),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_447),
.A2(n_371),
.B1(n_405),
.B2(n_378),
.Y(n_489)
);

BUFx4f_ASAP7_75t_L g490 ( 
.A(n_447),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_445),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_429),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_470),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_435),
.B(n_384),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_470),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_445),
.Y(n_496)
);

INVx3_ASAP7_75t_SL g497 ( 
.A(n_429),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_421),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_435),
.B(n_414),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_421),
.Y(n_500)
);

BUFx2_ASAP7_75t_SL g501 ( 
.A(n_446),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_433),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_424),
.B(n_464),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_433),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_446),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_441),
.A2(n_361),
.B1(n_396),
.B2(n_392),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_470),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_460),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_441),
.B(n_397),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_470),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_425),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_426),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_470),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_451),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_450),
.B(n_388),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_428),
.A2(n_402),
.B1(n_397),
.B2(n_406),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_446),
.Y(n_517)
);

BUFx24_ASAP7_75t_L g518 ( 
.A(n_455),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_426),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_449),
.B(n_409),
.Y(n_520)
);

INVx6_ASAP7_75t_L g521 ( 
.A(n_446),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_516),
.A2(n_409),
.B1(n_452),
.B2(n_374),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_473),
.A2(n_357),
.B(n_459),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_487),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_478),
.A2(n_443),
.B1(n_452),
.B2(n_434),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g526 ( 
.A1(n_506),
.A2(n_468),
.B1(n_467),
.B2(n_465),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_494),
.A2(n_443),
.B1(n_428),
.B2(n_434),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_487),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_498),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_508),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_497),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_502),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_478),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_485),
.A2(n_452),
.B1(n_455),
.B2(n_422),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_490),
.A2(n_409),
.B1(n_452),
.B2(n_494),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_502),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_SL g537 ( 
.A1(n_506),
.A2(n_485),
.B1(n_499),
.B2(n_407),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_497),
.Y(n_538)
);

INVx6_ASAP7_75t_L g539 ( 
.A(n_499),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_491),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_509),
.A2(n_455),
.B1(n_430),
.B2(n_359),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_509),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_474),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_483),
.A2(n_359),
.B1(n_402),
.B2(n_419),
.Y(n_544)
);

INVx6_ASAP7_75t_L g545 ( 
.A(n_491),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_483),
.A2(n_419),
.B1(n_348),
.B2(n_388),
.Y(n_546)
);

NAND2x1p5_ASAP7_75t_L g547 ( 
.A(n_491),
.B(n_449),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_488),
.A2(n_348),
.B1(n_469),
.B2(n_461),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_504),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_504),
.Y(n_550)
);

BUFx8_ASAP7_75t_L g551 ( 
.A(n_512),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_505),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_479),
.Y(n_553)
);

OAI22xp33_ASAP7_75t_L g554 ( 
.A1(n_497),
.A2(n_460),
.B1(n_409),
.B2(n_472),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_488),
.A2(n_469),
.B1(n_461),
.B2(n_409),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_474),
.Y(n_556)
);

BUFx12f_ASAP7_75t_L g557 ( 
.A(n_512),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_504),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_492),
.A2(n_409),
.B1(n_442),
.B2(n_444),
.Y(n_559)
);

INVx6_ASAP7_75t_L g560 ( 
.A(n_486),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_518),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_514),
.Y(n_562)
);

CKINVDCx11_ASAP7_75t_R g563 ( 
.A(n_500),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_490),
.A2(n_374),
.B1(n_431),
.B2(n_401),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_511),
.A2(n_417),
.B1(n_427),
.B2(n_374),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_549),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_551),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_526),
.A2(n_349),
.B1(n_454),
.B2(n_456),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_539),
.A2(n_462),
.B1(n_362),
.B2(n_363),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_542),
.B(n_514),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_542),
.B(n_475),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_533),
.B(n_515),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_540),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_527),
.B(n_503),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_535),
.B(n_390),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_524),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_551),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_528),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_539),
.A2(n_537),
.B1(n_525),
.B2(n_535),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_550),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_534),
.A2(n_362),
.B1(n_363),
.B2(n_453),
.Y(n_581)
);

OAI222xp33_ASAP7_75t_L g582 ( 
.A1(n_522),
.A2(n_511),
.B1(n_480),
.B2(n_489),
.C1(n_513),
.C2(n_495),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_541),
.A2(n_490),
.B1(n_394),
.B2(n_510),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_546),
.A2(n_490),
.B1(n_475),
.B2(n_476),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_548),
.A2(n_495),
.B1(n_476),
.B2(n_493),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_532),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_522),
.A2(n_394),
.B1(n_493),
.B2(n_507),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_L g588 ( 
.A1(n_561),
.A2(n_476),
.B1(n_475),
.B2(n_495),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_559),
.A2(n_510),
.B1(n_493),
.B2(n_507),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_SL g590 ( 
.A1(n_561),
.A2(n_513),
.B1(n_507),
.B2(n_510),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_564),
.A2(n_513),
.B1(n_404),
.B2(n_501),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_563),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_536),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_544),
.B(n_519),
.Y(n_594)
);

BUFx4f_ASAP7_75t_SL g595 ( 
.A(n_557),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_SL g596 ( 
.A1(n_564),
.A2(n_538),
.B1(n_531),
.B2(n_529),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_565),
.A2(n_386),
.B1(n_379),
.B2(n_385),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_554),
.A2(n_420),
.B1(n_423),
.B2(n_519),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_543),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_555),
.A2(n_420),
.B1(n_520),
.B2(n_471),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_523),
.A2(n_379),
.B1(n_386),
.B2(n_377),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_556),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_523),
.A2(n_377),
.B1(n_385),
.B2(n_373),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_562),
.A2(n_377),
.B1(n_385),
.B2(n_373),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_552),
.A2(n_404),
.B(n_420),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_558),
.Y(n_606)
);

CKINVDCx11_ASAP7_75t_R g607 ( 
.A(n_553),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_560),
.A2(n_372),
.B1(n_381),
.B2(n_367),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_560),
.A2(n_372),
.B1(n_381),
.B2(n_383),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_552),
.A2(n_381),
.B1(n_383),
.B2(n_368),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_530),
.A2(n_381),
.B1(n_368),
.B2(n_370),
.Y(n_611)
);

CKINVDCx11_ASAP7_75t_R g612 ( 
.A(n_553),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_553),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_545),
.A2(n_368),
.B1(n_370),
.B2(n_463),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_574),
.A2(n_579),
.B1(n_568),
.B2(n_596),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_590),
.A2(n_401),
.B1(n_520),
.B2(n_391),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_584),
.A2(n_545),
.B1(n_520),
.B2(n_501),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_588),
.B(n_591),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_589),
.A2(n_391),
.B1(n_393),
.B2(n_395),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_583),
.A2(n_370),
.B1(n_382),
.B2(n_376),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_569),
.A2(n_571),
.B1(n_587),
.B2(n_581),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_598),
.A2(n_395),
.B1(n_391),
.B2(n_393),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_602),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_571),
.A2(n_585),
.B1(n_597),
.B2(n_594),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_575),
.A2(n_376),
.B1(n_366),
.B2(n_451),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_572),
.B(n_570),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_601),
.A2(n_423),
.B1(n_466),
.B2(n_395),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_575),
.A2(n_376),
.B1(n_366),
.B2(n_466),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_611),
.A2(n_376),
.B1(n_366),
.B2(n_423),
.Y(n_629)
);

AOI222xp33_ASAP7_75t_L g630 ( 
.A1(n_582),
.A2(n_595),
.B1(n_570),
.B2(n_577),
.C1(n_603),
.C2(n_593),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_572),
.A2(n_366),
.B1(n_437),
.B2(n_457),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_567),
.A2(n_393),
.B1(n_545),
.B2(n_471),
.Y(n_632)
);

OAI222xp33_ASAP7_75t_L g633 ( 
.A1(n_592),
.A2(n_448),
.B1(n_458),
.B2(n_477),
.C1(n_496),
.C2(n_482),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_576),
.B(n_412),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_SL g635 ( 
.A1(n_577),
.A2(n_540),
.B1(n_547),
.B2(n_491),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_567),
.A2(n_600),
.B1(n_608),
.B2(n_609),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_578),
.A2(n_365),
.B1(n_517),
.B2(n_448),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_586),
.A2(n_365),
.B1(n_517),
.B2(n_482),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_604),
.A2(n_365),
.B1(n_517),
.B2(n_482),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_602),
.Y(n_640)
);

AOI221xp5_ASAP7_75t_L g641 ( 
.A1(n_605),
.A2(n_412),
.B1(n_380),
.B2(n_398),
.C(n_411),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_566),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_599),
.B(n_477),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_614),
.A2(n_612),
.B1(n_607),
.B2(n_613),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_566),
.B(n_412),
.Y(n_645)
);

OAI221xp5_ASAP7_75t_SL g646 ( 
.A1(n_610),
.A2(n_380),
.B1(n_482),
.B2(n_477),
.C(n_496),
.Y(n_646)
);

OAI222xp33_ASAP7_75t_L g647 ( 
.A1(n_592),
.A2(n_477),
.B1(n_496),
.B2(n_505),
.C1(n_547),
.C2(n_491),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_580),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_607),
.A2(n_365),
.B1(n_496),
.B2(n_505),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_SL g650 ( 
.A1(n_573),
.A2(n_491),
.B1(n_484),
.B2(n_481),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_626),
.B(n_580),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_615),
.B(n_606),
.Y(n_652)
);

NOR3xp33_ASAP7_75t_L g653 ( 
.A(n_615),
.B(n_612),
.C(n_573),
.Y(n_653)
);

OAI21xp33_ASAP7_75t_L g654 ( 
.A1(n_618),
.A2(n_606),
.B(n_398),
.Y(n_654)
);

OAI221xp5_ASAP7_75t_SL g655 ( 
.A1(n_630),
.A2(n_621),
.B1(n_636),
.B2(n_624),
.C(n_644),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_623),
.B(n_573),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_623),
.B(n_479),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_640),
.B(n_479),
.Y(n_658)
);

NAND3xp33_ASAP7_75t_L g659 ( 
.A(n_618),
.B(n_200),
.C(n_484),
.Y(n_659)
);

NOR3xp33_ASAP7_75t_L g660 ( 
.A(n_632),
.B(n_633),
.C(n_616),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g661 ( 
.A1(n_617),
.A2(n_484),
.B(n_481),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_646),
.A2(n_521),
.B1(n_486),
.B2(n_505),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_640),
.B(n_479),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_642),
.B(n_479),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_622),
.A2(n_521),
.B1(n_486),
.B2(n_365),
.Y(n_665)
);

OA211x2_ASAP7_75t_L g666 ( 
.A1(n_641),
.A2(n_649),
.B(n_637),
.C(n_638),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_634),
.A2(n_521),
.B1(n_486),
.B2(n_218),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_642),
.B(n_479),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_639),
.A2(n_635),
.B1(n_631),
.B2(n_620),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_627),
.B(n_481),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_627),
.B(n_484),
.C(n_481),
.Y(n_671)
);

OA21x2_ASAP7_75t_L g672 ( 
.A1(n_647),
.A2(n_410),
.B(n_521),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_650),
.B(n_481),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_648),
.B(n_643),
.Y(n_674)
);

NAND4xp25_ASAP7_75t_SL g675 ( 
.A(n_625),
.B(n_51),
.C(n_53),
.D(n_54),
.Y(n_675)
);

OAI211xp5_ASAP7_75t_SL g676 ( 
.A1(n_628),
.A2(n_449),
.B(n_58),
.C(n_59),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_629),
.A2(n_484),
.B1(n_481),
.B2(n_440),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_648),
.B(n_484),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_SL g679 ( 
.A1(n_659),
.A2(n_643),
.B1(n_619),
.B2(n_645),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_L g680 ( 
.A(n_653),
.B(n_205),
.C(n_221),
.Y(n_680)
);

AO21x2_ASAP7_75t_L g681 ( 
.A1(n_653),
.A2(n_410),
.B(n_60),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_655),
.B(n_56),
.C(n_61),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_656),
.B(n_674),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_663),
.B(n_62),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_651),
.B(n_63),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_657),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_652),
.B(n_65),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_658),
.B(n_67),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_661),
.B(n_68),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_666),
.A2(n_675),
.B1(n_660),
.B2(n_669),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_660),
.B(n_221),
.C(n_210),
.Y(n_691)
);

NAND3xp33_ASAP7_75t_L g692 ( 
.A(n_654),
.B(n_671),
.C(n_676),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_664),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_673),
.B(n_70),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_668),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_695),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_683),
.B(n_672),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_686),
.Y(n_698)
);

NOR3xp33_ASAP7_75t_SL g699 ( 
.A(n_691),
.B(n_677),
.C(n_662),
.Y(n_699)
);

INVxp67_ASAP7_75t_SL g700 ( 
.A(n_695),
.Y(n_700)
);

NAND4xp75_ASAP7_75t_L g701 ( 
.A(n_690),
.B(n_670),
.C(n_672),
.D(n_678),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_693),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_693),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_683),
.B(n_667),
.Y(n_704)
);

NAND4xp75_ASAP7_75t_L g705 ( 
.A(n_689),
.B(n_665),
.C(n_72),
.D(n_73),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_686),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_698),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_704),
.B(n_687),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_702),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_698),
.Y(n_710)
);

XNOR2x1_ASAP7_75t_L g711 ( 
.A(n_701),
.B(n_685),
.Y(n_711)
);

OA22x2_ASAP7_75t_L g712 ( 
.A1(n_711),
.A2(n_697),
.B1(n_700),
.B2(n_696),
.Y(n_712)
);

OA22x2_ASAP7_75t_L g713 ( 
.A1(n_707),
.A2(n_697),
.B1(n_696),
.B2(n_706),
.Y(n_713)
);

XNOR2x1_ASAP7_75t_L g714 ( 
.A(n_708),
.B(n_701),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_710),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_713),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_714),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_715),
.Y(n_718)
);

AOI322xp5_ASAP7_75t_L g719 ( 
.A1(n_712),
.A2(n_682),
.A3(n_699),
.B1(n_689),
.B2(n_679),
.C1(n_694),
.C2(n_709),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_718),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_716),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_717),
.A2(n_705),
.B1(n_681),
.B2(n_694),
.Y(n_722)
);

OAI22x1_ASAP7_75t_L g723 ( 
.A1(n_722),
.A2(n_716),
.B1(n_719),
.B2(n_680),
.Y(n_723)
);

AO22x2_ASAP7_75t_L g724 ( 
.A1(n_721),
.A2(n_709),
.B1(n_705),
.B2(n_692),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_720),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_721),
.Y(n_726)
);

NOR2x1_ASAP7_75t_L g727 ( 
.A(n_726),
.B(n_681),
.Y(n_727)
);

NOR2x1_ASAP7_75t_L g728 ( 
.A(n_725),
.B(n_684),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_723),
.B(n_703),
.Y(n_729)
);

NAND4xp25_ASAP7_75t_SL g730 ( 
.A(n_724),
.B(n_684),
.C(n_665),
.D(n_688),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_726),
.Y(n_731)
);

AOI221xp5_ASAP7_75t_L g732 ( 
.A1(n_723),
.A2(n_695),
.B1(n_221),
.B2(n_75),
.C(n_77),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_723),
.B(n_695),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_731),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_733),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_729),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_728),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_730),
.A2(n_365),
.B1(n_436),
.B2(n_440),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_732),
.B(n_71),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_727),
.A2(n_365),
.B1(n_436),
.B2(n_210),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_L g741 ( 
.A1(n_735),
.A2(n_737),
.B1(n_739),
.B2(n_736),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_734),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_738),
.B(n_74),
.Y(n_743)
);

AND4x1_ASAP7_75t_L g744 ( 
.A(n_740),
.B(n_81),
.C(n_82),
.D(n_83),
.Y(n_744)
);

AO22x2_ASAP7_75t_L g745 ( 
.A1(n_735),
.A2(n_84),
.B1(n_88),
.B2(n_89),
.Y(n_745)
);

OR3x2_ASAP7_75t_L g746 ( 
.A(n_737),
.B(n_90),
.C(n_91),
.Y(n_746)
);

AO22x2_ASAP7_75t_L g747 ( 
.A1(n_735),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_735),
.A2(n_365),
.B1(n_210),
.B2(n_98),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_742),
.Y(n_749)
);

AO22x1_ASAP7_75t_L g750 ( 
.A1(n_743),
.A2(n_95),
.B1(n_97),
.B2(n_101),
.Y(n_750)
);

AO22x1_ASAP7_75t_L g751 ( 
.A1(n_746),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_751)
);

OA22x2_ASAP7_75t_L g752 ( 
.A1(n_748),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_745),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_747),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_741),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_755),
.A2(n_744),
.B1(n_110),
.B2(n_111),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_749),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_753),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_754),
.A2(n_109),
.B1(n_112),
.B2(n_114),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_752),
.Y(n_760)
);

OAI211xp5_ASAP7_75t_SL g761 ( 
.A1(n_751),
.A2(n_115),
.B(n_118),
.C(n_119),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_757),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_760),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_758),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_763),
.A2(n_756),
.B1(n_761),
.B2(n_759),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_764),
.A2(n_750),
.B1(n_121),
.B2(n_122),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_L g767 ( 
.A1(n_762),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_765),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_766),
.B1(n_767),
.B2(n_130),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_769),
.Y(n_770)
);

AOI221x1_ASAP7_75t_L g771 ( 
.A1(n_770),
.A2(n_125),
.B1(n_129),
.B2(n_132),
.C(n_133),
.Y(n_771)
);

AOI211xp5_ASAP7_75t_L g772 ( 
.A1(n_771),
.A2(n_134),
.B(n_135),
.C(n_137),
.Y(n_772)
);


endmodule