module real_aes_8346_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_17;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_20;
wire n_18;
wire n_21;
wire n_7;
wire n_8;
wire n_10;
INVx1_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_1), .B(n_14), .Y(n_18) );
INVx1_ASAP7_75t_L g21 ( .A(n_1), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g6 ( .A1(n_2), .A2(n_7), .B1(n_19), .B2(n_20), .Y(n_6) );
INVxp67_ASAP7_75t_L g19 ( .A(n_2), .Y(n_19) );
NAND3xp33_ASAP7_75t_SL g9 ( .A(n_3), .B(n_10), .C(n_11), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_4), .Y(n_10) );
INVx1_ASAP7_75t_L g17 ( .A(n_5), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g7 ( .A(n_8), .Y(n_7) );
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_14), .B(n_18), .Y(n_8) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
CKINVDCx16_ASAP7_75t_R g14 ( .A(n_15), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
NOR2xp33_ASAP7_75t_SL g20 ( .A(n_16), .B(n_21), .Y(n_20) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
endmodule