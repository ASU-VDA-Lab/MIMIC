module fake_jpeg_21950_n_108 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_29),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_18),
.Y(n_28)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_1),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_23),
.B1(n_14),
.B2(n_17),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_13),
.B1(n_17),
.B2(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_16),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_50),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_12),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_12),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_25),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_36),
.B1(n_27),
.B2(n_21),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_64),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_21),
.B1(n_13),
.B2(n_14),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_40),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_22),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_29),
.C(n_26),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_48),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_34),
.B1(n_33),
.B2(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_75),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_74),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_48),
.C(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_40),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_59),
.B1(n_52),
.B2(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_81),
.C(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_42),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_42),
.B(n_41),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_19),
.B(n_1),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_34),
.B1(n_33),
.B2(n_41),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_71),
.B(n_74),
.C(n_22),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_86),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_80),
.C(n_78),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_66),
.C(n_71),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_90),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_82),
.B1(n_76),
.B2(n_83),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_65),
.C(n_22),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_2),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_19),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_3),
.B(n_5),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_100),
.B(n_7),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_6),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_93),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_99),
.Y(n_104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_105),
.B(n_102),
.C(n_8),
.D(n_19),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_92),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_92),
.Y(n_108)
);


endmodule