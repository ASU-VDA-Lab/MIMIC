module real_jpeg_4505_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_0),
.B(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_0),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_0),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_0),
.B(n_237),
.Y(n_236)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_2),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_2),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_2),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_2),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g295 ( 
.A(n_2),
.B(n_83),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_2),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_2),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_2),
.B(n_395),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_3),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_4),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_4),
.Y(n_141)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_4),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_5),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_5),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_5),
.B(n_122),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_5),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_5),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_5),
.B(n_61),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_5),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_5),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_6),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_6),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_6),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_6),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_6),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_6),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_6),
.B(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_8),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_8),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_8),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_8),
.B(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_8),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_8),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_8),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_8),
.B(n_331),
.Y(n_330)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_9),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_9),
.Y(n_429)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_10),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_12),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_12),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_12),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_12),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_12),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_12),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_12),
.B(n_420),
.Y(n_419)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_13),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_13),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_13),
.Y(n_324)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_14),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_15),
.B(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_15),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_15),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_15),
.B(n_180),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_15),
.B(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_16),
.Y(n_186)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_16),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_16),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_17),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_17),
.B(n_30),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_17),
.B(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_17),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_17),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_17),
.B(n_414),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_504),
.B(n_506),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_68),
.B(n_105),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_21),
.B(n_68),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.C(n_32),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_24),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_32),
.B1(n_44),
.B2(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_24),
.B(n_227),
.Y(n_226)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_27),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_27),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_27),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_28),
.A2(n_29),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_28),
.A2(n_29),
.B1(n_329),
.B2(n_335),
.Y(n_328)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_29),
.B(n_330),
.C(n_334),
.Y(n_485)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_31),
.Y(n_246)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_32),
.A2(n_54),
.B1(n_59),
.B2(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_32),
.A2(n_54),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_32),
.B(n_149),
.C(n_154),
.Y(n_248)
);

OR2x2_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_36),
.Y(n_135)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_36),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_36),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_60),
.Y(n_59)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_37),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_37),
.B(n_323),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_41),
.A2(n_42),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_41),
.A2(n_42),
.B1(n_347),
.B2(n_350),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_41),
.B(n_343),
.C(n_350),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_42),
.B(n_306),
.C(n_310),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_44),
.B(n_228),
.C(n_230),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_45),
.A2(n_46),
.B1(n_72),
.B2(n_73),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_59),
.C(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_47),
.Y(n_177)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.C(n_58),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_50),
.A2(n_51),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_59),
.C(n_64),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_99),
.B1(n_117),
.B2(n_120),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_59),
.B(n_117),
.C(n_121),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_59),
.A2(n_99),
.B1(n_480),
.B2(n_481),
.Y(n_479)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_62),
.B(n_169),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_63),
.Y(n_372)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_63),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_65),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_64),
.A2(n_65),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_64),
.B(n_193),
.C(n_289),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_100),
.C(n_101),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_69),
.B(n_501),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_86),
.C(n_96),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_70),
.B(n_492),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_82),
.C(n_84),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_72),
.A2(n_73),
.B1(n_131),
.B2(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_72),
.A2(n_73),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_128),
.C(n_131),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_73),
.B(n_193),
.C(n_322),
.Y(n_484)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_86),
.B(n_96),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.C(n_92),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_87),
.A2(n_89),
.B1(n_90),
.B2(n_475),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_87),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_89),
.A2(n_90),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_90),
.B(n_138),
.C(n_236),
.Y(n_310)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_92),
.B(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_100),
.B(n_101),
.Y(n_501)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_499),
.B(n_503),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_467),
.B(n_496),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_351),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_278),
.B(n_312),
.C(n_313),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_249),
.B(n_277),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_111),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_220),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_112),
.B(n_220),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_173),
.C(n_204),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_113),
.B(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_145),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_114),
.B(n_146),
.C(n_156),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_127),
.C(n_136),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_115),
.B(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx8_ASAP7_75t_L g363 ( 
.A(n_126),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g426 ( 
.A(n_126),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_127),
.A2(n_136),
.B1(n_137),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_127),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_128),
.B(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_130),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_131),
.Y(n_258)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_135),
.Y(n_270)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_138),
.A2(n_235),
.B1(n_236),
.B2(n_238),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_138),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_138),
.A2(n_142),
.B1(n_143),
.B2(n_238),
.Y(n_271)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_141),
.Y(n_417)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_156),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_154),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_150),
.B(n_193),
.Y(n_367)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_152),
.Y(n_237)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_152),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_152),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_158),
.B(n_159),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_157),
.B(n_164),
.C(n_168),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_173),
.B(n_204),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_188),
.C(n_190),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_174),
.A2(n_188),
.B1(n_189),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_174),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_179),
.C(n_183),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_176),
.B(n_425),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_176),
.B(n_432),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_182),
.B1(n_183),
.B2(n_187),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_182),
.A2(n_183),
.B1(n_294),
.B2(n_297),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_183),
.B(n_236),
.C(n_295),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_185),
.Y(n_366)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_186),
.Y(n_409)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_190),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_197),
.C(n_200),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_191),
.A2(n_192),
.B1(n_454),
.B2(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_193),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_193),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_193),
.A2(n_286),
.B1(n_322),
.B2(n_325),
.Y(n_321)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_196),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_455)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_219),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_207),
.C(n_219),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_214),
.C(n_217),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_214),
.A2(n_330),
.B1(n_333),
.B2(n_334),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_214),
.Y(n_334)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_221),
.B(n_223),
.C(n_239),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_239),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_232),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_225),
.B(n_226),
.C(n_232),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_235),
.A2(n_236),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_235),
.A2(n_236),
.B1(n_359),
.B2(n_360),
.Y(n_396)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_236),
.B(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_240),
.B(n_242),
.C(n_243),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_245),
.B(n_247),
.C(n_302),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_275),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_250),
.B(n_275),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_255),
.C(n_272),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_251),
.A2(n_252),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_255),
.B(n_272),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.C(n_271),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_256),
.B(n_449),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_259),
.B(n_271),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_265),
.C(n_266),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_260),
.A2(n_261),
.B1(n_266),
.B2(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_265),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_266),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_267),
.B(n_371),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_267),
.B(n_428),
.Y(n_427)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_279),
.B(n_314),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_281),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_315),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_281),
.B(n_315),
.Y(n_466)
);

FAx1_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_298),
.CI(n_311),
.CON(n_281),
.SN(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_293),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_285),
.C(n_293),
.Y(n_338)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_295),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_301),
.C(n_303),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_310),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_316),
.B(n_318),
.C(n_336),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_336),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_326),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_319),
.B(n_327),
.C(n_328),
.Y(n_476)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

INVx8_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_329),
.Y(n_335)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_330),
.Y(n_333)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_337),
.B(n_341),
.C(n_342),
.Y(n_486)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

AO22x1_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_345),
.B2(n_346),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_347),
.Y(n_350)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OAI31xp33_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_463),
.A3(n_464),
.B(n_466),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_457),
.B(n_462),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_444),
.B(n_456),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_397),
.B(n_443),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_383),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_356),
.B(n_383),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_368),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_357),
.B(n_369),
.C(n_380),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_364),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_358),
.B(n_365),
.C(n_367),
.Y(n_452)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_380),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_373),
.C(n_375),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_370),
.B(n_385),
.Y(n_384)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_373),
.A2(n_374),
.B1(n_375),
.B2(n_376),
.Y(n_385)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx8_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.C(n_396),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_384),
.B(n_440),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_386),
.A2(n_387),
.B1(n_396),
.B2(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_393),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_388),
.A2(n_389),
.B1(n_393),
.B2(n_394),
.Y(n_410)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_396),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_437),
.B(n_442),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_422),
.B(n_436),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_411),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_411),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_410),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_408),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_402),
.B(n_408),
.C(n_410),
.Y(n_438)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx5_ASAP7_75t_SL g404 ( 
.A(n_405),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_418),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_412),
.A2(n_413),
.B1(n_418),
.B2(n_419),
.Y(n_434)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx6_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx8_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_430),
.B(n_435),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_427),
.Y(n_423)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_434),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_431),
.B(n_434),
.Y(n_435)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_439),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_446),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_447),
.A2(n_448),
.B1(n_450),
.B2(n_451),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_452),
.C(n_453),
.Y(n_461)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_461),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_458),
.B(n_461),
.Y(n_462)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_459),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_493),
.Y(n_467)
);

OAI21xp33_ASAP7_75t_L g496 ( 
.A1(n_468),
.A2(n_497),
.B(n_498),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_487),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_469),
.B(n_487),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_477),
.C(n_486),
.Y(n_469)
);

FAx1_ASAP7_75t_SL g495 ( 
.A(n_470),
.B(n_477),
.CI(n_486),
.CON(n_495),
.SN(n_495)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_476),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_473),
.C(n_476),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_482),
.B2(n_483),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_484),
.C(n_485),
.Y(n_490)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_490),
.C(n_491),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_495),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_494),
.B(n_495),
.Y(n_497)
);

BUFx24_ASAP7_75t_SL g510 ( 
.A(n_495),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_502),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_500),
.B(n_502),
.Y(n_503)
);

INVx6_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx13_ASAP7_75t_L g508 ( 
.A(n_505),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_509),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);


endmodule