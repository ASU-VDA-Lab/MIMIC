module real_jpeg_23417_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_0),
.A2(n_57),
.B1(n_60),
.B2(n_63),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_0),
.A2(n_63),
.B1(n_66),
.B2(n_71),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_0),
.A2(n_41),
.B1(n_43),
.B2(n_63),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_0),
.A2(n_27),
.B1(n_35),
.B2(n_63),
.Y(n_224)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_2),
.A2(n_66),
.B1(n_71),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_41),
.B1(n_43),
.B2(n_88),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_2),
.A2(n_58),
.B1(n_88),
.B2(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_2),
.A2(n_27),
.B1(n_35),
.B2(n_88),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_3),
.B(n_136),
.Y(n_191)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_3),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_3),
.B(n_65),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_3),
.B(n_41),
.C(n_84),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_3),
.A2(n_66),
.B1(n_71),
.B2(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_3),
.B(n_127),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_3),
.A2(n_41),
.B1(n_43),
.B2(n_215),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_3),
.B(n_27),
.C(n_46),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_3),
.A2(n_26),
.B(n_276),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_6),
.A2(n_57),
.B1(n_76),
.B2(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_6),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_6),
.A2(n_66),
.B1(n_71),
.B2(n_164),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_6),
.A2(n_41),
.B1(n_43),
.B2(n_164),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_6),
.A2(n_27),
.B1(n_35),
.B2(n_164),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_8),
.A2(n_40),
.B1(n_66),
.B2(n_71),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_8),
.A2(n_40),
.B1(n_137),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_27),
.B1(n_35),
.B2(n_40),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_9),
.A2(n_57),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_9),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_9),
.A2(n_66),
.B1(n_71),
.B2(n_75),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_9),
.A2(n_41),
.B1(n_43),
.B2(n_75),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_9),
.A2(n_27),
.B1(n_35),
.B2(n_75),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_12),
.A2(n_57),
.B1(n_76),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_12),
.A2(n_66),
.B1(n_71),
.B2(n_112),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_12),
.A2(n_41),
.B1(n_43),
.B2(n_112),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_12),
.A2(n_27),
.B1(n_35),
.B2(n_112),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_14),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_14),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_14),
.A2(n_36),
.B1(n_66),
.B2(n_71),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_14),
.A2(n_36),
.B1(n_60),
.B2(n_61),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_15),
.A2(n_41),
.B1(n_43),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_15),
.A2(n_27),
.B1(n_35),
.B2(n_50),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_15),
.A2(n_50),
.B1(n_66),
.B2(n_71),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_15),
.A2(n_50),
.B1(n_60),
.B2(n_61),
.Y(n_344)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_16),
.Y(n_225)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_16),
.Y(n_290)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_354),
.B(n_357),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_349),
.B(n_353),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_336),
.B(n_348),
.Y(n_19)
);

OAI31xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_139),
.A3(n_154),
.B(n_333),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_116),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_22),
.B(n_116),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_79),
.C(n_95),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_23),
.A2(n_79),
.B1(n_80),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_23),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_52),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_24),
.A2(n_25),
.B(n_54),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_25),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_25),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_25),
.A2(n_37),
.B1(n_38),
.B2(n_53),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_26),
.A2(n_34),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_26),
.A2(n_31),
.B1(n_100),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_26),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_26),
.A2(n_188),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_26),
.B(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_26),
.A2(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_48)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_28),
.Y(n_189)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_32),
.B(n_277),
.Y(n_276)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_33),
.B(n_215),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_35),
.B(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_39),
.A2(n_44),
.B1(n_51),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_41),
.A2(n_43),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_41),
.B(n_283),
.Y(n_282)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_44),
.A2(n_51),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_44),
.B(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_44),
.A2(n_51),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_48),
.A2(n_91),
.B1(n_106),
.B2(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_48),
.A2(n_174),
.B(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_48),
.A2(n_211),
.B(n_249),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_48),
.B(n_215),
.Y(n_296)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_51),
.B(n_212),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_64),
.B(n_72),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_56),
.A2(n_64),
.B1(n_113),
.B2(n_135),
.Y(n_134)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_59),
.B1(n_69),
.B2(n_70),
.Y(n_78)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_60),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_74),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_64),
.A2(n_113),
.B1(n_135),
.B2(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_64),
.A2(n_72),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_65),
.A2(n_77),
.B1(n_111),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_65),
.A2(n_77),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_65),
.A2(n_77),
.B1(n_344),
.B2(n_351),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_65),
.A2(n_77),
.B(n_351),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_65)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_71),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g192 ( 
.A(n_66),
.B(n_70),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_66),
.B(n_240),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI32xp33_ASAP7_75t_L g190 ( 
.A1(n_69),
.A2(n_71),
.A3(n_76),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_77),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_77),
.A2(n_115),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_90),
.B(n_94),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_90),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_89),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_82),
.A2(n_83),
.B1(n_129),
.B2(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_82),
.A2(n_181),
.B(n_183),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_82),
.A2(n_183),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_83),
.A2(n_108),
.B(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_83),
.A2(n_167),
.B(n_220),
.Y(n_219)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_91),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_91),
.A2(n_264),
.B(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_93),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_95),
.A2(n_96),
.B1(n_328),
.B2(n_330),
.Y(n_327)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.C(n_109),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_97),
.A2(n_98),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_99),
.Y(n_176)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_107),
.B(n_109),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B(n_114),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_119),
.C(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_134),
.B2(n_138),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_131),
.C(n_134),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_126),
.B(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_126),
.A2(n_127),
.B1(n_182),
.B2(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_126),
.A2(n_127),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_127),
.B(n_168),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_131),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_131),
.B(n_146),
.C(n_151),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_138),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_134),
.B(n_142),
.C(n_145),
.Y(n_337)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_140),
.A2(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_153),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_141),
.B(n_153),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_147),
.Y(n_343)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_152),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_326),
.B(n_332),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_200),
.B(n_325),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_193),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_157),
.B(n_193),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_175),
.C(n_177),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_158),
.A2(n_159),
.B1(n_175),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_169),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_165),
.C(n_169),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_163),
.Y(n_179)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_170),
.B(n_173),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_185)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_175),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_177),
.B(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_184),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_180),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_184),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_190),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_190),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_186),
.A2(n_287),
.B1(n_289),
.B2(n_291),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_195),
.B(n_196),
.C(n_199),
.Y(n_331)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_232),
.B(n_319),
.C(n_324),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_226),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_226),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_217),
.C(n_218),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_203),
.A2(n_204),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_213),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_209),
.C(n_213),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_217),
.B(n_218),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.C(n_223),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_225),
.A2(n_288),
.B(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_227),
.B(n_230),
.C(n_231),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_313),
.B(n_318),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_265),
.B(n_312),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_254),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_237),
.B(n_254),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_247),
.C(n_251),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_238),
.B(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_241),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B(n_245),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_247),
.A2(n_251),
.B1(n_252),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_250),
.Y(n_263)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_255),
.B(n_261),
.C(n_262),
.Y(n_317)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_306),
.B(n_311),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_284),
.B(n_305),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_278),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_278),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_274),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_273),
.C(n_274),
.Y(n_310)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_275),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_282),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_294),
.B(n_304),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_292),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_292),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_299),
.B(n_303),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_297),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_310),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_317),
.Y(n_318)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_321),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_331),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_331),
.Y(n_332)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_328),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_338),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_347),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_342),
.B1(n_345),
.B2(n_346),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_340),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_342),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_345),
.C(n_347),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_352),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_350),
.B(n_355),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_350),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_356),
.B(n_359),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_358),
.Y(n_357)
);


endmodule