module fake_jpeg_3524_n_218 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_218);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_218;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

INVxp33_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_40),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_80),
.Y(n_87)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_67),
.Y(n_91)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_84),
.Y(n_95)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_83),
.A2(n_63),
.B1(n_60),
.B2(n_58),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_58),
.B1(n_66),
.B2(n_54),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_63),
.B1(n_66),
.B2(n_54),
.Y(n_89)
);

HAxp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_56),
.CON(n_90),
.SN(n_90)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_70),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_61),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_52),
.B1(n_53),
.B2(n_73),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_69),
.B1(n_78),
.B2(n_62),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_68),
.Y(n_106)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_104),
.Y(n_135)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_103),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_80),
.B1(n_82),
.B2(n_72),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_113),
.B1(n_87),
.B2(n_2),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_110),
.C(n_8),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_80),
.B1(n_68),
.B2(n_57),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_71),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_55),
.B(n_62),
.C(n_70),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_0),
.B(n_4),
.C(n_5),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_70),
.B1(n_2),
.B2(n_3),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_115),
.C(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_120),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_117),
.B(n_133),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_129),
.B1(n_10),
.B2(n_13),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_104),
.Y(n_120)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_6),
.B(n_7),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_107),
.B(n_11),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_9),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_132),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_99),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_127),
.B(n_8),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_143),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_10),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_107),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_148),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_111),
.B(n_112),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_156),
.B(n_157),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_48),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_159),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_13),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_151),
.B(n_152),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_14),
.B(n_16),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_17),
.B(n_18),
.Y(n_157)
);

AO22x1_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_36),
.B1(n_46),
.B2(n_21),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_123),
.C(n_124),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_147),
.C(n_150),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_158),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_162),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_144),
.A2(n_124),
.B1(n_19),
.B2(n_18),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_167),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_172),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_153),
.B(n_34),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_174),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_47),
.B1(n_39),
.B2(n_41),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_176),
.A2(n_157),
.B(n_145),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_146),
.C(n_162),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_150),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_166),
.Y(n_192)
);

BUFx12f_ASAP7_75t_SL g183 ( 
.A(n_165),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_191),
.Y(n_199)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_194),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_188),
.B1(n_165),
.B2(n_178),
.Y(n_193)
);

NOR2xp67_ASAP7_75t_SL g201 ( 
.A(n_193),
.B(n_196),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_164),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_164),
.B1(n_137),
.B2(n_175),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_181),
.A2(n_175),
.B1(n_176),
.B2(n_148),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_198),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_180),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_186),
.C(n_168),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_203),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_159),
.C(n_163),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_199),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_205),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_204),
.B(n_192),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_206),
.C(n_198),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_211),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_201),
.C(n_187),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_159),
.Y(n_213)
);

HAxp5_ASAP7_75t_SL g214 ( 
.A(n_213),
.B(n_183),
.CON(n_214),
.SN(n_214)
);

OAI311xp33_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_170),
.A3(n_173),
.B1(n_177),
.C1(n_45),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_37),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_42),
.B(n_44),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_208),
.Y(n_218)
);


endmodule