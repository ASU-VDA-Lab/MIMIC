module fake_jpeg_30337_n_244 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_244);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_96;

INVxp67_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_52),
.Y(n_71)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_27),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_58),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_0),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_60),
.Y(n_70)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_8),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_30),
.B(n_9),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_76),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_86),
.B1(n_39),
.B2(n_34),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_36),
.B1(n_42),
.B2(n_34),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_26),
.B1(n_44),
.B2(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_33),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_80),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_58),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_25),
.C(n_19),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_45),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_42),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_38),
.B1(n_25),
.B2(n_22),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_33),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_56),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_19),
.Y(n_104)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_61),
.B1(n_55),
.B2(n_63),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_94),
.A2(n_98),
.B1(n_102),
.B2(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_117),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_57),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_106),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_49),
.B1(n_50),
.B2(n_47),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_65),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_104),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_87),
.B1(n_79),
.B2(n_74),
.Y(n_126)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g141 ( 
.A(n_107),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_91),
.B1(n_73),
.B2(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_40),
.B1(n_37),
.B2(n_2),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_115),
.B(n_118),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_40),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_112),
.B(n_116),
.Y(n_124)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_82),
.Y(n_123)
);

NAND2x1_ASAP7_75t_SL g115 ( 
.A(n_81),
.B(n_40),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_40),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_70),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_67),
.A2(n_37),
.B1(n_3),
.B2(n_5),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_120),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_69),
.Y(n_121)
);

CKINVDCx12_ASAP7_75t_R g127 ( 
.A(n_121),
.Y(n_127)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_67),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_123),
.B(n_130),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_126),
.A2(n_108),
.B1(n_140),
.B2(n_102),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_95),
.B(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_99),
.B(n_14),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_100),
.B(n_18),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_145),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_159),
.B1(n_139),
.B2(n_125),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_106),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_106),
.C(n_97),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_154),
.C(n_155),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_151),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_108),
.C(n_96),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_105),
.C(n_110),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_115),
.B(n_117),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_92),
.C(n_115),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_142),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_120),
.B1(n_94),
.B2(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_172),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_131),
.B1(n_134),
.B2(n_139),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_170),
.B1(n_147),
.B2(n_149),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_132),
.B1(n_135),
.B2(n_133),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_133),
.B1(n_124),
.B2(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_184),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_179),
.B1(n_186),
.B2(n_167),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_138),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_147),
.B1(n_155),
.B2(n_156),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_157),
.B(n_154),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_162),
.B(n_167),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_132),
.C(n_124),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_188),
.C(n_143),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_150),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_166),
.B1(n_174),
.B2(n_172),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_128),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_162),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_192),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_186),
.B1(n_183),
.B2(n_187),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_184),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_196),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_177),
.B(n_185),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_183),
.B(n_175),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_188),
.B(n_153),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_198),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_128),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_197),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_207),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_165),
.B1(n_129),
.B2(n_143),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_198),
.Y(n_208)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_212),
.C(n_129),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_165),
.B(n_128),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_211),
.A2(n_113),
.B(n_114),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_119),
.C(n_137),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_136),
.Y(n_214)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_217),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_111),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_203),
.C(n_209),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_221),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_93),
.CI(n_5),
.CON(n_221),
.SN(n_221)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_208),
.B(n_202),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_224),
.B(n_213),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_215),
.A2(n_202),
.B(n_204),
.Y(n_224)
);

OAI21x1_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_209),
.B(n_10),
.Y(n_226)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_226),
.A2(n_217),
.B(n_10),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_220),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_219),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_230),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_231),
.A2(n_232),
.B(n_11),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_221),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_221),
.C(n_225),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_235),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_225),
.B(n_216),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_74),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_236),
.C(n_79),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_241),
.B1(n_12),
.B2(n_7),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);


endmodule