module fake_jpeg_29504_n_421 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_421);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_421;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_133;
wire n_132;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_48),
.Y(n_140)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_53),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_21),
.B(n_22),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_55),
.B(n_56),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_14),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_1),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_84),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_31),
.Y(n_65)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_70),
.Y(n_114)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_23),
.B(n_30),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_74),
.Y(n_121)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_23),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_79),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_83),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_88),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_42),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_87),
.B(n_25),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_14),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_90),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_20),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_78),
.B1(n_79),
.B2(n_77),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_92),
.A2(n_97),
.B1(n_104),
.B2(n_108),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_27),
.C(n_16),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_95),
.B(n_58),
.C(n_59),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_91),
.B1(n_60),
.B2(n_63),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_47),
.A2(n_16),
.B1(n_27),
.B2(n_28),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_48),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_109),
.B1(n_124),
.B2(n_141),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_49),
.A2(n_28),
.B1(n_38),
.B2(n_18),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_25),
.B1(n_30),
.B2(n_34),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_65),
.A2(n_39),
.B1(n_20),
.B2(n_33),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_116),
.A2(n_130),
.B1(n_131),
.B2(n_142),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_51),
.A2(n_18),
.B1(n_44),
.B2(n_33),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_67),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_75),
.A2(n_45),
.B1(n_41),
.B2(n_36),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_80),
.B(n_41),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_110),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_65),
.A2(n_84),
.B1(n_62),
.B2(n_90),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_68),
.A2(n_36),
.B1(n_34),
.B2(n_9),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_83),
.A2(n_1),
.B(n_2),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_86),
.A2(n_69),
.B1(n_85),
.B2(n_57),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_72),
.A2(n_8),
.B1(n_9),
.B2(n_4),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_55),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_144),
.B(n_170),
.Y(n_213)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_146),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_148),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_82),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_149),
.B(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_150),
.B(n_152),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_107),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_157),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_154),
.B(n_185),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_81),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_159),
.Y(n_195)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_76),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_120),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_112),
.B(n_114),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_162),
.B(n_168),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_100),
.Y(n_167)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_113),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_8),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_95),
.B(n_66),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_174),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_119),
.B(n_61),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_96),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_184),
.Y(n_207)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_118),
.A2(n_89),
.B1(n_3),
.B2(n_5),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_135),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_2),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_5),
.B(n_6),
.Y(n_215)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_102),
.B(n_3),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_147),
.A2(n_105),
.B1(n_103),
.B2(n_128),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_147),
.A2(n_103),
.B1(n_128),
.B2(n_111),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_147),
.A2(n_126),
.B1(n_136),
.B2(n_133),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_144),
.A2(n_126),
.B1(n_135),
.B2(n_102),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_135),
.B1(n_127),
.B2(n_137),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_183),
.B1(n_158),
.B2(n_149),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_183),
.B(n_154),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_127),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_155),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_172),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_250),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_224),
.A2(n_235),
.B1(n_248),
.B2(n_249),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_225),
.A2(n_189),
.B(n_5),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_213),
.B(n_148),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_226),
.B(n_230),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_184),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_227),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_188),
.A2(n_151),
.B1(n_180),
.B2(n_145),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_238),
.B1(n_214),
.B2(n_215),
.Y(n_258)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_185),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_231),
.B(n_244),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_188),
.C(n_195),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_236),
.C(n_246),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_200),
.A2(n_145),
.B1(n_185),
.B2(n_137),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_158),
.C(n_149),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_218),
.A2(n_185),
.B1(n_163),
.B2(n_160),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_117),
.Y(n_239)
);

AO22x1_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_193),
.B1(n_238),
.B2(n_224),
.Y(n_261)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_192),
.B(n_143),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_242),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_190),
.B(n_167),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_245),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_161),
.C(n_157),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_166),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_251),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_167),
.B(n_177),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_187),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_211),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_199),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_216),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_223),
.A2(n_201),
.B1(n_210),
.B2(n_203),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_256),
.A2(n_258),
.B1(n_264),
.B2(n_272),
.Y(n_293)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_261),
.A2(n_245),
.B1(n_243),
.B2(n_125),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_193),
.C(n_220),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_234),
.C(n_250),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_223),
.A2(n_209),
.B1(n_211),
.B2(n_220),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_228),
.A2(n_212),
.B1(n_197),
.B2(n_125),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_268),
.A2(n_253),
.B(n_229),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_236),
.A2(n_202),
.B1(n_197),
.B2(n_212),
.Y(n_272)
);

OAI32xp33_ASAP7_75t_L g274 ( 
.A1(n_231),
.A2(n_217),
.A3(n_208),
.B1(n_194),
.B2(n_191),
.Y(n_274)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_239),
.A2(n_202),
.B1(n_189),
.B2(n_194),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_275),
.A2(n_208),
.B1(n_233),
.B2(n_165),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_225),
.Y(n_300)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_282),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_241),
.Y(n_283)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_283),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_286),
.C(n_299),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_246),
.C(n_230),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_282),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_288),
.B(n_296),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_239),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_289),
.B(n_306),
.Y(n_330)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_290),
.Y(n_310)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_281),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_294),
.Y(n_309)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_281),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_255),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_305),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_232),
.C(n_240),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_300),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_242),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_301),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_302),
.A2(n_266),
.B(n_275),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_252),
.C(n_251),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_273),
.C(n_272),
.Y(n_321)
);

XOR2x2_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_247),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_263),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_270),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_307),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_199),
.B1(n_169),
.B2(n_171),
.Y(n_308)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_285),
.A2(n_258),
.B1(n_266),
.B2(n_261),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_315),
.A2(n_328),
.B1(n_289),
.B2(n_300),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_290),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_317),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_318),
.B(n_320),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_284),
.B(n_273),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_326),
.C(n_293),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_292),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_322),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_303),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_305),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_299),
.C(n_293),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_327),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_285),
.A2(n_261),
.B1(n_256),
.B2(n_264),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_319),
.A2(n_291),
.B1(n_294),
.B2(n_302),
.Y(n_333)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_287),
.Y(n_334)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_334),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_323),
.A2(n_287),
.B1(n_295),
.B2(n_297),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

INVx3_ASAP7_75t_SL g336 ( 
.A(n_313),
.Y(n_336)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_310),
.Y(n_338)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_346),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_326),
.C(n_312),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_343),
.A2(n_350),
.B1(n_351),
.B2(n_325),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_345),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_305),
.C(n_274),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_329),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_349),
.Y(n_354)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_348),
.Y(n_357)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_330),
.A2(n_305),
.B1(n_306),
.B2(n_269),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_330),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_332),
.B(n_327),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_353),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_364),
.C(n_338),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g356 ( 
.A(n_343),
.B(n_315),
.CI(n_320),
.CON(n_356),
.SN(n_356)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_360),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_321),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_341),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_312),
.C(n_324),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_337),
.B(n_316),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_365),
.B(n_368),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_344),
.A2(n_328),
.B(n_331),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_370),
.B(n_374),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g371 ( 
.A(n_353),
.B(n_318),
.CI(n_334),
.CON(n_371),
.SN(n_371)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_371),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_368),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_372),
.B(n_379),
.C(n_382),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_367),
.A2(n_325),
.B1(n_339),
.B2(n_346),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_375),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_345),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_354),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_369),
.A2(n_358),
.B1(n_357),
.B2(n_363),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_376),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_369),
.A2(n_350),
.B1(n_336),
.B2(n_340),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_378),
.A2(n_280),
.B(n_356),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_348),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_267),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_381),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_377),
.A2(n_358),
.B(n_362),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_385),
.A2(n_392),
.B(n_390),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_377),
.A2(n_356),
.B1(n_359),
.B2(n_362),
.Y(n_386)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_386),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_383),
.A2(n_363),
.B1(n_359),
.B2(n_314),
.Y(n_388)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_388),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_389),
.B(n_390),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_371),
.A2(n_316),
.B1(n_364),
.B2(n_267),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_269),
.C(n_265),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_394),
.B(n_379),
.C(n_372),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_279),
.C(n_259),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_384),
.Y(n_398)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_398),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_393),
.A2(n_395),
.B(n_385),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_399),
.B(n_393),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_380),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_404),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_181),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_259),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_405),
.A2(n_134),
.B(n_132),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_402),
.A2(n_394),
.B1(n_391),
.B2(n_265),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_406),
.B(n_410),
.C(n_396),
.Y(n_412)
);

NAND2x1_ASAP7_75t_L g409 ( 
.A(n_403),
.B(n_279),
.Y(n_409)
);

OAI21xp33_ASAP7_75t_SL g414 ( 
.A1(n_409),
.A2(n_411),
.B(n_134),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_412),
.A2(n_413),
.B(n_410),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_408),
.A2(n_400),
.B(n_397),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_414),
.A2(n_415),
.B(n_407),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_416),
.B(n_417),
.C(n_411),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_409),
.C(n_132),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_419),
.B(n_6),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_6),
.Y(n_421)
);


endmodule