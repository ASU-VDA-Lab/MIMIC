module fake_jpeg_16036_n_85 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_85);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_85;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx3_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx3_ASAP7_75t_SL g18 ( 
.A(n_16),
.Y(n_18)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_21),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_0),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_23),
.B1(n_17),
.B2(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_30),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_23),
.A3(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_20),
.B1(n_19),
.B2(n_11),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_19),
.B1(n_12),
.B2(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_11),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_14),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_27),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_46),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_9),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_9),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_51),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_58),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_26),
.C(n_25),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_45),
.B1(n_41),
.B2(n_24),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_59),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_56),
.A2(n_24),
.B1(n_46),
.B2(n_12),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_64),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_24),
.B1(n_13),
.B2(n_3),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_58),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_13),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_66),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_62),
.A3(n_61),
.B1(n_59),
.B2(n_52),
.C1(n_60),
.C2(n_24),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_74),
.B(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_76),
.B(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_1),
.Y(n_77)
);

AOI322xp5_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_76),
.C2(n_75),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_82),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_78),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_2),
.Y(n_85)
);


endmodule