module fake_jpeg_27243_n_83 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_83);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_83;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx3_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_14),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_14),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_28),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_15),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_15),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_18),
.B(n_17),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_41),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_19),
.B1(n_24),
.B2(n_12),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_8),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_13),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_51),
.C(n_50),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_9),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_53),
.A2(n_9),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_12),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_60),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_43),
.B(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_39),
.C(n_11),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_39),
.Y(n_67)
);

AOI322xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_6),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_45),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_56),
.C(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_67),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_58),
.B1(n_45),
.B2(n_57),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_56),
.B1(n_24),
.B2(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_8),
.B(n_3),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_65),
.C(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_74),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_73),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_70),
.B1(n_71),
.B2(n_24),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_78),
.B(n_79),
.Y(n_80)
);

NAND4xp25_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_77),
.C(n_75),
.D(n_6),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_5),
.B(n_7),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_0),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_0),
.Y(n_83)
);


endmodule