module fake_jpeg_18208_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_43),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_26),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_30),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_27),
.B1(n_16),
.B2(n_21),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_48),
.B1(n_46),
.B2(n_44),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_27),
.B1(n_16),
.B2(n_20),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_53),
.A2(n_72),
.B1(n_31),
.B2(n_28),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_67),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_21),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_24),
.B1(n_19),
.B2(n_29),
.Y(n_103)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_37),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_18),
.C(n_37),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_42),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_38),
.A2(n_16),
.B1(n_20),
.B2(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_79),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_78),
.B(n_82),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_88),
.B1(n_93),
.B2(n_96),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_83),
.Y(n_128)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_54),
.A2(n_33),
.B1(n_32),
.B2(n_48),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_60),
.A2(n_33),
.B1(n_32),
.B2(n_34),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_41),
.B1(n_39),
.B2(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_112),
.Y(n_114)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_63),
.B1(n_69),
.B2(n_59),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_32),
.B1(n_33),
.B2(n_31),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_95),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_47),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_62),
.C(n_18),
.Y(n_129)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_58),
.B1(n_66),
.B2(n_52),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_56),
.B1(n_67),
.B2(n_51),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_100),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_46),
.B1(n_44),
.B2(n_34),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_101),
.A2(n_104),
.B1(n_109),
.B2(n_19),
.Y(n_146)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_107),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_105),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_52),
.A2(n_36),
.B1(n_23),
.B2(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_59),
.A2(n_36),
.B1(n_23),
.B2(n_29),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_37),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_22),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_56),
.A2(n_0),
.B(n_1),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_107),
.B1(n_89),
.B2(n_111),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_120),
.A2(n_126),
.B1(n_77),
.B2(n_94),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_146),
.B1(n_99),
.B2(n_103),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_62),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_132),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_57),
.B1(n_56),
.B2(n_62),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_103),
.C(n_77),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_22),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_13),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_141),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_80),
.A2(n_63),
.B1(n_69),
.B2(n_19),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_108),
.B1(n_106),
.B2(n_112),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_96),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_147),
.B(n_149),
.Y(n_152)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_145),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_22),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_147),
.Y(n_164)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_90),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_25),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_105),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_163),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_159),
.B1(n_161),
.B2(n_177),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_152),
.A2(n_3),
.B(n_5),
.Y(n_213)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_166),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_154),
.B(n_118),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_155),
.A2(n_119),
.B1(n_8),
.B2(n_9),
.Y(n_211)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_149),
.C(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_121),
.A2(n_106),
.B1(n_84),
.B2(n_73),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_92),
.C(n_24),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_18),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_182),
.B(n_128),
.Y(n_201)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_130),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_168),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_130),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_171),
.B1(n_175),
.B2(n_140),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_122),
.A2(n_75),
.B1(n_74),
.B2(n_35),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_25),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_35),
.B1(n_9),
.B2(n_12),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_121),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_180),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_35),
.B1(n_25),
.B2(n_18),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_179),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_18),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_114),
.B(n_35),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_127),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_140),
.B1(n_117),
.B2(n_135),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_0),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_200),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_152),
.A2(n_143),
.B1(n_128),
.B2(n_135),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_190),
.A2(n_197),
.B1(n_3),
.B2(n_5),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_208),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_148),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_194),
.B(n_213),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_143),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_195),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_198),
.C(n_175),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_126),
.C(n_133),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_5),
.Y(n_233)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_201),
.A2(n_165),
.B(n_182),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_203),
.B(n_209),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_157),
.B(n_134),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_205),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_158),
.B(n_117),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_145),
.B1(n_139),
.B2(n_138),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_212),
.B1(n_5),
.B2(n_7),
.Y(n_235)
);

AOI22x1_ASAP7_75t_L g208 ( 
.A1(n_155),
.A2(n_170),
.B1(n_171),
.B2(n_164),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_164),
.A2(n_118),
.B1(n_119),
.B2(n_4),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_180),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_12),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_214),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_227),
.C(n_204),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_163),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_229),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_241),
.B(n_201),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_173),
.B1(n_174),
.B2(n_160),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_231),
.B1(n_235),
.B2(n_212),
.Y(n_244)
);

A2O1A1O1Ixp25_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_165),
.B(n_173),
.C(n_166),
.D(n_153),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_210),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_169),
.C(n_12),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_193),
.B(n_6),
.Y(n_229)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_234),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_236),
.B(n_238),
.Y(n_258)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_185),
.B(n_7),
.C(n_13),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_237),
.B(n_14),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_186),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_189),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_187),
.B1(n_203),
.B2(n_207),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_249),
.B1(n_224),
.B2(n_239),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_244),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_246),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_261),
.B(n_225),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_194),
.C(n_205),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_253),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_221),
.A2(n_208),
.B1(n_207),
.B2(n_192),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_223),
.B(n_198),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_255),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_208),
.B(n_192),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_217),
.A2(n_222),
.B(n_221),
.Y(n_255)
);

AO22x2_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_191),
.B1(n_14),
.B2(n_15),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

XOR2x2_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_14),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_226),
.C(n_227),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_229),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_264),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_259),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_268),
.Y(n_293)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_226),
.C(n_220),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_270),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_228),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_250),
.B(n_230),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_279),
.Y(n_290)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_278),
.B1(n_249),
.B2(n_235),
.Y(n_283)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_215),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_217),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_260),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_254),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_216),
.C(n_234),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_262),
.C(n_245),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_287),
.C(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_284),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_250),
.C(n_257),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_244),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_291),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_260),
.C(n_251),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_274),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_260),
.C(n_251),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_297),
.B(n_302),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_288),
.B1(n_272),
.B2(n_292),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_298),
.A2(n_301),
.B1(n_299),
.B2(n_302),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_271),
.B1(n_266),
.B2(n_264),
.Y(n_299)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_282),
.B1(n_286),
.B2(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_232),
.C(n_294),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_290),
.C(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_308),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_298),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_310),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_303),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_300),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_306),
.B(n_309),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_311),
.B(n_296),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_317),
.B(n_296),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_321),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_323),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_322),
.B(n_315),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_318),
.C(n_307),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_308),
.Y(n_329)
);


endmodule