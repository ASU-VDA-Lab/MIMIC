module fake_aes_4033_n_31 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_31);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_2), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
OAI22xp5_ASAP7_75t_L g14 ( .A1(n_1), .A2(n_0), .B1(n_8), .B2(n_4), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_1), .B(n_3), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_13), .B(n_2), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_13), .B(n_15), .Y(n_19) );
BUFx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
INVxp67_ASAP7_75t_SL g22 ( .A(n_21), .Y(n_22) );
HB1xp67_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
AOI221xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_20), .B1(n_22), .B2(n_14), .C(n_17), .Y(n_24) );
INVxp67_ASAP7_75t_SL g25 ( .A(n_24), .Y(n_25) );
AOI221xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_17), .B1(n_16), .B2(n_12), .C(n_4), .Y(n_26) );
NAND4xp75_ASAP7_75t_L g27 ( .A(n_26), .B(n_16), .C(n_5), .D(n_7), .Y(n_27) );
INVx5_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
BUFx3_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
OAI22xp5_ASAP7_75t_SL g30 ( .A1(n_29), .A2(n_28), .B1(n_27), .B2(n_10), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_29), .B1(n_9), .B2(n_11), .Y(n_31) );
endmodule