module fake_jpeg_9399_n_286 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

NAND2x1_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_29),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_54),
.B(n_18),
.C(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_53),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_22),
.B1(n_30),
.B2(n_29),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_29),
.B1(n_22),
.B2(n_30),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_40),
.B1(n_39),
.B2(n_19),
.Y(n_79)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_60),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_22),
.B(n_16),
.C(n_21),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_31),
.B1(n_16),
.B2(n_21),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_25),
.B1(n_32),
.B2(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_28),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_64),
.B(n_32),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_28),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_71),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_26),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_79),
.B1(n_83),
.B2(n_86),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_37),
.C(n_41),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_57),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_85),
.B1(n_56),
.B2(n_25),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_53),
.B(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_45),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_89),
.Y(n_105)
);

AO22x2_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_26),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_0),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_25),
.Y(n_100)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_95),
.Y(n_140)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_94),
.B(n_102),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_101),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_49),
.B1(n_59),
.B2(n_46),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_85),
.B1(n_67),
.B2(n_49),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_111),
.Y(n_119)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_103),
.B(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_56),
.B(n_24),
.C(n_27),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_85),
.B(n_63),
.C(n_80),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_114),
.B1(n_116),
.B2(n_85),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_57),
.C(n_43),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_111),
.C(n_73),
.Y(n_125)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_116),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

AOI22x1_ASAP7_75t_SL g117 ( 
.A1(n_115),
.A2(n_85),
.B1(n_70),
.B2(n_83),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_126),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_142),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_127),
.B(n_11),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_145),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_112),
.B(n_71),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_134),
.B(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_63),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_139),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_83),
.B1(n_72),
.B2(n_85),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_138),
.B1(n_144),
.B2(n_121),
.Y(n_146)
);

BUFx12f_ASAP7_75t_SL g134 ( 
.A(n_100),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_94),
.A2(n_58),
.B1(n_49),
.B2(n_67),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_46),
.B1(n_88),
.B2(n_68),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_109),
.B(n_64),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_90),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_98),
.A2(n_68),
.B1(n_84),
.B2(n_90),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_155),
.B1(n_162),
.B2(n_168),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_93),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_147),
.A2(n_164),
.B(n_165),
.Y(n_179)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_107),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_151),
.A2(n_153),
.B1(n_160),
.B2(n_166),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_140),
.Y(n_153)
);

AOI22x1_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_100),
.B1(n_90),
.B2(n_102),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_64),
.Y(n_156)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_97),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_123),
.A2(n_101),
.B1(n_91),
.B2(n_68),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_76),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_145),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

AO22x1_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_57),
.B1(n_43),
.B2(n_26),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_89),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_170),
.A2(n_130),
.B1(n_12),
.B2(n_10),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_175),
.B(n_156),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_33),
.B1(n_27),
.B2(n_24),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_33),
.B1(n_23),
.B2(n_8),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_106),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_174),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_110),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_129),
.B(n_1),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_157),
.A2(n_125),
.B1(n_138),
.B2(n_126),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_178),
.B1(n_191),
.B2(n_193),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_170),
.A2(n_136),
.B1(n_119),
.B2(n_142),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_119),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_194),
.C(n_175),
.Y(n_212)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_9),
.B(n_15),
.C(n_14),
.D(n_13),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_186),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_168),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_196),
.B(n_175),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_174),
.B(n_147),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_130),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_168),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_3),
.C(n_4),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_195),
.B(n_171),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_152),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_164),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_166),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

OR2x4_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_155),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_218),
.B(n_220),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_208),
.A2(n_211),
.B1(n_213),
.B2(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_148),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_183),
.C(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_161),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_154),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_217),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_162),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_192),
.B(n_172),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_151),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_221),
.A2(n_222),
.B(n_152),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_203),
.B(n_202),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_222),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_179),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_200),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_177),
.B1(n_178),
.B2(n_199),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_232),
.B1(n_198),
.B2(n_154),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_199),
.B1(n_193),
.B2(n_180),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_208),
.C(n_207),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_235),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_215),
.C(n_214),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_219),
.A2(n_180),
.B1(n_149),
.B2(n_187),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_201),
.B1(n_155),
.B2(n_147),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_220),
.B1(n_219),
.B2(n_218),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_209),
.B(n_201),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_248),
.B(n_224),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_227),
.C(n_233),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_247),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_223),
.B(n_153),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_246),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_244),
.A2(n_232),
.B1(n_234),
.B2(n_226),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_210),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_204),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_224),
.B(n_230),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_250),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_249),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_5),
.C(n_6),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_228),
.C(n_225),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_158),
.C(n_5),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_257),
.Y(n_270)
);

XNOR2x1_ASAP7_75t_SL g258 ( 
.A(n_251),
.B(n_229),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_259),
.B1(n_244),
.B2(n_241),
.Y(n_265)
);

AO221x1_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_182),
.B1(n_231),
.B2(n_238),
.C(n_185),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_250),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_263),
.B(n_264),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_186),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_262),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_269),
.C(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_253),
.B(n_4),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_5),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_273),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_258),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_252),
.B1(n_257),
.B2(n_254),
.Y(n_275)
);

NOR2x1_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_6),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_252),
.B(n_266),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_280),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_273),
.B(n_274),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_281),
.A2(n_279),
.B(n_277),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_270),
.C(n_282),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_284),
.A2(n_270),
.B(n_6),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_7),
.Y(n_286)
);


endmodule