module fake_jpeg_4333_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_0),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_22),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_25),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_28),
.B1(n_15),
.B2(n_24),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_51),
.B1(n_26),
.B2(n_16),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_28),
.B1(n_24),
.B2(n_17),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_17),
.B1(n_24),
.B2(n_18),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_52),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_28),
.B1(n_27),
.B2(n_18),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_59),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_56),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_38),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_38),
.C(n_39),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_30),
.B(n_39),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_37),
.B1(n_40),
.B2(n_36),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_73),
.B1(n_47),
.B2(n_21),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_27),
.B(n_37),
.C(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_78),
.B(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_42),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_55),
.B1(n_59),
.B2(n_47),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_87),
.B1(n_89),
.B2(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_36),
.B1(n_40),
.B2(n_39),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_52),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_78),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_30),
.C(n_74),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_26),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_36),
.B1(n_40),
.B2(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_106),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_65),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_105),
.B(n_100),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_72),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_99),
.C(n_105),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_103),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_64),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_61),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_81),
.B(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_86),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_87),
.C(n_84),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_109),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_50),
.B(n_62),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_60),
.B(n_45),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_117),
.B(n_29),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_87),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_104),
.B1(n_98),
.B2(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_129),
.B1(n_130),
.B2(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_126),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_61),
.B1(n_63),
.B2(n_77),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_125),
.B1(n_29),
.B2(n_23),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_85),
.B1(n_82),
.B2(n_60),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_128),
.A2(n_21),
.B(n_22),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_70),
.B1(n_90),
.B2(n_58),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_97),
.B1(n_101),
.B2(n_70),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_101),
.C(n_22),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_136),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_113),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_35),
.C(n_56),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_134),
.C(n_142),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_35),
.C(n_88),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_129),
.A2(n_29),
.B1(n_26),
.B2(n_23),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_137),
.B(n_138),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_145),
.B1(n_114),
.B2(n_122),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_146),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_22),
.C(n_23),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_127),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_21),
.B1(n_16),
.B2(n_20),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_149),
.C(n_158),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_118),
.C(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_130),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_19),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_121),
.B(n_120),
.C(n_119),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_117),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_156),
.B(n_20),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_114),
.C(n_124),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_125),
.C(n_22),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_19),
.C(n_3),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_139),
.B(n_145),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_2),
.B(n_4),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_140),
.B1(n_142),
.B2(n_20),
.Y(n_163)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_160),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_168),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_20),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_5),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_19),
.B(n_3),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_2),
.B(n_3),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_172),
.A2(n_148),
.B(n_151),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_166),
.C(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_157),
.B(n_153),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_179),
.B(n_172),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_19),
.B1(n_4),
.B2(n_5),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_181),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_183),
.B(n_187),
.Y(n_190)
);

AOI31xp33_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_161),
.A3(n_165),
.B(n_170),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_188),
.C(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_171),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_168),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_191),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_175),
.C(n_176),
.Y(n_191)
);

OAI21x1_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_14),
.B(n_7),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_6),
.C(n_7),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_9),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_186),
.A2(n_8),
.B(n_9),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_194),
.A2(n_9),
.B(n_10),
.Y(n_197)
);

OAI321xp33_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_190),
.A3(n_185),
.B1(n_12),
.B2(n_13),
.C(n_11),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_198),
.A2(n_10),
.B(n_11),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_200),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_SL g202 ( 
.A(n_199),
.B(n_195),
.C(n_196),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_202),
.A2(n_201),
.B(n_10),
.Y(n_203)
);


endmodule