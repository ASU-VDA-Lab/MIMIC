module real_jpeg_15133_n_3 (n_1, n_0, n_2, n_3);

input n_1;
input n_0;
input n_2;

output n_3;

wire n_5;
wire n_4;
wire n_8;
wire n_11;
wire n_6;
wire n_7;
wire n_10;
wire n_9;

INVx2_ASAP7_75t_R g6 ( 
.A(n_0),
.Y(n_6)
);

OA22x2_ASAP7_75t_L g8 ( 
.A1(n_1),
.A2(n_2),
.B1(n_9),
.B2(n_10),
.Y(n_8)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g3 ( 
.A(n_4),
.B(n_11),
.Y(n_3)
);

INVx1_ASAP7_75t_L g4 ( 
.A(n_5),
.Y(n_4)
);

NOR2xp33_ASAP7_75t_L g5 ( 
.A(n_6),
.B(n_7),
.Y(n_5)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_6),
.B(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_SL g7 ( 
.A(n_8),
.Y(n_7)
);


endmodule