module fake_jpeg_21414_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_4),
.B(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_21),
.B1(n_15),
.B2(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_20),
.A2(n_26),
.B(n_17),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_24),
.Y(n_29)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_1),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_4),
.B1(n_10),
.B2(n_9),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_15),
.B1(n_26),
.B2(n_23),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_8),
.B(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_21),
.A2(n_16),
.B(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.C(n_29),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_34),
.B1(n_27),
.B2(n_28),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.C(n_37),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NOR3xp33_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_38),
.C(n_39),
.Y(n_46)
);


endmodule