module fake_jpeg_7690_n_235 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_235);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_235;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_32),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_59),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_18),
.B1(n_31),
.B2(n_26),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_46),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_24),
.B(n_23),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_58),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_64),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_33),
.A2(n_18),
.B1(n_31),
.B2(n_26),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g81 ( 
.A(n_53),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_18),
.B1(n_31),
.B2(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_60),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_22),
.B1(n_32),
.B2(n_17),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_22),
.B1(n_21),
.B2(n_23),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_22),
.B1(n_24),
.B2(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_30),
.B1(n_17),
.B2(n_25),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_65),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_30),
.B1(n_27),
.B2(n_25),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_0),
.C(n_2),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_19),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_68),
.B(n_79),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_77),
.Y(n_106)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_37),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_50),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_98),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_48),
.C(n_35),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_36),
.C(n_42),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_52),
.B1(n_27),
.B2(n_19),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_93),
.B1(n_102),
.B2(n_42),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_43),
.B1(n_67),
.B2(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_45),
.Y(n_98)
);

AOI32xp33_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_54),
.A3(n_45),
.B1(n_47),
.B2(n_65),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_85),
.B(n_88),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_82),
.B1(n_85),
.B2(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_50),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_59),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

BUFx4f_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_125),
.B1(n_99),
.B2(n_36),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_117),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_116),
.B(n_38),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_73),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_124),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_111),
.B1(n_110),
.B2(n_102),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_129),
.B1(n_104),
.B2(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_43),
.B1(n_88),
.B2(n_54),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_88),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_132),
.C(n_101),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_74),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_128),
.Y(n_148)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_56),
.B1(n_67),
.B2(n_76),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_133),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_52),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_110),
.B(n_98),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_152),
.B(n_154),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_149),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_143),
.B(n_146),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_95),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_142),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_124),
.B1(n_119),
.B2(n_125),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_105),
.B1(n_104),
.B2(n_44),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_89),
.Y(n_142)
);

AO21x1_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_107),
.B(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_51),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_155),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_147),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_106),
.B(n_97),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_42),
.C(n_38),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_44),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_38),
.C(n_39),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_34),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_161),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_112),
.B1(n_117),
.B2(n_128),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_168),
.B1(n_171),
.B2(n_104),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_63),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_164),
.B(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_44),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_141),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_166),
.A2(n_172),
.B1(n_173),
.B2(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_105),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_155),
.C(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_176),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_145),
.C(n_154),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_179),
.C(n_182),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_140),
.B1(n_138),
.B2(n_152),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_167),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_147),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_181),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_34),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_34),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_38),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_164),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_83),
.C(n_77),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_189),
.C(n_165),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_2),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_185),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_160),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_195),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_197),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_162),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_202),
.C(n_203),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_156),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_200),
.B(n_188),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_204),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_201),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_206),
.A2(n_210),
.B(n_211),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_190),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_203),
.C(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_185),
.Y(n_210)
);

NAND4xp25_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_181),
.C(n_183),
.D(n_14),
.Y(n_211)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_214),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_210),
.A2(n_156),
.B1(n_194),
.B2(n_13),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_219),
.C(n_208),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_205),
.A2(n_194),
.B(n_4),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_14),
.B(n_15),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_12),
.C(n_15),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_222),
.Y(n_226)
);

NOR2xp67_ASAP7_75t_SL g221 ( 
.A(n_216),
.B(n_207),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_221),
.A2(n_223),
.B(n_218),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_217),
.B(n_207),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_227),
.C(n_228),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_213),
.B(n_87),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_13),
.C(n_39),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_44),
.Y(n_229)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_39),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_231),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_230),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_232),
.C(n_7),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_6),
.B(n_8),
.Y(n_235)
);


endmodule