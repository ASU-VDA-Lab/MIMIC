module fake_jpeg_31323_n_69 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_32;
wire n_66;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_7),
.B(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_40),
.B1(n_45),
.B2(n_48),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_43),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_24),
.A2(n_6),
.B1(n_9),
.B2(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_6),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_26),
.B1(n_35),
.B2(n_21),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_26),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_35),
.B1(n_25),
.B2(n_23),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_58),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_49),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_51),
.C(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_55),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_28),
.Y(n_62)
);

AOI21x1_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_57),
.B(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_60),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_63),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_66),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_66),
.C(n_64),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_40),
.B(n_29),
.Y(n_69)
);


endmodule