module fake_ariane_1527_n_105 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_17, n_4, n_10, n_105);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_17;
input n_4;
input n_10;

output n_105;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_18;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_87;
wire n_81;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVxp67_ASAP7_75t_SL g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVxp67_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_0),
.Y(n_37)
);

AND2x6_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_6),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

AND2x4_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_23),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_20),
.C(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_52),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_34),
.B1(n_43),
.B2(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_50),
.B1(n_38),
.B2(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_56),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_54),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_48),
.B1(n_47),
.B2(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_61),
.B(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_73)
);

AOI221xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_66),
.B1(n_36),
.B2(n_40),
.C(n_18),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_36),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_38),
.B1(n_61),
.B2(n_59),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_4),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_45),
.Y(n_80)
);

OAI31xp33_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_38),
.A3(n_4),
.B(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_78),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_85),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

OAI31xp33_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_87),
.A3(n_83),
.B(n_81),
.Y(n_94)
);

NOR2xp67_ASAP7_75t_SL g95 ( 
.A(n_93),
.B(n_88),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_94),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_91),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

AOI31xp33_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_78),
.A3(n_80),
.B(n_13),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_51),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

OAI221xp5_ASAP7_75t_R g102 ( 
.A1(n_101),
.A2(n_99),
.B1(n_12),
.B2(n_16),
.C(n_17),
.Y(n_102)
);

OR3x2_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_8),
.C(n_38),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_49),
.B(n_51),
.Y(n_105)
);


endmodule