module fake_jpeg_1475_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_56),
.Y(n_71)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_53),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_1),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_53),
.B(n_51),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_58),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_54),
.C(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_81),
.Y(n_99)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_55),
.B1(n_65),
.B2(n_43),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_62),
.B1(n_63),
.B2(n_41),
.Y(n_87)
);

NAND2x1p5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_56),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_64),
.Y(n_86)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_38),
.B(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_59),
.B1(n_48),
.B2(n_42),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_84),
.B1(n_45),
.B2(n_52),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_42),
.B1(n_48),
.B2(n_40),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_39),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_2),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_83),
.B(n_9),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_97),
.B(n_96),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_45),
.B1(n_40),
.B2(n_52),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_98),
.B1(n_101),
.B2(n_7),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_47),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_47),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_39),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_96),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_38),
.B1(n_44),
.B2(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_83),
.B1(n_74),
.B2(n_6),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_37),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_36),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_105),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_114),
.B1(n_116),
.B2(n_15),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_4),
.C(n_5),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_112),
.B1(n_117),
.B2(n_83),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_7),
.CI(n_9),
.CON(n_109),
.SN(n_109)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_113),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_21),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_111),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_92),
.B1(n_99),
.B2(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_10),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_10),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_120)
);

OAI22x1_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_131),
.B1(n_103),
.B2(n_110),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_129),
.B1(n_123),
.B2(n_125),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_24),
.C(n_30),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_130),
.B(n_127),
.C(n_128),
.D(n_124),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_14),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_16),
.C(n_17),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_108),
.C(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_R g132 ( 
.A(n_130),
.B(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_134),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_136),
.B(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_125),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_123),
.C(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_136),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_143),
.Y(n_144)
);

AOI21x1_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_139),
.B(n_140),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_138),
.C(n_120),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_121),
.B1(n_126),
.B2(n_25),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_34),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_18),
.Y(n_150)
);


endmodule