module fake_jpeg_32165_n_146 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_146);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_34),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_31),
.A2(n_3),
.B(n_4),
.Y(n_55)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_5),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_19),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_21),
.C(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_67),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_4),
.B(n_8),
.Y(n_74)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_64),
.Y(n_83)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_29),
.B1(n_28),
.B2(n_24),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_42),
.B1(n_19),
.B2(n_44),
.Y(n_70)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_13),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_22),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_31),
.B(n_27),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_26),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_74),
.B1(n_80),
.B2(n_49),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_77),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_32),
.B1(n_24),
.B2(n_21),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_75),
.B1(n_81),
.B2(n_83),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_32),
.B1(n_14),
.B2(n_27),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_12),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_48),
.B1(n_56),
.B2(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_23),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_86),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_26),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_61),
.B(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_8),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_12),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_103),
.C(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_97),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_74),
.B1(n_86),
.B2(n_75),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_49),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_82),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_50),
.C(n_78),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_93),
.C(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_50),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_104),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_82),
.B(n_76),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_90),
.B(n_94),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_76),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_95),
.C(n_102),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_127),
.B(n_131),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_114),
.C(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_136),
.Y(n_139)
);

OA21x2_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_126),
.B(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_137),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_128),
.A2(n_126),
.B1(n_111),
.B2(n_121),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_111),
.B1(n_115),
.B2(n_100),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_131),
.B(n_127),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_138),
.A2(n_134),
.B(n_136),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_135),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_139),
.C(n_142),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_137),
.C(n_98),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_99),
.Y(n_146)
);


endmodule