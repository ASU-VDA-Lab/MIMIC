module fake_jpeg_1093_n_127 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_55),
.Y(n_62)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_0),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_2),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_39),
.B1(n_48),
.B2(n_38),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_35),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_67),
.Y(n_71)
);

BUFx2_ASAP7_75t_SL g66 ( 
.A(n_50),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_47),
.B(n_3),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_6),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_51),
.B1(n_50),
.B2(n_40),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_75),
.B1(n_58),
.B2(n_42),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_79),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_49),
.C(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_76),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_51),
.B1(n_40),
.B2(n_43),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_20),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_35),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_43),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_94)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_54),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_6),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_7),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_100),
.B1(n_32),
.B2(n_34),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_104),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_100)
);

XNOR2x1_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_16),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_19),
.B(n_23),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_105),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_24),
.C(n_26),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_29),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_111),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_106),
.B(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_31),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_116),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_102),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_120),
.A2(n_121),
.B1(n_113),
.B2(n_109),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_113),
.B(n_95),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_119),
.C(n_101),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_108),
.C(n_98),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_99),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_117),
.Y(n_127)
);


endmodule