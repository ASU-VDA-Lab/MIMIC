module real_jpeg_31199_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_0),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_0),
.Y(n_176)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_0),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_0),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_1),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_1),
.B(n_482),
.Y(n_481)
);

OAI22x1_ASAP7_75t_SL g52 ( 
.A1(n_2),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_2),
.Y(n_58)
);

AO22x1_ASAP7_75t_SL g180 ( 
.A1(n_2),
.A2(n_32),
.B1(n_58),
.B2(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_2),
.A2(n_58),
.B1(n_71),
.B2(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_2),
.B(n_111),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_SL g406 ( 
.A(n_2),
.B(n_401),
.Y(n_406)
);

OAI32xp33_ASAP7_75t_L g421 ( 
.A1(n_2),
.A2(n_422),
.A3(n_424),
.B1(n_427),
.B2(n_431),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_3),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_3),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_3),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_4),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_4),
.Y(n_101)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_5),
.Y(n_181)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_5),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_6),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_6),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_6),
.A2(n_203),
.B1(n_300),
.B2(n_302),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_6),
.A2(n_203),
.B1(n_379),
.B2(n_382),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_6),
.A2(n_203),
.B1(n_391),
.B2(n_393),
.Y(n_390)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_7),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_8),
.A2(n_65),
.B1(n_70),
.B2(n_74),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_8),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_8),
.A2(n_59),
.B1(n_74),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_8),
.A2(n_74),
.B1(n_255),
.B2(n_258),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_9),
.Y(n_94)
);

AO22x2_ASAP7_75t_SL g104 ( 
.A1(n_10),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_10),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_10),
.A2(n_109),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_10),
.A2(n_109),
.B1(n_160),
.B2(n_163),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_10),
.A2(n_109),
.B1(n_225),
.B2(n_228),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_11),
.Y(n_118)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_12),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_13),
.Y(n_88)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_13),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_479),
.B(n_481),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_236),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_235),
.Y(n_16)
);

INVxp33_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_195),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_19),
.B(n_195),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_166),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_150),
.B2(n_165),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_112),
.Y(n_22)
);

XNOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_63),
.Y(n_23)
);

MAJx2_ASAP7_75t_L g329 ( 
.A(n_24),
.B(n_330),
.C(n_332),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_24),
.A2(n_25),
.B1(n_330),
.B2(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_42),
.B(n_52),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_26),
.B(n_52),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_26),
.B(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_26),
.B(n_378),
.Y(n_409)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_27),
.B(n_58),
.Y(n_449)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_28),
.B(n_159),
.Y(n_192)
);

OAI22x1_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_35),
.B2(n_39),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_34),
.Y(n_178)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_41),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_41),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_42),
.B(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_42),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_42),
.B(n_52),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_42),
.B(n_378),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_46),
.Y(n_51)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_57),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_58),
.A2(n_134),
.B(n_137),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_58),
.B(n_138),
.Y(n_137)
);

NOR2xp67_ASAP7_75t_SL g346 ( 
.A(n_58),
.B(n_149),
.Y(n_346)
);

AOI32xp33_ASAP7_75t_L g399 ( 
.A1(n_58),
.A2(n_400),
.A3(n_402),
.B1(n_405),
.B2(n_406),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_58),
.B(n_428),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_58),
.B(n_168),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_62),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_75),
.B(n_102),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_69),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2x1_ASAP7_75t_L g155 ( 
.A(n_76),
.B(n_104),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_76),
.B(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g210 ( 
.A(n_77),
.B(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_77),
.A2(n_211),
.B(n_251),
.Y(n_250)
);

AO21x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_85),
.B(n_91),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_80),
.Y(n_278)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_85),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_87),
.Y(n_301)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_91)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_93),
.Y(n_433)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_102),
.B(n_298),
.Y(n_345)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g209 ( 
.A(n_103),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_111),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_106),
.Y(n_292)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_107),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_111),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_111),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_111),
.B(n_299),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_141),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_114),
.B(n_249),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_133),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_115),
.A2(n_116),
.B(n_133),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_115),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_115),
.B(n_142),
.Y(n_248)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_123),
.Y(n_115)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_L g249 ( 
.A(n_116),
.B(n_200),
.Y(n_249)
);

AO22x2_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_118),
.Y(n_281)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_128),
.B2(n_130),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_132),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_133),
.B(n_148),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_136),
.Y(n_206)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_136),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_137),
.Y(n_293)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_141),
.B(n_199),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_151),
.A2(n_152),
.B(n_156),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_155),
.B(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_157),
.B(n_377),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_158),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_158),
.B(n_216),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_158),
.B(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_162),
.Y(n_426)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_182),
.B(n_193),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_167),
.B(n_194),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_167),
.A2(n_184),
.B1(n_185),
.B2(n_312),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_167),
.A2(n_184),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_167),
.B(n_399),
.Y(n_470)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_173),
.B(n_179),
.Y(n_167)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_173),
.A2(n_254),
.B(n_261),
.Y(n_253)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_174),
.B(n_180),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_174),
.B(n_390),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_175),
.Y(n_262)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_178),
.Y(n_257)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_181),
.Y(n_260)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_181),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_181),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_182),
.A2(n_183),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_185),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_191),
.B(n_192),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_190),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_190),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_192),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_192),
.B(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_230),
.C(n_231),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_196),
.B(n_365),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_208),
.C(n_215),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_198),
.B(n_209),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_210),
.Y(n_412)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_211),
.Y(n_297)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_215),
.B(n_310),
.Y(n_309)
);

XNOR2x2_ASAP7_75t_SL g267 ( 
.A(n_217),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_218),
.B(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_223),
.A2(n_254),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_223),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_224),
.B(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_227),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_227),
.Y(n_395)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_230),
.Y(n_366)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2x1p5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_367),
.Y(n_237)
);

OAI21x1_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_320),
.B(n_357),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_306),
.Y(n_239)
);

INVxp33_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

AOI21x1_ASAP7_75t_L g355 ( 
.A1(n_241),
.A2(n_319),
.B(n_356),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_266),
.C(n_269),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_244),
.B(n_267),
.Y(n_337)
);

OAI22x1_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_252),
.B2(n_265),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2x2_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_247),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_250),
.Y(n_316)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_252),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_263),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_253),
.B(n_263),
.Y(n_334)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g348 ( 
.A(n_261),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_261),
.B(n_389),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_264),
.B(n_409),
.Y(n_440)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVxp33_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_270),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_294),
.C(n_304),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_271),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_272),
.B(n_275),
.Y(n_343)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_274),
.Y(n_445)
);

OAI31xp33_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_279),
.A3(n_282),
.B(n_286),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx4f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_291),
.B(n_293),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_295),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_304),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_305),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_313),
.B(n_319),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_308),
.B(n_313),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_313),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_314),
.B(n_360),
.C(n_362),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.C(n_317),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_352),
.B(n_355),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_338),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_322),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_335),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_323),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.C(n_333),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_351),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_334),
.Y(n_351)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_331),
.B(n_412),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_341),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_335),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_350),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_350),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.C(n_344),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_340),
.B(n_474),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_343),
.B(n_344),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.C(n_347),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_345),
.B(n_466),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_346),
.A2(n_347),
.B1(n_348),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_346),
.Y(n_467)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_349),
.B(n_444),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_355),
.A2(n_358),
.B(n_363),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_363),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_359),
.B(n_364),
.Y(n_478)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AOI31xp67_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_370),
.A3(n_477),
.B(n_478),
.Y(n_367)
);

OAI21x1_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_472),
.B(n_476),
.Y(n_370)
);

AOI21x1_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_461),
.B(n_471),
.Y(n_371)
);

AO21x1_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_414),
.B(n_460),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_396),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_374),
.B(n_396),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_385),
.C(n_387),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_376),
.A2(n_385),
.B1(n_386),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_390),
.B(n_445),
.Y(n_444)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_407),
.Y(n_396)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_397),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_408),
.A2(n_410),
.B1(n_411),
.B2(n_413),
.Y(n_407)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_408),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_410),
.B(n_413),
.C(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_415),
.A2(n_441),
.B(n_459),
.Y(n_414)
);

NOR2x1_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_419),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_416),
.B(n_419),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_439),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_420),
.A2(n_421),
.B1(n_439),
.B2(n_440),
.Y(n_446)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_436),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_442),
.A2(n_447),
.B(n_458),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_446),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_446),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_448),
.A2(n_451),
.B(n_457),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_450),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_456),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_464),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_464),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_468),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_465),
.B(n_469),
.C(n_470),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_475),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_473),
.B(n_475),
.Y(n_476)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);


endmodule