module fake_ibex_1313_n_762 (n_85, n_128, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_55, n_130, n_63, n_98, n_129, n_29, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_112, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_101, n_113, n_96, n_68, n_117, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_762);

input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_101;
input n_113;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_762;

wire n_151;
wire n_599;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_638;
wire n_398;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_421;
wire n_738;
wire n_475;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_375;
wire n_317;
wire n_340;
wire n_708;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_170;
wire n_144;
wire n_270;
wire n_383;
wire n_346;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_750;
wire n_746;
wire n_136;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_474;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_141;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_689;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_618;
wire n_488;
wire n_139;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_137;
wire n_679;
wire n_338;
wire n_173;
wire n_696;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_718;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_567;
wire n_516;
wire n_548;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_444;
wire n_200;
wire n_562;
wire n_506;
wire n_564;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_410;
wire n_308;
wire n_675;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_135;
wire n_520;
wire n_684;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_138;
wire n_650;
wire n_409;
wire n_582;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_728;
wire n_670;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_752;
wire n_668;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_202;
wire n_231;
wire n_298;
wire n_159;
wire n_587;
wire n_760;
wire n_751;
wire n_160;
wire n_657;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_1),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_36),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_108),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_15),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_99),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_100),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_41),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_79),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_12),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_14),
.Y(n_145)
);

BUFx10_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_34),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_85),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_32),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_114),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_98),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_56),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_29),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_89),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_57),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_7),
.Y(n_161)
);

NOR2xp67_ASAP7_75t_L g162 ( 
.A(n_24),
.B(n_42),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_12),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_23),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_13),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_14),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_40),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_29),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_92),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_64),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_44),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_103),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_39),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_69),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_68),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_47),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_9),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_63),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_59),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_61),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_19),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_37),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_66),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_35),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_17),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_82),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_6),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_1),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_91),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_84),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_73),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_58),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_70),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_118),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_52),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_104),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_43),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_38),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_109),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_28),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_78),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_81),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_112),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_86),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_49),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_45),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_54),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_5),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_94),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_33),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_90),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_31),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_17),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_83),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_62),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_152),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_0),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_152),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_136),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_132),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_234)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_2),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_152),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_138),
.A2(n_199),
.B1(n_222),
.B2(n_158),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_134),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_133),
.Y(n_241)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_3),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_147),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_146),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_152),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_147),
.Y(n_248)
);

BUFx8_ASAP7_75t_SL g249 ( 
.A(n_161),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_164),
.B(n_4),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_171),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_145),
.B(n_5),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g254 ( 
.A1(n_186),
.A2(n_74),
.B(n_131),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_134),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_168),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g257 ( 
.A1(n_186),
.A2(n_210),
.B(n_188),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_170),
.Y(n_258)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_171),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_6),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_135),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_205),
.B(n_8),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_171),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_144),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_166),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_134),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_181),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_205),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_171),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_134),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_184),
.A2(n_11),
.B1(n_15),
.B2(n_16),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_134),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_181),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_134),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_188),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g277 ( 
.A(n_187),
.B(n_16),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_187),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_148),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_195),
.B(n_18),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_195),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_191),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_192),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_150),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_156),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_157),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_163),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_191),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_226),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_213),
.A2(n_165),
.B1(n_198),
.B2(n_220),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_169),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_173),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_175),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_177),
.Y(n_295)
);

OA21x2_ASAP7_75t_L g296 ( 
.A1(n_178),
.A2(n_80),
.B(n_130),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_179),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_180),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_183),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_191),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_242),
.B(n_167),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_231),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_231),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_235),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_277),
.B(n_185),
.Y(n_309)
);

OR2x6_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_162),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_235),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_277),
.B(n_189),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_267),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_280),
.B(n_241),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_230),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_235),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_267),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_253),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_280),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_245),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_273),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_L g325 ( 
.A1(n_238),
.A2(n_137),
.B1(n_174),
.B2(n_212),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_241),
.B(n_193),
.Y(n_326)
);

BUFx10_ASAP7_75t_L g327 ( 
.A(n_259),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_230),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_275),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_244),
.Y(n_331)
);

AO22x2_ASAP7_75t_L g332 ( 
.A1(n_272),
.A2(n_229),
.B1(n_224),
.B2(n_200),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_249),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_275),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_257),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_257),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_248),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_SL g338 ( 
.A(n_263),
.B(n_214),
.Y(n_338)
);

NAND2xp33_ASAP7_75t_L g339 ( 
.A(n_263),
.B(n_191),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_257),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_276),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_276),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_262),
.B(n_201),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_256),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_233),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_230),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_232),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_258),
.Y(n_349)
);

AOI21x1_ASAP7_75t_L g350 ( 
.A1(n_254),
.A2(n_203),
.B(n_211),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_281),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_245),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_248),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_232),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_259),
.B(n_204),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_259),
.B(n_206),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_266),
.B(n_215),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_281),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_265),
.B(n_139),
.Y(n_359)
);

AO21x2_ASAP7_75t_L g360 ( 
.A1(n_254),
.A2(n_218),
.B(n_217),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_234),
.A2(n_219),
.B1(n_227),
.B2(n_225),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_236),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_244),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_236),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_279),
.A2(n_172),
.B1(n_143),
.B2(n_182),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_252),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_252),
.Y(n_367)
);

CKINVDCx6p67_ASAP7_75t_R g368 ( 
.A(n_251),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_249),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_252),
.Y(n_370)
);

INVx8_ASAP7_75t_L g371 ( 
.A(n_233),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_252),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_252),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_298),
.B(n_140),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_284),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_285),
.B(n_141),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_260),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_260),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_290),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_274),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_278),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_286),
.Y(n_382)
);

CKINVDCx6p67_ASAP7_75t_R g383 ( 
.A(n_278),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_337),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_305),
.A2(n_287),
.B1(n_292),
.B2(n_297),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_337),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_315),
.A2(n_296),
.B(n_243),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_344),
.B(n_376),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_341),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_305),
.A2(n_299),
.B1(n_295),
.B2(n_294),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_335),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_301),
.A2(n_286),
.B1(n_291),
.B2(n_294),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_304),
.A2(n_291),
.B1(n_250),
.B2(n_261),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_268),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_307),
.A2(n_237),
.B1(n_239),
.B2(n_268),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_344),
.B(n_374),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_345),
.B(n_239),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_375),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_382),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_319),
.B(n_239),
.Y(n_400)
);

BUFx5_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_312),
.A2(n_237),
.B1(n_283),
.B2(n_296),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_327),
.B(n_142),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_359),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_353),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_381),
.B(n_149),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_349),
.B(n_151),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_321),
.B(n_22),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_317),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_315),
.A2(n_202),
.B1(n_154),
.B2(n_155),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_357),
.B(n_153),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_355),
.B(n_159),
.Y(n_414)
);

OR2x6_ASAP7_75t_L g415 ( 
.A(n_371),
.B(n_223),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_368),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_356),
.B(n_160),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_351),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_302),
.B(n_176),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_190),
.Y(n_421)
);

A2O1A1Ixp33_ASAP7_75t_L g422 ( 
.A1(n_320),
.A2(n_247),
.B(n_289),
.C(n_197),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_309),
.B(n_194),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_L g424 ( 
.A(n_369),
.B(n_247),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_383),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_352),
.B(n_325),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_313),
.B(n_208),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_365),
.B(n_209),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_336),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_333),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_326),
.B(n_247),
.Y(n_431)
);

NOR3xp33_ASAP7_75t_L g432 ( 
.A(n_361),
.B(n_338),
.C(n_326),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_331),
.B(n_289),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_338),
.A2(n_310),
.B1(n_346),
.B2(n_339),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_339),
.B(n_363),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_340),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_346),
.B(n_246),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_303),
.B(n_282),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_332),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_332),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_360),
.A2(n_322),
.B1(n_306),
.B2(n_328),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_308),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_333),
.Y(n_444)
);

NAND3xp33_ASAP7_75t_L g445 ( 
.A(n_310),
.B(n_318),
.C(n_334),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_308),
.Y(n_446)
);

O2A1O1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_310),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_311),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_314),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_323),
.B(n_260),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_324),
.B(n_264),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_404),
.B(n_324),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_429),
.A2(n_379),
.B1(n_328),
.B2(n_334),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_404),
.B(n_330),
.Y(n_454)
);

CKINVDCx8_ASAP7_75t_R g455 ( 
.A(n_430),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_388),
.B(n_379),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_416),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_393),
.B(n_350),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_437),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_434),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_442),
.A2(n_402),
.B(n_396),
.Y(n_461)
);

INVx11_ASAP7_75t_L g462 ( 
.A(n_444),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_393),
.B(n_26),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_402),
.B(n_264),
.C(n_270),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_440),
.B(n_26),
.Y(n_465)
);

INVxp33_ASAP7_75t_SL g466 ( 
.A(n_438),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_389),
.B(n_27),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_385),
.B(n_27),
.Y(n_468)
);

BUFx4f_ASAP7_75t_L g469 ( 
.A(n_415),
.Y(n_469)
);

INVx11_ASAP7_75t_L g470 ( 
.A(n_424),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_410),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_413),
.B(n_30),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_385),
.B(n_30),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_264),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_415),
.A2(n_445),
.B1(n_395),
.B2(n_411),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_400),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_392),
.A2(n_288),
.B1(n_300),
.B2(n_354),
.Y(n_479)
);

O2A1O1Ixp33_ASAP7_75t_L g480 ( 
.A1(n_432),
.A2(n_377),
.B(n_372),
.C(n_370),
.Y(n_480)
);

INVx5_ASAP7_75t_L g481 ( 
.A(n_391),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_449),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_412),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_392),
.B(n_300),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_394),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_398),
.Y(n_488)
);

A2O1A1Ixp33_ASAP7_75t_L g489 ( 
.A1(n_435),
.A2(n_362),
.B(n_347),
.C(n_367),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_435),
.A2(n_443),
.B(n_446),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_409),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_449),
.Y(n_492)
);

OAI321xp33_ASAP7_75t_L g493 ( 
.A1(n_447),
.A2(n_366),
.A3(n_364),
.B1(n_378),
.B2(n_373),
.C(n_348),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_418),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_433),
.A2(n_391),
.B(n_427),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_423),
.B(n_46),
.Y(n_496)
);

AO21x1_ASAP7_75t_L g497 ( 
.A1(n_450),
.A2(n_451),
.B(n_399),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_405),
.Y(n_498)
);

O2A1O1Ixp33_ASAP7_75t_SL g499 ( 
.A1(n_422),
.A2(n_48),
.B(n_50),
.C(n_51),
.Y(n_499)
);

A2O1A1Ixp33_ASAP7_75t_L g500 ( 
.A1(n_408),
.A2(n_390),
.B(n_420),
.C(n_419),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_431),
.A2(n_417),
.B1(n_414),
.B2(n_406),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_448),
.A2(n_348),
.B1(n_329),
.B2(n_316),
.Y(n_502)
);

AO21x1_ASAP7_75t_L g503 ( 
.A1(n_439),
.A2(n_53),
.B(n_55),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_421),
.A2(n_60),
.B(n_65),
.Y(n_504)
);

O2A1O1Ixp33_ASAP7_75t_SL g505 ( 
.A1(n_403),
.A2(n_72),
.B(n_75),
.C(n_76),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_456),
.B(n_407),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_452),
.B(n_401),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_469),
.Y(n_508)
);

BUFx12f_ASAP7_75t_L g509 ( 
.A(n_471),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_454),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_485),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_462),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_488),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_469),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_514)
);

AO31x2_ASAP7_75t_L g515 ( 
.A1(n_489),
.A2(n_101),
.A3(n_102),
.B(n_107),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_460),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_495),
.A2(n_113),
.B(n_116),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_486),
.B(n_487),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_467),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_478),
.B(n_457),
.Y(n_520)
);

O2A1O1Ixp5_ASAP7_75t_L g521 ( 
.A1(n_501),
.A2(n_464),
.B(n_496),
.C(n_461),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_453),
.A2(n_490),
.B1(n_463),
.B2(n_494),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_475),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_485),
.Y(n_524)
);

AO31x2_ASAP7_75t_L g525 ( 
.A1(n_476),
.A2(n_484),
.A3(n_479),
.B(n_504),
.Y(n_525)
);

OAI21x1_ASAP7_75t_SL g526 ( 
.A1(n_490),
.A2(n_473),
.B(n_468),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_485),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_483),
.B(n_465),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_455),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_474),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_481),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_477),
.B(n_482),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_492),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_499),
.A2(n_481),
.B(n_493),
.Y(n_534)
);

AO32x2_ASAP7_75t_L g535 ( 
.A1(n_505),
.A2(n_470),
.A3(n_502),
.B1(n_476),
.B2(n_501),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_458),
.A2(n_442),
.B(n_387),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_452),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_456),
.B(n_404),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_491),
.B(n_425),
.Y(n_539)
);

OA21x2_ASAP7_75t_L g540 ( 
.A1(n_464),
.A2(n_442),
.B(n_461),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_452),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_452),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_458),
.A2(n_442),
.B(n_387),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_455),
.Y(n_544)
);

NAND2x1p5_ASAP7_75t_L g545 ( 
.A(n_469),
.B(n_416),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_469),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_452),
.Y(n_547)
);

AO31x2_ASAP7_75t_L g548 ( 
.A1(n_497),
.A2(n_503),
.A3(n_458),
.B(n_489),
.Y(n_548)
);

AO31x2_ASAP7_75t_L g549 ( 
.A1(n_497),
.A2(n_503),
.A3(n_458),
.B(n_489),
.Y(n_549)
);

AO31x2_ASAP7_75t_L g550 ( 
.A1(n_497),
.A2(n_503),
.A3(n_458),
.B(n_489),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_456),
.B(n_404),
.Y(n_551)
);

OAI21x1_ASAP7_75t_SL g552 ( 
.A1(n_490),
.A2(n_461),
.B(n_459),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_458),
.A2(n_442),
.B(n_387),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_469),
.A2(n_452),
.B1(n_454),
.B2(n_466),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_456),
.B(n_404),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_458),
.A2(n_442),
.B(n_387),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_456),
.B(n_404),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_462),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_452),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_469),
.B(n_416),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_456),
.B(n_404),
.Y(n_561)
);

NOR2x1_ASAP7_75t_SL g562 ( 
.A(n_452),
.B(n_415),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_469),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_458),
.A2(n_437),
.B(n_436),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_491),
.B(n_425),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_456),
.B(n_404),
.Y(n_566)
);

A2O1A1Ixp33_ASAP7_75t_L g567 ( 
.A1(n_480),
.A2(n_500),
.B(n_472),
.C(n_461),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_456),
.B(n_404),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_458),
.A2(n_442),
.B(n_387),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_458),
.A2(n_442),
.B(n_387),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_456),
.B(n_404),
.Y(n_571)
);

AO31x2_ASAP7_75t_L g572 ( 
.A1(n_497),
.A2(n_503),
.A3(n_458),
.B(n_489),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_510),
.A2(n_559),
.B1(n_547),
.B2(n_537),
.Y(n_573)
);

OAI21x1_ASAP7_75t_SL g574 ( 
.A1(n_562),
.A2(n_526),
.B(n_552),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_513),
.Y(n_575)
);

CKINVDCx6p67_ASAP7_75t_R g576 ( 
.A(n_529),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_518),
.Y(n_577)
);

INVx8_ASAP7_75t_L g578 ( 
.A(n_512),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_541),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_567),
.A2(n_521),
.B(n_536),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_542),
.A2(n_554),
.B1(n_522),
.B2(n_516),
.Y(n_581)
);

NOR2xp67_ASAP7_75t_L g582 ( 
.A(n_558),
.B(n_509),
.Y(n_582)
);

OA21x2_ASAP7_75t_L g583 ( 
.A1(n_543),
.A2(n_553),
.B(n_556),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_508),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_555),
.B(n_568),
.Y(n_585)
);

INVx3_ASAP7_75t_SL g586 ( 
.A(n_544),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_519),
.B(n_538),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_551),
.B(n_557),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_520),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_546),
.Y(n_590)
);

OA21x2_ASAP7_75t_L g591 ( 
.A1(n_569),
.A2(n_570),
.B(n_534),
.Y(n_591)
);

BUFx8_ASAP7_75t_L g592 ( 
.A(n_539),
.Y(n_592)
);

OAI22xp33_ASAP7_75t_L g593 ( 
.A1(n_561),
.A2(n_566),
.B1(n_571),
.B2(n_528),
.Y(n_593)
);

INVx8_ASAP7_75t_L g594 ( 
.A(n_565),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_520),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_506),
.B(n_564),
.Y(n_596)
);

NAND2x1p5_ASAP7_75t_L g597 ( 
.A(n_563),
.B(n_531),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_545),
.B(n_560),
.Y(n_598)
);

A2O1A1Ixp33_ASAP7_75t_L g599 ( 
.A1(n_507),
.A2(n_523),
.B(n_517),
.C(n_532),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_530),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_533),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_511),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_515),
.Y(n_603)
);

AOI222xp33_ASAP7_75t_L g604 ( 
.A1(n_514),
.A2(n_527),
.B1(n_511),
.B2(n_524),
.C1(n_535),
.C2(n_540),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_548),
.A2(n_572),
.B(n_549),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g606 ( 
.A1(n_550),
.A2(n_549),
.B(n_525),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_537),
.B(n_541),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_508),
.B(n_546),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_555),
.B(n_568),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_537),
.B(n_541),
.Y(n_610)
);

OAI21x1_ASAP7_75t_SL g611 ( 
.A1(n_562),
.A2(n_526),
.B(n_552),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_555),
.B(n_568),
.Y(n_612)
);

INVx8_ASAP7_75t_L g613 ( 
.A(n_512),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_510),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_512),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_537),
.B(n_541),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_555),
.B(n_568),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_510),
.A2(n_559),
.B1(n_537),
.B2(n_542),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_555),
.B(n_568),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_510),
.A2(n_559),
.B1(n_537),
.B2(n_542),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_510),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_513),
.Y(n_622)
);

BUFx12f_ASAP7_75t_L g623 ( 
.A(n_512),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_537),
.B(n_541),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_555),
.A2(n_432),
.B1(n_460),
.B2(n_568),
.Y(n_625)
);

NAND2x1p5_ASAP7_75t_L g626 ( 
.A(n_508),
.B(n_546),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_531),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_596),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_577),
.B(n_585),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_575),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_L g631 ( 
.A1(n_573),
.A2(n_618),
.B1(n_620),
.B2(n_621),
.Y(n_631)
);

BUFx4f_ASAP7_75t_L g632 ( 
.A(n_626),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_622),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_574),
.B(n_611),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_R g635 ( 
.A(n_578),
.B(n_613),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_614),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_621),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_573),
.B(n_618),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_579),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_607),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_607),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_588),
.B(n_609),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_612),
.B(n_617),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_619),
.B(n_624),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_593),
.A2(n_581),
.B(n_599),
.Y(n_645)
);

INVx3_ASAP7_75t_SL g646 ( 
.A(n_578),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_625),
.A2(n_624),
.B1(n_610),
.B2(n_616),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_583),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_627),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_587),
.A2(n_595),
.B1(n_589),
.B2(n_592),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_603),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_580),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_591),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_606),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_623),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_606),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_594),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_601),
.B(n_605),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_608),
.B(n_597),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_628),
.B(n_605),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_644),
.B(n_604),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_638),
.A2(n_631),
.B1(n_647),
.B2(n_645),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_651),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_640),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_637),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_629),
.B(n_592),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_658),
.B(n_604),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_636),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_658),
.B(n_602),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_654),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_641),
.Y(n_671)
);

NOR2x1_ASAP7_75t_L g672 ( 
.A(n_659),
.B(n_584),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_638),
.A2(n_608),
.B1(n_597),
.B2(n_590),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_652),
.B(n_600),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_656),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_634),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_630),
.B(n_584),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_633),
.B(n_598),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_634),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_634),
.B(n_582),
.Y(n_680)
);

NOR2xp67_ASAP7_75t_L g681 ( 
.A(n_673),
.B(n_649),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_663),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_664),
.B(n_633),
.Y(n_683)
);

NOR2xp67_ASAP7_75t_L g684 ( 
.A(n_673),
.B(n_649),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_671),
.B(n_639),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_661),
.B(n_648),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_674),
.B(n_639),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_668),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_661),
.A2(n_643),
.B1(n_642),
.B2(n_650),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_679),
.B(n_676),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_667),
.B(n_669),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_667),
.B(n_648),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_660),
.B(n_653),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_692),
.B(n_660),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_691),
.B(n_662),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_682),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_688),
.B(n_666),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_691),
.B(n_660),
.Y(n_698)
);

BUFx2_ASAP7_75t_SL g699 ( 
.A(n_681),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_693),
.B(n_670),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_685),
.Y(n_701)
);

AND2x4_ASAP7_75t_SL g702 ( 
.A(n_690),
.B(n_680),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_686),
.B(n_675),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_702),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_701),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_698),
.B(n_686),
.Y(n_706)
);

NOR2x1_ASAP7_75t_L g707 ( 
.A(n_699),
.B(n_672),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_702),
.B(n_700),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_698),
.B(n_687),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_696),
.Y(n_710)
);

NOR2x1_ASAP7_75t_L g711 ( 
.A(n_699),
.B(n_672),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_696),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_707),
.A2(n_681),
.B(n_684),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_705),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_706),
.B(n_695),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_708),
.B(n_704),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_706),
.B(n_694),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_710),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_708),
.B(n_694),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_704),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_712),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_718),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_721),
.B(n_703),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_715),
.B(n_709),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_716),
.B(n_708),
.Y(n_725)
);

OAI221xp5_ASAP7_75t_L g726 ( 
.A1(n_725),
.A2(n_720),
.B1(n_713),
.B2(n_714),
.C(n_689),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_SL g727 ( 
.A(n_723),
.B(n_635),
.C(n_719),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_SL g728 ( 
.A(n_724),
.B(n_646),
.Y(n_728)
);

AND4x1_ASAP7_75t_L g729 ( 
.A(n_728),
.B(n_646),
.C(n_697),
.D(n_711),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_726),
.Y(n_730)
);

NOR3x1_ASAP7_75t_L g731 ( 
.A(n_730),
.B(n_727),
.C(n_723),
.Y(n_731)
);

NOR2x1_ASAP7_75t_L g732 ( 
.A(n_729),
.B(n_646),
.Y(n_732)
);

OAI21xp33_ASAP7_75t_L g733 ( 
.A1(n_732),
.A2(n_716),
.B(n_722),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_731),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_734),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_733),
.B(n_655),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_736),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_736),
.Y(n_738)
);

OAI21xp5_ASAP7_75t_SL g739 ( 
.A1(n_735),
.A2(n_680),
.B(n_626),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_SL g740 ( 
.A1(n_737),
.A2(n_680),
.B(n_576),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_738),
.B(n_586),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_739),
.B(n_717),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_737),
.Y(n_743)
);

NOR2x1p5_ASAP7_75t_L g744 ( 
.A(n_737),
.B(n_615),
.Y(n_744)
);

AO22x2_ASAP7_75t_L g745 ( 
.A1(n_743),
.A2(n_615),
.B1(n_613),
.B2(n_578),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_741),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_744),
.Y(n_747)
);

CKINVDCx16_ASAP7_75t_R g748 ( 
.A(n_742),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_740),
.A2(n_632),
.B(n_716),
.Y(n_749)
);

OAI22x1_ASAP7_75t_L g750 ( 
.A1(n_744),
.A2(n_613),
.B1(n_643),
.B2(n_665),
.Y(n_750)
);

AO22x2_ASAP7_75t_L g751 ( 
.A1(n_743),
.A2(n_657),
.B1(n_719),
.B2(n_717),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_745),
.B(n_702),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_748),
.A2(n_632),
.B1(n_659),
.B2(n_683),
.Y(n_753)
);

AOI21xp33_ASAP7_75t_L g754 ( 
.A1(n_746),
.A2(n_747),
.B(n_750),
.Y(n_754)
);

INVx3_ASAP7_75t_SL g755 ( 
.A(n_751),
.Y(n_755)
);

OR2x6_ASAP7_75t_L g756 ( 
.A(n_752),
.B(n_749),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_755),
.A2(n_674),
.B1(n_679),
.B2(n_677),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_754),
.B(n_678),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_756),
.A2(n_753),
.B(n_632),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_758),
.A2(n_632),
.B(n_659),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_759),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_761),
.A2(n_760),
.B1(n_757),
.B2(n_659),
.Y(n_762)
);


endmodule