module real_jpeg_16523_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_249;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_243;
wire n_105;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_0),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_2),
.B(n_46),
.Y(n_45)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_2),
.B(n_67),
.Y(n_66)
);

NAND2x1_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_2),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_2),
.B(n_135),
.Y(n_134)
);

NAND2x1_ASAP7_75t_L g183 ( 
.A(n_2),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_3),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_3),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_3),
.B(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_4),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_4),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_4),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_4),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_4),
.B(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_7),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_7),
.Y(n_175)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_7),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_36),
.Y(n_35)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_8),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_8),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_8),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g172 ( 
.A(n_8),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_8),
.B(n_184),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

BUFx8_ASAP7_75t_L g184 ( 
.A(n_11),
.Y(n_184)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_11),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_232),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_231),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_197),
.Y(n_16)
);

OAI21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_160),
.B(n_196),
.Y(n_17)
);

AOI21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_112),
.B(n_159),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_20),
.B(n_73),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_43),
.C(n_59),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_21),
.B(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_22),
.Y(n_150)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_23),
.A2(n_35),
.B(n_42),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_24),
.A2(n_25),
.B1(n_108),
.B2(n_111),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_38),
.B(n_40),
.Y(n_37)
);

NAND2x1p5_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_38),
.Y(n_40)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_28),
.Y(n_139)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_28),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_29),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_29),
.Y(n_141)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_R g133 ( 
.A1(n_35),
.A2(n_134),
.B(n_136),
.C(n_142),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_35),
.B(n_134),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_35),
.A2(n_41),
.B1(n_134),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_38),
.A2(n_123),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_38),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_38),
.B(n_137),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_38),
.A2(n_129),
.B1(n_137),
.B2(n_140),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_40),
.B(n_78),
.C(n_84),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_43),
.A2(n_59),
.B1(n_60),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.C(n_54),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_44),
.A2(n_45),
.B1(n_54),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_44),
.A2(n_45),
.B1(n_172),
.B2(n_176),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_45),
.B(n_209),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_45),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_50),
.B1(n_91),
.B2(n_101),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_49),
.A2(n_50),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_50),
.A2(n_93),
.B(n_95),
.C(n_142),
.Y(n_167)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_53),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_54),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_54),
.A2(n_78),
.B1(n_86),
.B2(n_120),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_55),
.B(n_109),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_55),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_72),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_61),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_66),
.C(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_66),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_66),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_68),
.Y(n_193)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_69),
.A2(n_105),
.B1(n_171),
.B2(n_177),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_72),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_89),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_87),
.B2(n_88),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_76),
.B(n_87),
.C(n_89),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_86),
.B(n_120),
.C(n_204),
.Y(n_255)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_102),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_103),
.C(n_107),
.Y(n_164)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_100),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_92),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_92),
.B(n_149),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_92),
.B(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_93),
.B(n_134),
.C(n_183),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_94),
.Y(n_260)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_105),
.B(n_137),
.C(n_172),
.Y(n_228)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_108),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_108),
.A2(n_111),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_108),
.B(n_220),
.C(n_223),
.Y(n_262)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_122),
.B(n_123),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_131),
.B(n_158),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_117),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_127),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_127),
.B1(n_128),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_146),
.B(n_157),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_143),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_134),
.A2(n_155),
.B1(n_208),
.B2(n_213),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_134),
.B(n_210),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_140),
.B1(n_172),
.B2(n_176),
.Y(n_171)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_153),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_152),
.B(n_156),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_150),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_155),
.B(n_209),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_162),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_178),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_165),
.C(n_178),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_170),
.C(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_195),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_186),
.C(n_195),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_185),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_191),
.B(n_194),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_191),
.Y(n_194)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_194),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_199),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_216),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_200),
.B(n_217),
.C(n_230),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_214),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_206),
.C(n_214),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_230),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_226),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_228),
.C(n_229),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_267),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_266),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_266),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_253),
.Y(n_237)
);

XOR2x2_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_251),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_247),
.B2(n_248),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_265),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_263),
.B2(n_264),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_262),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_259),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);


endmodule