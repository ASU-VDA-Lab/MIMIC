module fake_aes_1655_n_728 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_728);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_728;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_565;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_195;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_16), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_29), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_54), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_15), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_47), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_43), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_53), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_75), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_31), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_52), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_56), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_33), .Y(n_92) );
BUFx2_ASAP7_75t_L g93 ( .A(n_13), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_7), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_45), .Y(n_95) );
BUFx3_ASAP7_75t_L g96 ( .A(n_68), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_2), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_38), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_48), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_71), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_27), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_35), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_25), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_65), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_69), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_62), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_59), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_8), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_26), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_58), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_63), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_7), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_14), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_14), .Y(n_115) );
INVxp33_ASAP7_75t_L g116 ( .A(n_21), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_72), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_15), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_19), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_26), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_11), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_13), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_30), .Y(n_123) );
INVxp33_ASAP7_75t_L g124 ( .A(n_9), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_61), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_42), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_3), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_23), .Y(n_128) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_74), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_6), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_108), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_82), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_90), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_93), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_108), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_82), .Y(n_136) );
OAI21x1_ASAP7_75t_L g137 ( .A1(n_90), .A2(n_34), .B(n_79), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_128), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_98), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_108), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_93), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_93), .B(n_0), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_83), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_98), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_85), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g148 ( .A(n_128), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_85), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_81), .Y(n_151) );
INVx6_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_116), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_86), .Y(n_154) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_86), .A2(n_36), .B(n_78), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_89), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_96), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
BUFx2_ASAP7_75t_L g159 ( .A(n_113), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_107), .Y(n_160) );
INVxp67_ASAP7_75t_L g161 ( .A(n_94), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g162 ( .A1(n_84), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_89), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_127), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_102), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_88), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_116), .B(n_4), .Y(n_167) );
NAND2xp33_ASAP7_75t_L g168 ( .A(n_91), .B(n_80), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_107), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_92), .Y(n_170) );
INVxp33_ASAP7_75t_L g171 ( .A(n_124), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_92), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_124), .B(n_5), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_107), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_87), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_153), .B(n_91), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_153), .B(n_95), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
OR2x2_ASAP7_75t_L g182 ( .A(n_171), .B(n_84), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_142), .A2(n_112), .B1(n_101), .B2(n_120), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_134), .B(n_95), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_133), .Y(n_186) );
OAI221xp5_ASAP7_75t_L g187 ( .A1(n_134), .A2(n_112), .B1(n_101), .B2(n_120), .C(n_130), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_142), .B(n_144), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_161), .B(n_130), .Y(n_189) );
BUFx2_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_159), .B(n_111), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_156), .B(n_111), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_175), .B(n_100), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_161), .B(n_100), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_150), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_142), .Y(n_196) );
AND2x6_ASAP7_75t_L g197 ( .A(n_142), .B(n_99), .Y(n_197) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_133), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_150), .Y(n_200) );
AO22x2_ASAP7_75t_L g201 ( .A1(n_167), .A2(n_129), .B1(n_126), .B2(n_99), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_143), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_144), .A2(n_104), .B(n_125), .C(n_126), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
INVxp67_ASAP7_75t_L g205 ( .A(n_167), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_146), .B(n_105), .Y(n_206) );
INVx5_ASAP7_75t_L g207 ( .A(n_152), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_146), .B(n_114), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_150), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_147), .B(n_105), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_147), .B(n_123), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_149), .B(n_115), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_149), .B(n_123), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_143), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_140), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_137), .Y(n_216) );
AND2x6_ASAP7_75t_L g217 ( .A(n_160), .B(n_106), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_131), .Y(n_218) );
NAND2x1p5_ASAP7_75t_L g219 ( .A(n_154), .B(n_106), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_131), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_140), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_173), .A2(n_115), .B1(n_97), .B2(n_122), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_157), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_154), .B(n_114), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_163), .B(n_117), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_135), .Y(n_227) );
AO22x2_ASAP7_75t_L g228 ( .A1(n_158), .A2(n_129), .B1(n_117), .B2(n_110), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_157), .Y(n_229) );
OR2x2_ASAP7_75t_L g230 ( .A(n_173), .B(n_94), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_135), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_136), .B(n_97), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_157), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_158), .B(n_118), .Y(n_234) );
NAND2xp33_ASAP7_75t_R g235 ( .A(n_165), .B(n_103), .Y(n_235) );
BUFx6f_ASAP7_75t_SL g236 ( .A(n_166), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_166), .B(n_110), .Y(n_237) );
INVx4_ASAP7_75t_L g238 ( .A(n_160), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_170), .B(n_118), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_157), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_170), .B(n_125), .Y(n_241) );
NAND2xp33_ASAP7_75t_L g242 ( .A(n_172), .B(n_125), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_215), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_183), .A2(n_141), .B1(n_145), .B2(n_139), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_219), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_216), .Y(n_246) );
INVxp67_ASAP7_75t_SL g247 ( .A(n_219), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_190), .Y(n_248) );
AND2x6_ASAP7_75t_L g249 ( .A(n_188), .B(n_160), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_178), .B(n_172), .Y(n_250) );
CKINVDCx8_ASAP7_75t_R g251 ( .A(n_190), .Y(n_251) );
NOR2xp33_ASAP7_75t_R g252 ( .A(n_236), .B(n_164), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_215), .Y(n_253) );
NOR3xp33_ASAP7_75t_SL g254 ( .A(n_235), .B(n_148), .C(n_162), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_228), .A2(n_140), .B1(n_160), .B2(n_109), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_215), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_219), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_188), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_216), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_189), .B(n_140), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_201), .B(n_162), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_239), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_189), .B(n_141), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_236), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g265 ( .A(n_198), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_201), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_230), .B(n_168), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_188), .B(n_152), .Y(n_268) );
INVx6_ASAP7_75t_L g269 ( .A(n_196), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_239), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_188), .B(n_152), .Y(n_271) );
OAI21xp33_ASAP7_75t_SL g272 ( .A1(n_196), .A2(n_137), .B(n_122), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_230), .B(n_152), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_205), .B(n_103), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_182), .B(n_151), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_239), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_181), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_201), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_236), .Y(n_279) );
OR2x4_ASAP7_75t_L g280 ( .A(n_182), .B(n_148), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_228), .A2(n_109), .B1(n_119), .B2(n_121), .Y(n_281) );
NOR3xp33_ASAP7_75t_SL g282 ( .A(n_187), .B(n_119), .C(n_121), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_197), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_239), .Y(n_284) );
NOR3xp33_ASAP7_75t_SL g285 ( .A(n_226), .B(n_138), .C(n_6), .Y(n_285) );
NAND2xp33_ASAP7_75t_SL g286 ( .A(n_196), .B(n_104), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_196), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_228), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_208), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_215), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_208), .Y(n_292) );
INVxp67_ASAP7_75t_SL g293 ( .A(n_221), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_212), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_212), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_201), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_225), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_225), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_234), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_183), .A2(n_104), .B1(n_169), .B2(n_157), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_234), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_197), .B(n_137), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_180), .A2(n_174), .B1(n_169), .B2(n_155), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_185), .B(n_5), .Y(n_304) );
NOR2xp33_ASAP7_75t_R g305 ( .A(n_197), .B(n_8), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_194), .B(n_174), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_191), .B(n_174), .Y(n_307) );
INVx2_ASAP7_75t_SL g308 ( .A(n_197), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_197), .B(n_174), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_197), .Y(n_310) );
INVx5_ASAP7_75t_L g311 ( .A(n_217), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_176), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_181), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_197), .B(n_174), .Y(n_314) );
INVxp67_ASAP7_75t_L g315 ( .A(n_247), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_262), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_272), .A2(n_203), .B(n_227), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_290), .B(n_193), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_248), .Y(n_319) );
CKINVDCx11_ASAP7_75t_R g320 ( .A(n_251), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_292), .B(n_232), .Y(n_321) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_245), .B(n_238), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_265), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_251), .B(n_232), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_288), .Y(n_325) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_303), .A2(n_213), .B(n_206), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_267), .B(n_228), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_270), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_294), .B(n_222), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_275), .B(n_222), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_281), .A2(n_210), .B1(n_211), .B2(n_241), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_263), .B(n_192), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_263), .A2(n_242), .B1(n_217), .B2(n_237), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_263), .B(n_214), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_284), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_297), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_280), .B(n_238), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_267), .B(n_217), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_250), .B(n_217), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_269), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_281), .A2(n_204), .B1(n_202), .B2(n_199), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_298), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_299), .B(n_221), .Y(n_345) );
INVxp67_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_311), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_302), .A2(n_216), .B(n_238), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_248), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_311), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_255), .A2(n_204), .B1(n_202), .B2(n_199), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_257), .A2(n_217), .B1(n_220), .B2(n_218), .Y(n_353) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_266), .B(n_238), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_278), .A2(n_296), .B1(n_258), .B2(n_289), .Y(n_355) );
BUFx12f_ASAP7_75t_L g356 ( .A(n_264), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_258), .B(n_217), .Y(n_357) );
CKINVDCx6p67_ASAP7_75t_R g358 ( .A(n_261), .Y(n_358) );
OR2x6_ASAP7_75t_L g359 ( .A(n_261), .B(n_216), .Y(n_359) );
BUFx12f_ASAP7_75t_L g360 ( .A(n_264), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_260), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_311), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_288), .Y(n_363) );
OAI21xp33_ASAP7_75t_L g364 ( .A1(n_255), .A2(n_218), .B(n_231), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_261), .A2(n_217), .B1(n_220), .B2(n_231), .Y(n_365) );
INVxp67_ASAP7_75t_L g366 ( .A(n_274), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_302), .B(n_227), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_252), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_302), .A2(n_221), .B(n_176), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_286), .A2(n_221), .B(n_155), .Y(n_370) );
INVx5_ASAP7_75t_L g371 ( .A(n_347), .Y(n_371) );
INVx4_ASAP7_75t_L g372 ( .A(n_347), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_316), .Y(n_373) );
OAI22xp33_ASAP7_75t_SL g374 ( .A1(n_359), .A2(n_261), .B1(n_279), .B2(n_244), .Y(n_374) );
NAND3x1_ASAP7_75t_L g375 ( .A(n_358), .B(n_254), .C(n_300), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_347), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_322), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_327), .A2(n_312), .B1(n_273), .B2(n_283), .Y(n_378) );
AOI22xp33_ASAP7_75t_SL g379 ( .A1(n_324), .A2(n_252), .B1(n_305), .B2(n_279), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_320), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_315), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_322), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g383 ( .A1(n_331), .A2(n_280), .B1(n_283), .B2(n_310), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_328), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_366), .B(n_307), .Y(n_385) );
BUFx10_ASAP7_75t_L g386 ( .A(n_354), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_330), .B(n_249), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_335), .B(n_286), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_330), .B(n_282), .Y(n_389) );
AOI22xp33_ASAP7_75t_SL g390 ( .A1(n_319), .A2(n_305), .B1(n_249), .B2(n_308), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_325), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_333), .A2(n_249), .B1(n_288), .B2(n_269), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_346), .B(n_269), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_323), .B(n_268), .Y(n_394) );
INVx3_ASAP7_75t_SL g395 ( .A(n_349), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_363), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_321), .B(n_271), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_337), .A2(n_285), .B1(n_293), .B2(n_243), .C(n_253), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_361), .B(n_186), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_329), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_368), .A2(n_249), .B1(n_308), .B2(n_311), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_367), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_315), .B(n_186), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_321), .B(n_249), .Y(n_404) );
OR2x6_ASAP7_75t_L g405 ( .A(n_359), .B(n_246), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_402), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_402), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_380), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_402), .Y(n_409) );
AOI222xp33_ASAP7_75t_L g410 ( .A1(n_389), .A2(n_338), .B1(n_344), .B2(n_352), .C1(n_318), .C2(n_327), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_381), .A2(n_359), .B1(n_355), .B2(n_332), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_381), .B(n_343), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_389), .A2(n_332), .B1(n_318), .B2(n_336), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_378), .A2(n_388), .B1(n_387), .B2(n_385), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_399), .B(n_369), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_371), .Y(n_416) );
OAI22xp33_ASAP7_75t_SL g417 ( .A1(n_378), .A2(n_334), .B1(n_369), .B2(n_367), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_374), .A2(n_345), .B1(n_364), .B2(n_317), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_390), .A2(n_365), .B1(n_343), .B2(n_351), .Y(n_419) );
AOI221x1_ASAP7_75t_L g420 ( .A1(n_374), .A2(n_370), .B1(n_317), .B2(n_348), .C(n_351), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_391), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_395), .Y(n_422) );
OA21x2_ASAP7_75t_L g423 ( .A1(n_373), .A2(n_370), .B(n_348), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_387), .A2(n_345), .B1(n_339), .B2(n_326), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_398), .B(n_169), .C(n_174), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_391), .Y(n_426) );
AOI322xp5_ASAP7_75t_L g427 ( .A1(n_383), .A2(n_356), .A3(n_360), .B1(n_214), .B2(n_306), .C1(n_16), .C2(n_17), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_377), .Y(n_428) );
OAI21xp33_ASAP7_75t_L g429 ( .A1(n_403), .A2(n_340), .B(n_341), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_388), .A2(n_326), .B1(n_214), .B2(n_340), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_377), .B(n_362), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g432 ( .A1(n_373), .A2(n_341), .B1(n_214), .B2(n_342), .C(n_357), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_385), .Y(n_433) );
OAI21x1_ASAP7_75t_L g434 ( .A1(n_375), .A2(n_155), .B(n_309), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_403), .A2(n_397), .B1(n_384), .B2(n_400), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_410), .A2(n_386), .B1(n_384), .B2(n_400), .Y(n_436) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_427), .B(n_377), .C(n_382), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_413), .A2(n_379), .B1(n_397), .B2(n_404), .C(n_394), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_421), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_416), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_416), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_406), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_410), .A2(n_386), .B1(n_395), .B2(n_399), .Y(n_443) );
NAND2xp33_ASAP7_75t_R g444 ( .A(n_422), .B(n_155), .Y(n_444) );
OAI22xp5_ASAP7_75t_SL g445 ( .A1(n_413), .A2(n_395), .B1(n_382), .B2(n_405), .Y(n_445) );
NOR2x1_ASAP7_75t_L g446 ( .A(n_416), .B(n_405), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_412), .B(n_382), .Y(n_447) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_407), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_427), .B(n_169), .C(n_393), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_421), .Y(n_450) );
OAI22xp33_ASAP7_75t_L g451 ( .A1(n_412), .A2(n_405), .B1(n_386), .B2(n_372), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_411), .A2(n_386), .B1(n_392), .B2(n_394), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_415), .B(n_391), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_407), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_412), .B(n_406), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_425), .A2(n_375), .B(n_353), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_435), .A2(n_405), .B1(n_396), .B2(n_372), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_409), .B(n_396), .Y(n_459) );
NOR2xp33_ASAP7_75t_R g460 ( .A(n_408), .B(n_371), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_409), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_409), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_411), .A2(n_405), .B1(n_396), .B2(n_342), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_419), .A2(n_372), .B1(n_401), .B2(n_376), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_425), .A2(n_376), .B(n_357), .C(n_371), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_421), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_419), .A2(n_372), .B1(n_371), .B2(n_376), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_428), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_426), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_426), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_431), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_415), .B(n_376), .Y(n_472) );
BUFx3_ASAP7_75t_L g473 ( .A(n_440), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_454), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_455), .B(n_414), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_455), .B(n_433), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_442), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_439), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_472), .B(n_415), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_472), .B(n_428), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_442), .Y(n_481) );
AO22x1_ASAP7_75t_L g482 ( .A1(n_458), .A2(n_433), .B1(n_428), .B2(n_431), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_454), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_449), .A2(n_414), .B1(n_417), .B2(n_418), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_447), .B(n_428), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_439), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_472), .B(n_428), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_439), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_436), .B(n_435), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_462), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_462), .Y(n_491) );
OAI33xp33_ASAP7_75t_L g492 ( .A1(n_449), .A2(n_417), .A3(n_429), .B1(n_11), .B2(n_12), .B3(n_17), .Y(n_492) );
NAND2xp67_ASAP7_75t_L g493 ( .A(n_459), .B(n_426), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_450), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_448), .Y(n_495) );
OAI31xp33_ASAP7_75t_L g496 ( .A1(n_438), .A2(n_436), .A3(n_443), .B(n_451), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_438), .B(n_9), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_448), .B(n_424), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_453), .B(n_418), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_450), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_459), .B(n_424), .Y(n_501) );
NAND3xp33_ASAP7_75t_SL g502 ( .A(n_460), .B(n_432), .C(n_430), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_459), .B(n_430), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_466), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_466), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_445), .B(n_10), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_461), .B(n_423), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_452), .A2(n_429), .B1(n_432), .B2(n_423), .C(n_314), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_453), .B(n_420), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_450), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_469), .Y(n_511) );
AND2x4_ASAP7_75t_SL g512 ( .A(n_441), .B(n_431), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_447), .B(n_420), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g514 ( .A1(n_445), .A2(n_431), .B1(n_434), .B2(n_371), .C1(n_19), .C2(n_20), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_440), .Y(n_515) );
AOI22x1_ASAP7_75t_L g516 ( .A1(n_441), .A2(n_431), .B1(n_169), .B2(n_362), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_461), .B(n_423), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_469), .B(n_423), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_469), .B(n_423), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_470), .B(n_434), .Y(n_520) );
OAI31xp33_ASAP7_75t_SL g521 ( .A1(n_458), .A2(n_434), .A3(n_12), .B(n_18), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_470), .B(n_371), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_456), .B(n_10), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_437), .A2(n_246), .B1(n_259), .B2(n_287), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_518), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_479), .B(n_470), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_479), .B(n_456), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_474), .B(n_456), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_518), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_478), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_491), .B(n_456), .Y(n_531) );
NAND5xp2_ASAP7_75t_SL g532 ( .A(n_496), .B(n_464), .C(n_467), .D(n_463), .E(n_457), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_495), .B(n_471), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_476), .B(n_471), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_478), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_503), .B(n_467), .Y(n_536) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_497), .A2(n_437), .B1(n_451), .B2(n_457), .C(n_169), .Y(n_537) );
OAI33xp33_ASAP7_75t_L g538 ( .A1(n_489), .A2(n_18), .A3(n_20), .B1(n_21), .B2(n_22), .B3(n_23), .Y(n_538) );
NOR2xp33_ASAP7_75t_R g539 ( .A(n_473), .B(n_440), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_476), .B(n_441), .Y(n_540) );
OAI33xp33_ASAP7_75t_L g541 ( .A1(n_477), .A2(n_24), .A3(n_25), .B1(n_27), .B2(n_223), .B3(n_184), .Y(n_541) );
NAND4xp25_ASAP7_75t_SL g542 ( .A(n_514), .B(n_446), .C(n_465), .D(n_444), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_493), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_477), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_481), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_481), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_503), .B(n_468), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_478), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_495), .B(n_483), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_501), .B(n_468), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_501), .B(n_468), .Y(n_551) );
NAND2xp33_ASAP7_75t_SL g552 ( .A(n_523), .B(n_441), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_507), .B(n_468), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_504), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_475), .B(n_504), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_507), .B(n_446), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_514), .B(n_184), .C(n_195), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_473), .B(n_66), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_505), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_480), .B(n_24), .Y(n_560) );
NAND2xp33_ASAP7_75t_SL g561 ( .A(n_523), .B(n_259), .Y(n_561) );
NOR2xp33_ASAP7_75t_R g562 ( .A(n_473), .B(n_350), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_521), .B(n_506), .C(n_496), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_480), .B(n_223), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_475), .B(n_184), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_515), .B(n_28), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_499), .B(n_195), .Y(n_567) );
BUFx4f_ASAP7_75t_SL g568 ( .A(n_515), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_487), .B(n_223), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_487), .B(n_32), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_493), .Y(n_571) );
NAND3xp33_ASAP7_75t_SL g572 ( .A(n_484), .B(n_195), .C(n_200), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_499), .B(n_200), .Y(n_573) );
NAND2xp33_ASAP7_75t_R g574 ( .A(n_517), .B(n_37), .Y(n_574) );
NAND2x1_ASAP7_75t_L g575 ( .A(n_510), .B(n_246), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_483), .B(n_200), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_490), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_490), .B(n_209), .Y(n_578) );
BUFx2_ASAP7_75t_L g579 ( .A(n_517), .Y(n_579) );
BUFx3_ASAP7_75t_L g580 ( .A(n_512), .Y(n_580) );
BUFx3_ASAP7_75t_L g581 ( .A(n_512), .Y(n_581) );
NAND2xp33_ASAP7_75t_R g582 ( .A(n_519), .B(n_39), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_486), .Y(n_583) );
AOI211xp5_ASAP7_75t_L g584 ( .A1(n_521), .A2(n_209), .B(n_224), .C(n_229), .Y(n_584) );
AOI31xp33_ASAP7_75t_L g585 ( .A1(n_582), .A2(n_492), .A3(n_502), .B(n_524), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g586 ( .A1(n_563), .A2(n_524), .B(n_522), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_537), .A2(n_522), .B1(n_485), .B2(n_498), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_577), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_574), .A2(n_482), .B1(n_498), .B2(n_513), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_579), .Y(n_590) );
OAI21xp33_ASAP7_75t_L g591 ( .A1(n_542), .A2(n_509), .B(n_513), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_555), .B(n_509), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_568), .A2(n_516), .B1(n_485), .B2(n_519), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_538), .A2(n_482), .B1(n_508), .B2(n_510), .C(n_511), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_550), .B(n_512), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_549), .Y(n_596) );
OAI21xp5_ASAP7_75t_SL g597 ( .A1(n_560), .A2(n_520), .B(n_486), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_580), .A2(n_520), .B1(n_488), .B2(n_511), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_560), .A2(n_552), .B1(n_541), .B2(n_540), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_549), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_552), .A2(n_511), .B(n_500), .C(n_494), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_544), .B(n_500), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g603 ( .A1(n_580), .A2(n_516), .B1(n_500), .B2(n_494), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_545), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_526), .B(n_494), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_571), .A2(n_486), .B1(n_488), .B2(n_209), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_525), .B(n_488), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_525), .B(n_229), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_543), .B(n_40), .Y(n_609) );
AO22x1_ASAP7_75t_L g610 ( .A1(n_581), .A2(n_362), .B1(n_350), .B2(n_287), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_546), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_570), .A2(n_224), .B1(n_229), .B2(n_177), .Y(n_612) );
AOI322xp5_ASAP7_75t_L g613 ( .A1(n_536), .A2(n_224), .A3(n_179), .B1(n_177), .B2(n_233), .C1(n_240), .C2(n_253), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_554), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_559), .Y(n_615) );
AOI222xp33_ASAP7_75t_L g616 ( .A1(n_536), .A2(n_179), .B1(n_233), .B2(n_240), .C1(n_291), .C2(n_243), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_539), .B(n_350), .Y(n_617) );
INVx3_ASAP7_75t_L g618 ( .A(n_581), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_529), .B(n_41), .Y(n_619) );
NOR3xp33_ASAP7_75t_SL g620 ( .A(n_557), .B(n_44), .C(n_46), .Y(n_620) );
AOI32xp33_ASAP7_75t_L g621 ( .A1(n_561), .A2(n_291), .A3(n_256), .B1(n_181), .B2(n_313), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_562), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_550), .B(n_49), .Y(n_623) );
NAND4xp25_ASAP7_75t_SL g624 ( .A(n_584), .B(n_50), .C(n_51), .D(n_55), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_579), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_527), .Y(n_626) );
AO21x1_ASAP7_75t_L g627 ( .A1(n_561), .A2(n_57), .B(n_60), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_534), .Y(n_628) );
OAI21xp5_ASAP7_75t_SL g629 ( .A1(n_558), .A2(n_259), .B(n_246), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_565), .B(n_287), .C(n_259), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_551), .B(n_64), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_570), .A2(n_256), .B1(n_287), .B2(n_277), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_532), .A2(n_313), .B1(n_277), .B2(n_207), .C(n_73), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_529), .B(n_67), .Y(n_634) );
INVxp67_ASAP7_75t_SL g635 ( .A(n_533), .Y(n_635) );
INVx1_ASAP7_75t_SL g636 ( .A(n_528), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_556), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_528), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_596), .B(n_600), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_629), .A2(n_575), .B(n_532), .Y(n_640) );
XNOR2xp5_ASAP7_75t_L g641 ( .A(n_622), .B(n_556), .Y(n_641) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_585), .A2(n_533), .B1(n_531), .B2(n_575), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_590), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_626), .B(n_551), .Y(n_644) );
INVxp67_ASAP7_75t_L g645 ( .A(n_635), .Y(n_645) );
INVx3_ASAP7_75t_L g646 ( .A(n_618), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_607), .Y(n_647) );
AOI21xp33_ASAP7_75t_L g648 ( .A1(n_591), .A2(n_566), .B(n_567), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_604), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_636), .B(n_531), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_637), .B(n_553), .Y(n_651) );
NOR2x1_ASAP7_75t_L g652 ( .A(n_617), .B(n_558), .Y(n_652) );
AO22x1_ASAP7_75t_L g653 ( .A1(n_618), .A2(n_586), .B1(n_598), .B2(n_625), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_611), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_588), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_614), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_638), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_628), .B(n_547), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_615), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_597), .A2(n_558), .B(n_570), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_595), .B(n_553), .Y(n_661) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_593), .B(n_624), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_605), .B(n_547), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_589), .B(n_548), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_598), .B(n_548), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_592), .B(n_564), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_607), .B(n_583), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_627), .B(n_583), .Y(n_668) );
INVx3_ASAP7_75t_L g669 ( .A(n_602), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_608), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_586), .B(n_535), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_599), .B(n_569), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_608), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_594), .B(n_569), .Y(n_674) );
OAI21xp33_ASAP7_75t_L g675 ( .A1(n_633), .A2(n_573), .B(n_564), .Y(n_675) );
XNOR2xp5_ASAP7_75t_L g676 ( .A(n_587), .B(n_572), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_639), .B(n_535), .Y(n_677) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_660), .A2(n_587), .B(n_621), .Y(n_678) );
OAI21xp33_ASAP7_75t_L g679 ( .A1(n_662), .A2(n_601), .B(n_620), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_653), .A2(n_609), .B1(n_603), .B2(n_619), .C(n_623), .Y(n_680) );
AOI321xp33_ASAP7_75t_L g681 ( .A1(n_674), .A2(n_631), .A3(n_619), .B1(n_606), .B2(n_632), .C(n_634), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_671), .B(n_530), .Y(n_682) );
NOR2x1_ASAP7_75t_L g683 ( .A(n_641), .B(n_630), .Y(n_683) );
INVx1_ASAP7_75t_SL g684 ( .A(n_641), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_672), .A2(n_616), .B1(n_612), .B2(n_610), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_671), .B(n_530), .Y(n_686) );
XNOR2xp5_ASAP7_75t_L g687 ( .A(n_676), .B(n_578), .Y(n_687) );
NAND3x2_ASAP7_75t_L g688 ( .A(n_650), .B(n_613), .C(n_70), .Y(n_688) );
AOI32xp33_ASAP7_75t_L g689 ( .A1(n_642), .A2(n_652), .A3(n_646), .B1(n_661), .B2(n_665), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_653), .A2(n_576), .B1(n_207), .B2(n_77), .C(n_76), .Y(n_690) );
BUFx2_ASAP7_75t_L g691 ( .A(n_646), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_676), .A2(n_207), .B(n_640), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_669), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_663), .B(n_207), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_645), .A2(n_207), .B1(n_666), .B2(n_643), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_669), .B(n_657), .Y(n_696) );
INVx2_ASAP7_75t_SL g697 ( .A(n_677), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_678), .A2(n_664), .B1(n_658), .B2(n_665), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_688), .A2(n_648), .B1(n_675), .B2(n_670), .Y(n_699) );
INVxp33_ASAP7_75t_SL g700 ( .A(n_687), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_689), .A2(n_655), .B1(n_659), .B2(n_656), .C(n_649), .Y(n_701) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_683), .B(n_668), .Y(n_702) );
INVx2_ASAP7_75t_SL g703 ( .A(n_691), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_679), .A2(n_669), .B1(n_650), .B2(n_649), .C(n_654), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_696), .Y(n_705) );
NOR2xp33_ASAP7_75t_R g706 ( .A(n_687), .B(n_684), .Y(n_706) );
OAI211xp5_ASAP7_75t_SL g707 ( .A1(n_692), .A2(n_644), .B(n_673), .C(n_639), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_695), .A2(n_647), .B1(n_651), .B2(n_673), .C(n_661), .Y(n_708) );
NOR2xp67_ASAP7_75t_L g709 ( .A(n_693), .B(n_647), .Y(n_709) );
NAND3xp33_ASAP7_75t_SL g710 ( .A(n_690), .B(n_667), .C(n_651), .Y(n_710) );
NAND4xp75_ASAP7_75t_L g711 ( .A(n_680), .B(n_685), .C(n_694), .D(n_686), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_682), .A2(n_689), .B1(n_684), .B2(n_678), .C(n_679), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_694), .A2(n_678), .B1(n_684), .B2(n_683), .Y(n_713) );
NOR3x2_ASAP7_75t_L g714 ( .A(n_681), .B(n_688), .C(n_679), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_712), .A2(n_701), .B1(n_700), .B2(n_713), .C(n_706), .Y(n_715) );
NOR2x1_ASAP7_75t_L g716 ( .A(n_702), .B(n_711), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_698), .B(n_708), .Y(n_717) );
XOR2x2_ASAP7_75t_L g718 ( .A(n_710), .B(n_714), .Y(n_718) );
NAND4xp75_ASAP7_75t_L g719 ( .A(n_703), .B(n_705), .C(n_709), .D(n_697), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_717), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_718), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_715), .A2(n_704), .B1(n_707), .B2(n_699), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_720), .Y(n_723) );
INVxp33_ASAP7_75t_L g724 ( .A(n_721), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_723), .Y(n_725) );
INVx4_ASAP7_75t_L g726 ( .A(n_723), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_726), .A2(n_716), .B1(n_724), .B2(n_722), .Y(n_727) );
O2A1O1Ixp5_ASAP7_75t_L g728 ( .A1(n_727), .A2(n_726), .B(n_725), .C(n_719), .Y(n_728) );
endmodule