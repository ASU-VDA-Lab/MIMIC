module fake_jpeg_25703_n_322 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_38),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_34),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_9),
.B(n_15),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_14),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_64),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_57),
.Y(n_76)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_26),
.B1(n_23),
.B2(n_32),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_25),
.B1(n_18),
.B2(n_30),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_25),
.B1(n_18),
.B2(n_30),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_67),
.B1(n_17),
.B2(n_32),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_17),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_63),
.Y(n_85)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_66),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_24),
.B1(n_34),
.B2(n_31),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_87),
.Y(n_114)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_77),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_22),
.B1(n_33),
.B2(n_29),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_78),
.A2(n_83),
.B1(n_53),
.B2(n_45),
.Y(n_123)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_17),
.A3(n_32),
.B1(n_28),
.B2(n_20),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_29),
.A3(n_20),
.B1(n_28),
.B2(n_22),
.Y(n_109)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_84),
.Y(n_108)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_91),
.B1(n_94),
.B2(n_48),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_22),
.B1(n_33),
.B2(n_29),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_46),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_36),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_22),
.B1(n_33),
.B2(n_20),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_27),
.Y(n_98)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

AO22x2_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_98),
.A2(n_110),
.B1(n_123),
.B2(n_74),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_76),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_20),
.B(n_28),
.Y(n_150)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_113),
.Y(n_153)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_85),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_66),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_117),
.B(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_58),
.B1(n_69),
.B2(n_45),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_119),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_66),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_79),
.C(n_87),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_58),
.B1(n_45),
.B2(n_64),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_55),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_124),
.B(n_70),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_124),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_138),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_139),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_120),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_42),
.C(n_43),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_98),
.C(n_49),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_117),
.A2(n_80),
.B1(n_93),
.B2(n_96),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_130),
.A2(n_133),
.B1(n_146),
.B2(n_154),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_53),
.B1(n_73),
.B2(n_84),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_73),
.B1(n_71),
.B2(n_58),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_149),
.B1(n_100),
.B2(n_97),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_71),
.B(n_1),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_141),
.B(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_114),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_20),
.B(n_29),
.C(n_35),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_148),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_81),
.B1(n_77),
.B2(n_74),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_151),
.B(n_102),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_106),
.A2(n_42),
.B1(n_43),
.B2(n_40),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_166),
.C(n_169),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_109),
.B1(n_100),
.B2(n_123),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_160),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_172),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_171),
.B1(n_177),
.B2(n_133),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_153),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_145),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_116),
.C(n_103),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_97),
.B1(n_122),
.B2(n_99),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_148),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_101),
.C(n_99),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_183),
.B(n_136),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_131),
.A2(n_101),
.B1(n_49),
.B2(n_33),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_49),
.C(n_27),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_143),
.C(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_27),
.B1(n_19),
.B2(n_46),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_147),
.B1(n_27),
.B2(n_35),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_144),
.B(n_9),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_182),
.B(n_184),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_27),
.B(n_1),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_137),
.B(n_27),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_153),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_195),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_129),
.C(n_150),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_189),
.B(n_7),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_190),
.A2(n_210),
.B1(n_156),
.B2(n_161),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_180),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_179),
.A2(n_130),
.B1(n_128),
.B2(n_142),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_200),
.A2(n_211),
.B1(n_174),
.B2(n_156),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_205),
.C(n_207),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_202),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_203),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_125),
.C(n_149),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_143),
.B(n_137),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_209),
.B(n_162),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_141),
.C(n_138),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_141),
.C(n_128),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_189),
.C(n_207),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_35),
.B1(n_7),
.B2(n_10),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_221),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_159),
.B1(n_171),
.B2(n_158),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_220),
.B1(n_228),
.B2(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_232),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_223),
.C(n_205),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_158),
.B1(n_174),
.B2(n_162),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_170),
.C(n_183),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_198),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_236),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_208),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_230),
.B(n_233),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_7),
.B(n_14),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_231),
.B(n_204),
.Y(n_240)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_6),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_234),
.B(n_237),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_200),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_240),
.A2(n_244),
.B1(n_231),
.B2(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_251),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

AOI211xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_212),
.B(n_187),
.C(n_194),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_226),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_245),
.B(n_248),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_254),
.B1(n_220),
.B2(n_236),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_190),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_223),
.Y(n_266)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_188),
.C(n_186),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_257),
.C(n_230),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_186),
.C(n_211),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_259),
.B(n_263),
.Y(n_283)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_273),
.C(n_268),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_272),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_233),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_247),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_213),
.C(n_235),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_270),
.C(n_273),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_213),
.C(n_10),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_239),
.A2(n_16),
.B1(n_13),
.B2(n_12),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_274),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_16),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_16),
.C(n_11),
.Y(n_273)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_244),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_280),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_259),
.A2(n_258),
.B(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_278),
.B(n_279),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_261),
.C(n_265),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_238),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_281),
.B(n_282),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_257),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_255),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_261),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_253),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_288),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_260),
.B1(n_267),
.B2(n_249),
.Y(n_289)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_282),
.A2(n_276),
.B1(n_283),
.B2(n_288),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_292),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_284),
.C(n_277),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_296),
.C(n_3),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_247),
.B1(n_11),
.B2(n_10),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_295),
.B(n_3),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_0),
.C(n_1),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_0),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_299),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_2),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_307),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_4),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_310),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_297),
.C(n_293),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_311),
.A2(n_306),
.B(n_305),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g312 ( 
.A1(n_304),
.A2(n_290),
.B(n_4),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_303),
.C(n_302),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_316),
.C(n_314),
.Y(n_318)
);

O2A1O1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_317),
.B(n_313),
.C(n_309),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_4),
.B(n_5),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_4),
.B1(n_5),
.B2(n_245),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_5),
.Y(n_322)
);


endmodule