module fake_netlist_1_7113_n_936 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_936);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_936;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_624;
wire n_255;
wire n_426;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_241;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_235;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_622;
wire n_549;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_58), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_15), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_64), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_98), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_107), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_78), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_80), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_23), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_53), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_50), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_81), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_97), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_51), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_28), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_19), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_49), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_22), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_45), .Y(n_131) );
CKINVDCx14_ASAP7_75t_R g132 ( .A(n_44), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_96), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_108), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_41), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_59), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_25), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_38), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_12), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_54), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_13), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_11), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_12), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_43), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_109), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_88), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_84), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_37), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_23), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_71), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_14), .Y(n_152) );
INVx1_ASAP7_75t_SL g153 ( .A(n_77), .Y(n_153) );
BUFx3_ASAP7_75t_L g154 ( .A(n_5), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_15), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_99), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_63), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_132), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_127), .B(n_0), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_113), .Y(n_160) );
INVxp67_ASAP7_75t_L g161 ( .A(n_154), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_154), .B(n_0), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_127), .B(n_1), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_154), .B(n_1), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_128), .Y(n_165) );
INVx2_ASAP7_75t_SL g166 ( .A(n_115), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
BUFx12f_ASAP7_75t_L g168 ( .A(n_128), .Y(n_168) );
INVx5_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_115), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_115), .B(n_2), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_128), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_131), .B(n_2), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_128), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_119), .Y(n_177) );
BUFx12f_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_131), .B(n_3), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_117), .B(n_3), .Y(n_180) );
NOR2xp33_ASAP7_75t_SL g181 ( .A(n_153), .B(n_147), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_171), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_158), .B(n_120), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_158), .A2(n_138), .B1(n_140), .B2(n_143), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_171), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_170), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_158), .A2(n_162), .B1(n_164), .B2(n_171), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_162), .A2(n_145), .B1(n_130), .B2(n_144), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_161), .B(n_126), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_162), .A2(n_150), .B1(n_152), .B2(n_155), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_162), .A2(n_155), .B1(n_137), .B2(n_133), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_162), .A2(n_137), .B1(n_122), .B2(n_135), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_161), .B(n_117), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_159), .A2(n_149), .B1(n_114), .B2(n_142), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_171), .B(n_124), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_170), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_171), .A2(n_114), .B1(n_142), .B2(n_124), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_159), .A2(n_114), .B1(n_142), .B2(n_129), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_170), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_159), .B(n_114), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_161), .B(n_129), .Y(n_201) );
OA22x2_ASAP7_75t_L g202 ( .A1(n_171), .A2(n_139), .B1(n_141), .B2(n_148), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_171), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
AO22x2_ASAP7_75t_L g205 ( .A1(n_162), .A2(n_139), .B1(n_141), .B2(n_148), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_166), .B(n_168), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_164), .Y(n_207) );
OAI22xp5_ASAP7_75t_SL g208 ( .A1(n_177), .A2(n_114), .B1(n_142), .B2(n_156), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_177), .B(n_164), .Y(n_209) );
BUFx10_ASAP7_75t_L g210 ( .A(n_164), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_177), .B(n_114), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_166), .B(n_147), .Y(n_212) );
AO22x2_ASAP7_75t_L g213 ( .A1(n_164), .A2(n_156), .B1(n_5), .B2(n_6), .Y(n_213) );
OAI22xp5_ASAP7_75t_SL g214 ( .A1(n_160), .A2(n_142), .B1(n_156), .B2(n_151), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_164), .A2(n_142), .B1(n_157), .B2(n_146), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_164), .A2(n_136), .B1(n_125), .B2(n_123), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_181), .A2(n_121), .B1(n_118), .B2(n_116), .Y(n_217) );
OAI22xp33_ASAP7_75t_R g218 ( .A1(n_180), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_218) );
OR2x6_ASAP7_75t_L g219 ( .A(n_163), .B(n_134), .Y(n_219) );
OAI22xp33_ASAP7_75t_L g220 ( .A1(n_163), .A2(n_134), .B1(n_7), .B2(n_8), .Y(n_220) );
AO22x2_ASAP7_75t_L g221 ( .A1(n_166), .A2(n_4), .B1(n_8), .B2(n_9), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_170), .Y(n_222) );
OAI22xp5_ASAP7_75t_SL g223 ( .A1(n_160), .A2(n_134), .B1(n_10), .B2(n_11), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_181), .A2(n_134), .B1(n_10), .B2(n_13), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_181), .A2(n_9), .B1(n_14), .B2(n_16), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_168), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_180), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_166), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_182), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_182), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_204), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_228), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_185), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_219), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_203), .Y(n_235) );
NOR2xp33_ASAP7_75t_SL g236 ( .A(n_209), .B(n_163), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_207), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_189), .B(n_173), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_187), .B(n_173), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_213), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_210), .Y(n_241) );
INVx4_ASAP7_75t_SL g242 ( .A(n_219), .Y(n_242) );
NAND2x1p5_ASAP7_75t_L g243 ( .A(n_195), .B(n_170), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_192), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_183), .B(n_173), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_213), .Y(n_246) );
AND2x2_ASAP7_75t_SL g247 ( .A(n_195), .B(n_179), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_200), .B(n_179), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_213), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_219), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_186), .Y(n_252) );
XNOR2x2_ASAP7_75t_L g253 ( .A(n_221), .B(n_179), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_196), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_199), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_222), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_202), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_202), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_205), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_205), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_205), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_212), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_212), .Y(n_263) );
INVx4_ASAP7_75t_L g264 ( .A(n_226), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_197), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_226), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_197), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_193), .B(n_176), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_221), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_221), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_206), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_193), .Y(n_272) );
XOR2xp5_ASAP7_75t_L g273 ( .A(n_191), .B(n_17), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_201), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_184), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_201), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_190), .B(n_176), .Y(n_277) );
XNOR2x2_ASAP7_75t_L g278 ( .A(n_227), .B(n_167), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_206), .B(n_176), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_211), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_188), .B(n_176), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_215), .A2(n_176), .B(n_167), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_198), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g284 ( .A1(n_216), .A2(n_167), .B(n_169), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_220), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_220), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_217), .B(n_168), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_208), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_198), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_225), .B(n_18), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_214), .B(n_168), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_224), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_223), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_194), .B(n_19), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_260), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_284), .A2(n_167), .B(n_194), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_242), .B(n_20), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_242), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_243), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_247), .B(n_168), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_247), .B(n_239), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_238), .B(n_20), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_242), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_247), .B(n_178), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_239), .B(n_178), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_238), .B(n_21), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_243), .Y(n_307) );
INVx4_ASAP7_75t_L g308 ( .A(n_242), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_243), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_234), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_254), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_245), .B(n_21), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_231), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_254), .Y(n_314) );
AND2x4_ASAP7_75t_SL g315 ( .A(n_260), .B(n_218), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_254), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_272), .A2(n_167), .B(n_169), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_260), .B(n_178), .Y(n_318) );
INVxp33_ASAP7_75t_L g319 ( .A(n_248), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_242), .B(n_22), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_277), .B(n_178), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_229), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_277), .B(n_24), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_259), .B(n_24), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_277), .B(n_25), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_272), .B(n_178), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_277), .B(n_26), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_274), .B(n_26), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_274), .B(n_27), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_294), .B(n_27), .Y(n_330) );
AND2x2_ASAP7_75t_SL g331 ( .A(n_259), .B(n_165), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_234), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_276), .B(n_262), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_234), .Y(n_334) );
INVx4_ASAP7_75t_L g335 ( .A(n_250), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_294), .B(n_28), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_250), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_229), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_294), .B(n_29), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_294), .B(n_29), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_231), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_290), .B(n_30), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_230), .Y(n_343) );
NAND2x1p5_ASAP7_75t_L g344 ( .A(n_261), .B(n_169), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_230), .Y(n_345) );
AND2x2_ASAP7_75t_SL g346 ( .A(n_261), .B(n_165), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_290), .B(n_30), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_232), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_250), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_348), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_348), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_348), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_348), .Y(n_353) );
OR2x6_ASAP7_75t_L g354 ( .A(n_308), .B(n_240), .Y(n_354) );
OR2x6_ASAP7_75t_SL g355 ( .A(n_328), .B(n_269), .Y(n_355) );
AND2x6_ASAP7_75t_L g356 ( .A(n_298), .B(n_240), .Y(n_356) );
AND2x6_ASAP7_75t_L g357 ( .A(n_298), .B(n_246), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_348), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_297), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_348), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_313), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_333), .B(n_276), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_319), .B(n_236), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_295), .Y(n_364) );
CKINVDCx8_ASAP7_75t_R g365 ( .A(n_297), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_308), .Y(n_366) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_308), .B(n_264), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_319), .B(n_342), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_299), .Y(n_369) );
BUFx2_ASAP7_75t_SL g370 ( .A(n_308), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_313), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_333), .B(n_293), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_319), .B(n_273), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_333), .B(n_293), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_333), .B(n_262), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_313), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_342), .B(n_281), .Y(n_377) );
CKINVDCx8_ASAP7_75t_R g378 ( .A(n_297), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_342), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_295), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_301), .B(n_302), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_313), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_341), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_379), .A2(n_273), .B1(n_347), .B2(n_342), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_350), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_366), .Y(n_386) );
INVx2_ASAP7_75t_SL g387 ( .A(n_366), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_366), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_359), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_350), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_353), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_353), .Y(n_392) );
BUFx12f_ASAP7_75t_L g393 ( .A(n_366), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_351), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_353), .Y(n_395) );
INVx6_ASAP7_75t_L g396 ( .A(n_366), .Y(n_396) );
BUFx8_ASAP7_75t_L g397 ( .A(n_359), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_366), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_351), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_366), .Y(n_400) );
BUFx8_ASAP7_75t_L g401 ( .A(n_352), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_358), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_362), .B(n_301), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_362), .B(n_301), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_358), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_352), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_358), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_360), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_360), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_360), .B(n_308), .Y(n_410) );
CKINVDCx11_ASAP7_75t_R g411 ( .A(n_365), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_361), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_365), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_401), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g415 ( .A1(n_384), .A2(n_365), .B1(n_378), .B2(n_375), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_385), .Y(n_416) );
AOI22xp33_ASAP7_75t_SL g417 ( .A1(n_401), .A2(n_315), .B1(n_347), .B2(n_342), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_385), .Y(n_418) );
INVx4_ASAP7_75t_L g419 ( .A(n_393), .Y(n_419) );
CKINVDCx11_ASAP7_75t_R g420 ( .A(n_393), .Y(n_420) );
NAND2x1p5_ASAP7_75t_L g421 ( .A(n_410), .B(n_369), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_395), .Y(n_422) );
CKINVDCx11_ASAP7_75t_R g423 ( .A(n_393), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_401), .A2(n_315), .B1(n_290), .B2(n_347), .Y(n_424) );
OAI22xp5_ASAP7_75t_SL g425 ( .A1(n_384), .A2(n_244), .B1(n_378), .B2(n_373), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_390), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_392), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_390), .B(n_368), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_394), .Y(n_429) );
INVx6_ASAP7_75t_L g430 ( .A(n_401), .Y(n_430) );
BUFx8_ASAP7_75t_SL g431 ( .A(n_389), .Y(n_431) );
INVx6_ASAP7_75t_L g432 ( .A(n_401), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_394), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_395), .A2(n_375), .B(n_249), .Y(n_434) );
INVx6_ASAP7_75t_L g435 ( .A(n_397), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_399), .Y(n_436) );
INVx8_ASAP7_75t_L g437 ( .A(n_410), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_413), .A2(n_378), .B1(n_355), .B2(n_381), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_397), .Y(n_439) );
BUFx4f_ASAP7_75t_SL g440 ( .A(n_397), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_392), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_403), .B(n_381), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_392), .Y(n_443) );
CKINVDCx6p67_ASAP7_75t_R g444 ( .A(n_411), .Y(n_444) );
CKINVDCx11_ASAP7_75t_R g445 ( .A(n_411), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_386), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_386), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_397), .A2(n_315), .B1(n_290), .B2(n_347), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_399), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_403), .A2(n_315), .B1(n_347), .B2(n_377), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_397), .A2(n_315), .B1(n_327), .B2(n_323), .Y(n_451) );
OAI22x1_ASAP7_75t_L g452 ( .A1(n_406), .A2(n_297), .B1(n_330), .B2(n_336), .Y(n_452) );
AOI22xp33_ASAP7_75t_SL g453 ( .A1(n_389), .A2(n_315), .B1(n_253), .B2(n_325), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_406), .B(n_368), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_389), .A2(n_327), .B1(n_323), .B2(n_325), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_392), .Y(n_456) );
BUFx12f_ASAP7_75t_L g457 ( .A(n_413), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_404), .A2(n_327), .B1(n_323), .B2(n_325), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_427), .Y(n_459) );
BUFx12f_ASAP7_75t_L g460 ( .A(n_420), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_430), .A2(n_432), .B1(n_414), .B2(n_438), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_427), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_415), .A2(n_325), .B1(n_327), .B2(n_323), .Y(n_463) );
OAI21xp5_ASAP7_75t_SL g464 ( .A1(n_417), .A2(n_336), .B(n_330), .Y(n_464) );
INVxp67_ASAP7_75t_L g465 ( .A(n_431), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_423), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_445), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_415), .A2(n_325), .B1(n_327), .B2(n_323), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_430), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_440), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_416), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_430), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_440), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_438), .A2(n_278), .B1(n_297), .B2(n_377), .Y(n_474) );
OAI22xp33_ASAP7_75t_L g475 ( .A1(n_450), .A2(n_355), .B1(n_373), .B2(n_404), .Y(n_475) );
BUFx8_ASAP7_75t_SL g476 ( .A(n_414), .Y(n_476) );
OAI21xp33_ASAP7_75t_L g477 ( .A1(n_453), .A2(n_336), .B(n_330), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_417), .A2(n_340), .B1(n_339), .B2(n_336), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_424), .A2(n_355), .B1(n_330), .B2(n_339), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_430), .A2(n_253), .B1(n_370), .B2(n_330), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_427), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_430), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_441), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_441), .B(n_391), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_441), .B(n_391), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_425), .A2(n_340), .B1(n_339), .B2(n_336), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_425), .A2(n_278), .B1(n_297), .B2(n_339), .Y(n_487) );
OAI21xp5_ASAP7_75t_SL g488 ( .A1(n_414), .A2(n_340), .B(n_339), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_432), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_453), .A2(n_297), .B1(n_340), .B2(n_320), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_414), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_416), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_448), .A2(n_297), .B1(n_340), .B2(n_320), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_418), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_451), .A2(n_297), .B1(n_320), .B2(n_363), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_428), .B(n_412), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_446), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_418), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_432), .A2(n_320), .B1(n_335), .B2(n_410), .Y(n_499) );
OA222x2_ASAP7_75t_L g500 ( .A1(n_439), .A2(n_354), .B1(n_412), .B2(n_249), .C1(n_246), .C2(n_270), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_422), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_426), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_443), .B(n_391), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_443), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_432), .A2(n_320), .B1(n_335), .B2(n_410), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_432), .A2(n_370), .B1(n_396), .B2(n_302), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_439), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_426), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_455), .A2(n_369), .B1(n_410), .B2(n_328), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_443), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_450), .A2(n_335), .B1(n_302), .B2(n_306), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_439), .A2(n_335), .B1(n_302), .B2(n_306), .Y(n_512) );
OAI21xp33_ASAP7_75t_L g513 ( .A1(n_452), .A2(n_329), .B(n_328), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_458), .A2(n_369), .B1(n_328), .B2(n_329), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_435), .A2(n_335), .B1(n_306), .B2(n_302), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_435), .A2(n_396), .B1(n_306), .B2(n_356), .Y(n_516) );
INVx4_ASAP7_75t_L g517 ( .A(n_435), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_435), .A2(n_329), .B1(n_383), .B2(n_371), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_435), .A2(n_335), .B1(n_306), .B2(n_372), .Y(n_519) );
INVx2_ASAP7_75t_SL g520 ( .A(n_437), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_419), .A2(n_329), .B1(n_383), .B2(n_371), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_456), .B(n_386), .Y(n_522) );
OAI21xp5_ASAP7_75t_SL g523 ( .A1(n_421), .A2(n_298), .B(n_312), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_444), .A2(n_335), .B1(n_374), .B2(n_372), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_429), .Y(n_525) );
OAI21xp33_ASAP7_75t_L g526 ( .A1(n_452), .A2(n_433), .B(n_429), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_444), .A2(n_335), .B1(n_374), .B2(n_285), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_419), .A2(n_382), .B1(n_376), .B2(n_361), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_444), .A2(n_335), .B1(n_286), .B2(n_285), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_419), .A2(n_382), .B1(n_376), .B2(n_354), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_419), .A2(n_354), .B1(n_408), .B2(n_407), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_456), .B(n_402), .Y(n_532) );
OAI221xp5_ASAP7_75t_SL g533 ( .A1(n_488), .A2(n_312), .B1(n_286), .B2(n_433), .C(n_436), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_489), .A2(n_437), .B1(n_457), .B2(n_421), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_475), .A2(n_452), .B1(n_437), .B2(n_454), .Y(n_535) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_489), .A2(n_437), .B1(n_457), .B2(n_421), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_489), .A2(n_437), .B1(n_457), .B2(n_421), .Y(n_537) );
AOI22xp33_ASAP7_75t_SL g538 ( .A1(n_489), .A2(n_517), .B1(n_520), .B2(n_472), .Y(n_538) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_517), .A2(n_437), .B1(n_449), .B2(n_436), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_477), .A2(n_428), .B1(n_454), .B2(n_442), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_477), .A2(n_442), .B1(n_356), .B2(n_357), .Y(n_541) );
AOI221xp5_ASAP7_75t_L g542 ( .A1(n_479), .A2(n_449), .B1(n_312), .B2(n_281), .C(n_321), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_517), .A2(n_422), .B1(n_396), .B2(n_388), .Y(n_543) );
NAND2xp33_ASAP7_75t_SL g544 ( .A(n_470), .B(n_456), .Y(n_544) );
NAND2xp33_ASAP7_75t_R g545 ( .A(n_466), .B(n_31), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_471), .B(n_446), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_461), .A2(n_357), .B1(n_356), .B2(n_354), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_517), .A2(n_396), .B1(n_398), .B2(n_388), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_474), .A2(n_357), .B1(n_356), .B2(n_354), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_487), .A2(n_357), .B1(n_356), .B2(n_354), .Y(n_550) );
OAI221xp5_ASAP7_75t_SL g551 ( .A1(n_488), .A2(n_312), .B1(n_301), .B2(n_269), .C(n_270), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_463), .A2(n_468), .B1(n_490), .B2(n_480), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_520), .A2(n_396), .B1(n_388), .B2(n_386), .Y(n_553) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_523), .B(n_408), .C(n_407), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_496), .B(n_409), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_486), .A2(n_356), .B1(n_357), .B2(n_324), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_486), .A2(n_356), .B1(n_357), .B2(n_324), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_509), .A2(n_356), .B1(n_357), .B2(n_324), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_511), .A2(n_356), .B1(n_357), .B2(n_324), .Y(n_559) );
AOI222xp33_ASAP7_75t_L g560 ( .A1(n_460), .A2(n_312), .B1(n_324), .B2(n_409), .C1(n_275), .C2(n_288), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_472), .A2(n_357), .B1(n_324), .B2(n_396), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_472), .A2(n_324), .B1(n_434), .B2(n_387), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_524), .A2(n_324), .B1(n_434), .B2(n_387), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_464), .A2(n_405), .B1(n_402), .B2(n_324), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_523), .B(n_388), .C(n_386), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_464), .A2(n_400), .B1(n_387), .B2(n_405), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_515), .A2(n_400), .B1(n_388), .B2(n_398), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_471), .B(n_402), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_499), .A2(n_400), .B1(n_386), .B2(n_398), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_505), .A2(n_388), .B1(n_386), .B2(n_398), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_527), .A2(n_388), .B1(n_386), .B2(n_398), .Y(n_571) );
OAI222xp33_ASAP7_75t_L g572 ( .A1(n_507), .A2(n_405), .B1(n_308), .B2(n_298), .C1(n_367), .C2(n_303), .Y(n_572) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_465), .B(n_321), .C(n_258), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_478), .A2(n_398), .B1(n_388), .B2(n_308), .Y(n_574) );
NAND3xp33_ASAP7_75t_SL g575 ( .A(n_466), .B(n_308), .C(n_367), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_519), .A2(n_398), .B1(n_349), .B2(n_308), .Y(n_576) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_469), .A2(n_398), .B1(n_446), .B2(n_447), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_514), .A2(n_349), .B1(n_299), .B2(n_309), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_512), .A2(n_349), .B1(n_299), .B2(n_309), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_492), .B(n_446), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_493), .A2(n_349), .B1(n_299), .B2(n_309), .Y(n_581) );
INVx4_ASAP7_75t_L g582 ( .A(n_476), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_513), .A2(n_349), .B1(n_299), .B2(n_309), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_513), .A2(n_307), .B1(n_299), .B2(n_309), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_478), .A2(n_321), .B1(n_309), .B2(n_307), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_518), .A2(n_307), .B1(n_341), .B2(n_305), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_530), .A2(n_307), .B1(n_310), .B2(n_332), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_469), .A2(n_307), .B1(n_310), .B2(n_332), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g589 ( .A1(n_506), .A2(n_267), .B1(n_265), .B2(n_305), .C(n_280), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_469), .A2(n_482), .B1(n_516), .B2(n_529), .Y(n_590) );
OAI21xp5_ASAP7_75t_SL g591 ( .A1(n_531), .A2(n_303), .B(n_367), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_492), .B(n_446), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_501), .B(n_175), .C(n_174), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_522), .Y(n_594) );
NOR2xp67_ASAP7_75t_L g595 ( .A(n_482), .B(n_446), .Y(n_595) );
OAI211xp5_ASAP7_75t_L g596 ( .A1(n_491), .A2(n_303), .B(n_265), .C(n_267), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_494), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_482), .A2(n_307), .B1(n_332), .B2(n_310), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_495), .A2(n_331), .B1(n_346), .B2(n_447), .Y(n_599) );
INVx4_ASAP7_75t_L g600 ( .A(n_460), .Y(n_600) );
OAI211xp5_ASAP7_75t_L g601 ( .A1(n_526), .A2(n_305), .B(n_289), .C(n_282), .Y(n_601) );
OAI221xp5_ASAP7_75t_L g602 ( .A1(n_526), .A2(n_280), .B1(n_257), .B2(n_258), .C(n_289), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_528), .A2(n_332), .B1(n_310), .B2(n_334), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_521), .A2(n_332), .B1(n_310), .B2(n_334), .Y(n_604) );
AOI22xp33_ASAP7_75t_SL g605 ( .A1(n_473), .A2(n_447), .B1(n_331), .B2(n_346), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_494), .A2(n_332), .B1(n_310), .B2(n_334), .Y(n_606) );
NAND3xp33_ASAP7_75t_SL g607 ( .A(n_467), .B(n_31), .C(n_32), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_498), .A2(n_257), .B1(n_280), .B2(n_174), .C(n_175), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_498), .A2(n_332), .B1(n_310), .B2(n_337), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_502), .A2(n_332), .B1(n_310), .B2(n_337), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_502), .A2(n_332), .B1(n_310), .B2(n_337), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_508), .A2(n_447), .B1(n_331), .B2(n_346), .Y(n_612) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_467), .A2(n_447), .B1(n_337), .B2(n_341), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_508), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_525), .A2(n_447), .B1(n_331), .B2(n_346), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_525), .A2(n_331), .B1(n_346), .B2(n_341), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_522), .A2(n_337), .B1(n_296), .B2(n_346), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_532), .B(n_32), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_522), .A2(n_296), .B1(n_346), .B2(n_331), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_484), .B(n_33), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_497), .A2(n_296), .B1(n_331), .B2(n_283), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_459), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_497), .A2(n_296), .B1(n_283), .B2(n_318), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_484), .A2(n_318), .B1(n_345), .B2(n_322), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_497), .A2(n_296), .B1(n_283), .B2(n_318), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_462), .Y(n_626) );
NAND2xp33_ASAP7_75t_SL g627 ( .A(n_485), .B(n_295), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_485), .A2(n_296), .B1(n_283), .B2(n_291), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_497), .A2(n_345), .B1(n_343), .B2(n_338), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_503), .B(n_33), .Y(n_630) );
OAI21xp33_ASAP7_75t_L g631 ( .A1(n_503), .A2(n_165), .B(n_172), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_532), .B(n_34), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_462), .A2(n_343), .B1(n_338), .B2(n_345), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_481), .B(n_34), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_600), .B(n_35), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_545), .A2(n_510), .B1(n_504), .B2(n_483), .C(n_481), .Y(n_636) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_534), .A2(n_500), .B(n_483), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_535), .A2(n_500), .B1(n_345), .B2(n_322), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_554), .A2(n_165), .B(n_172), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_597), .B(n_35), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_597), .B(n_36), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_614), .B(n_36), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_614), .B(n_37), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_560), .B(n_165), .C(n_175), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_546), .B(n_165), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_555), .B(n_38), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_560), .B(n_165), .C(n_175), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_632), .B(n_39), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_593), .B(n_165), .C(n_175), .Y(n_649) );
NOR3xp33_ASAP7_75t_L g650 ( .A(n_607), .B(n_317), .C(n_292), .Y(n_650) );
NAND3xp33_ASAP7_75t_L g651 ( .A(n_593), .B(n_165), .C(n_175), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_536), .A2(n_311), .B1(n_314), .B2(n_316), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_546), .B(n_580), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_554), .B(n_364), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_580), .B(n_39), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_565), .B(n_364), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_592), .B(n_40), .Y(n_657) );
OAI221xp5_ASAP7_75t_SL g658 ( .A1(n_552), .A2(n_292), .B1(n_300), .B2(n_304), .C(n_338), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_592), .B(n_165), .Y(n_659) );
NOR3xp33_ASAP7_75t_L g660 ( .A(n_575), .B(n_317), .C(n_268), .Y(n_660) );
NAND4xp25_ASAP7_75t_L g661 ( .A(n_590), .B(n_304), .C(n_300), .D(n_317), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_573), .A2(n_172), .B1(n_174), .B2(n_175), .C(n_169), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_565), .B(n_172), .C(n_175), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_594), .B(n_172), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_540), .B(n_40), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_594), .B(n_172), .Y(n_666) );
OAI221xp5_ASAP7_75t_SL g667 ( .A1(n_591), .A2(n_300), .B1(n_304), .B2(n_322), .C(n_338), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_564), .A2(n_322), .B1(n_345), .B2(n_338), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_591), .B(n_172), .C(n_175), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_564), .A2(n_322), .B1(n_345), .B2(n_338), .Y(n_670) );
AND2x2_ASAP7_75t_SL g671 ( .A(n_582), .B(n_295), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_626), .B(n_172), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_538), .B(n_172), .C(n_175), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_533), .A2(n_174), .B1(n_169), .B2(n_317), .C(n_263), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_634), .B(n_174), .C(n_169), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_600), .B(n_582), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_626), .B(n_41), .Y(n_677) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_618), .B(n_174), .C(n_169), .Y(n_678) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_566), .A2(n_311), .B1(n_314), .B2(n_316), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_620), .B(n_630), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_539), .B(n_174), .C(n_169), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_622), .B(n_42), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_622), .B(n_174), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_549), .A2(n_322), .B1(n_343), .B2(n_174), .Y(n_684) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_600), .B(n_263), .C(n_343), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g686 ( .A(n_537), .B(n_601), .C(n_583), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_550), .A2(n_343), .B1(n_174), .B2(n_311), .Y(n_687) );
OAI21xp5_ASAP7_75t_SL g688 ( .A1(n_547), .A2(n_344), .B(n_300), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_551), .A2(n_169), .B1(n_233), .B2(n_304), .C(n_343), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_541), .A2(n_311), .B1(n_316), .B2(n_314), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_568), .B(n_42), .Y(n_691) );
OA21x2_ASAP7_75t_L g692 ( .A1(n_631), .A2(n_380), .B(n_364), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_582), .A2(n_344), .B1(n_233), .B2(n_169), .C(n_326), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_586), .B(n_43), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_586), .B(n_44), .Y(n_695) );
OAI21xp33_ASAP7_75t_SL g696 ( .A1(n_595), .A2(n_380), .B(n_46), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_543), .B(n_311), .C(n_316), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_595), .B(n_45), .Y(n_698) );
NOR3xp33_ASAP7_75t_L g699 ( .A(n_589), .B(n_326), .C(n_287), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_544), .B(n_380), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_584), .B(n_577), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_628), .B(n_46), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_548), .B(n_47), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_585), .A2(n_316), .B1(n_314), .B2(n_311), .Y(n_704) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_631), .A2(n_316), .B(n_314), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_553), .B(n_47), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_542), .A2(n_314), .B1(n_295), .B2(n_344), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_570), .B(n_48), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_569), .B(n_295), .C(n_255), .Y(n_709) );
AND2x2_ASAP7_75t_SL g710 ( .A(n_558), .B(n_295), .Y(n_710) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_596), .B(n_295), .C(n_255), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_571), .B(n_52), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_556), .A2(n_295), .B1(n_344), .B2(n_256), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_557), .A2(n_295), .B1(n_344), .B2(n_256), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g715 ( .A(n_567), .B(n_295), .C(n_252), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_562), .B(n_295), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_624), .B(n_55), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g718 ( .A(n_613), .B(n_326), .C(n_232), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_608), .B(n_295), .C(n_252), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_633), .B(n_295), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_624), .B(n_56), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_605), .A2(n_344), .B1(n_326), .B2(n_271), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_633), .B(n_57), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_559), .A2(n_344), .B1(n_271), .B2(n_251), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_563), .A2(n_574), .B1(n_576), .B2(n_578), .Y(n_725) );
NAND3xp33_ASAP7_75t_L g726 ( .A(n_544), .B(n_237), .C(n_235), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_585), .B(n_60), .Y(n_727) );
OAI21xp5_ASAP7_75t_SL g728 ( .A1(n_572), .A2(n_251), .B(n_279), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_623), .B(n_61), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_587), .B(n_62), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_625), .B(n_65), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_604), .B(n_66), .Y(n_732) );
AOI21xp5_ASAP7_75t_SL g733 ( .A1(n_599), .A2(n_67), .B(n_68), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_629), .B(n_69), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_561), .B(n_70), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_617), .B(n_72), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_603), .B(n_73), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_621), .B(n_74), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_627), .B(n_271), .Y(n_739) );
NOR3xp33_ASAP7_75t_SL g740 ( .A(n_637), .B(n_627), .C(n_599), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_636), .B(n_602), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_653), .B(n_579), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_685), .B(n_598), .C(n_588), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_653), .B(n_606), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_645), .B(n_581), .Y(n_745) );
NAND3xp33_ASAP7_75t_L g746 ( .A(n_669), .B(n_610), .C(n_609), .Y(n_746) );
AOI211xp5_ASAP7_75t_L g747 ( .A1(n_635), .A2(n_615), .B(n_612), .C(n_616), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_659), .B(n_611), .Y(n_748) );
INVx1_ASAP7_75t_SL g749 ( .A(n_676), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_686), .B(n_619), .C(n_237), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_644), .A2(n_235), .B1(n_241), .B2(n_266), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_659), .B(n_75), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_655), .B(n_76), .Y(n_753) );
NAND4xp75_ASAP7_75t_L g754 ( .A(n_671), .B(n_696), .C(n_701), .D(n_706), .Y(n_754) );
INVx1_ASAP7_75t_SL g755 ( .A(n_671), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_701), .B(n_82), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_664), .B(n_83), .Y(n_757) );
OR2x2_ASAP7_75t_L g758 ( .A(n_657), .B(n_86), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_647), .A2(n_264), .B1(n_87), .B2(n_89), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_680), .B(n_90), .Y(n_760) );
NAND3xp33_ASAP7_75t_L g761 ( .A(n_696), .B(n_264), .C(n_92), .Y(n_761) );
BUFx2_ASAP7_75t_L g762 ( .A(n_698), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_666), .B(n_91), .Y(n_763) );
NAND3xp33_ASAP7_75t_L g764 ( .A(n_638), .B(n_264), .C(n_94), .Y(n_764) );
NOR3xp33_ASAP7_75t_L g765 ( .A(n_665), .B(n_93), .C(n_95), .Y(n_765) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_673), .B(n_100), .C(n_101), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_661), .A2(n_102), .B1(n_103), .B2(n_104), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_698), .B(n_105), .Y(n_768) );
NAND4xp75_ASAP7_75t_L g769 ( .A(n_706), .B(n_106), .C(n_110), .D(n_111), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_699), .A2(n_112), .B1(n_689), .B2(n_725), .Y(n_770) );
OA211x2_ASAP7_75t_L g771 ( .A1(n_639), .A2(n_700), .B(n_654), .C(n_739), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_640), .B(n_641), .Y(n_772) );
AND2x4_ASAP7_75t_L g773 ( .A(n_656), .B(n_654), .Y(n_773) );
OAI211xp5_ASAP7_75t_L g774 ( .A1(n_728), .A2(n_688), .B(n_733), .C(n_667), .Y(n_774) );
NOR3xp33_ASAP7_75t_L g775 ( .A(n_648), .B(n_646), .C(n_694), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_639), .B(n_663), .Y(n_776) );
INVxp33_ASAP7_75t_L g777 ( .A(n_733), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_642), .B(n_643), .Y(n_778) );
OR2x2_ASAP7_75t_L g779 ( .A(n_656), .B(n_677), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_726), .A2(n_711), .B(n_681), .Y(n_780) );
AOI211x1_ASAP7_75t_L g781 ( .A1(n_693), .A2(n_695), .B(n_703), .C(n_702), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_672), .B(n_682), .Y(n_782) );
OR2x2_ASAP7_75t_L g783 ( .A(n_691), .B(n_683), .Y(n_783) );
OAI211xp5_ASAP7_75t_L g784 ( .A1(n_679), .A2(n_668), .B(n_670), .C(n_658), .Y(n_784) );
OR2x6_ASAP7_75t_L g785 ( .A(n_700), .B(n_739), .Y(n_785) );
AOI21xp33_ASAP7_75t_L g786 ( .A1(n_678), .A2(n_675), .B(n_735), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_717), .B(n_721), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_721), .B(n_736), .Y(n_788) );
BUFx3_ASAP7_75t_L g789 ( .A(n_697), .Y(n_789) );
AND2x4_ASAP7_75t_L g790 ( .A(n_712), .B(n_708), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_727), .B(n_710), .Y(n_791) );
OAI211xp5_ASAP7_75t_SL g792 ( .A1(n_674), .A2(n_662), .B(n_684), .C(n_687), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_705), .B(n_649), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_718), .A2(n_650), .B1(n_710), .B2(n_722), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_736), .B(n_729), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_651), .A2(n_705), .B(n_652), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_738), .A2(n_731), .B1(n_729), .B2(n_660), .Y(n_797) );
NOR3xp33_ASAP7_75t_L g798 ( .A(n_723), .B(n_732), .C(n_737), .Y(n_798) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_724), .A2(n_738), .B1(n_731), .B2(n_704), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_716), .A2(n_708), .B1(n_712), .B2(n_707), .Y(n_800) );
NAND3xp33_ASAP7_75t_L g801 ( .A(n_715), .B(n_709), .C(n_690), .Y(n_801) );
NAND4xp75_ASAP7_75t_L g802 ( .A(n_730), .B(n_734), .C(n_692), .D(n_720), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_719), .B(n_713), .Y(n_803) );
NOR3xp33_ASAP7_75t_L g804 ( .A(n_714), .B(n_607), .C(n_635), .Y(n_804) );
OR2x6_ASAP7_75t_L g805 ( .A(n_637), .B(n_554), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_644), .A2(n_647), .B1(n_560), .B2(n_661), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_653), .B(n_645), .Y(n_807) );
NAND3xp33_ASAP7_75t_L g808 ( .A(n_637), .B(n_636), .C(n_685), .Y(n_808) );
INVx2_ASAP7_75t_SL g809 ( .A(n_676), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_653), .Y(n_810) );
NAND3xp33_ASAP7_75t_SL g811 ( .A(n_637), .B(n_685), .C(n_635), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_653), .Y(n_812) );
NAND4xp75_ASAP7_75t_L g813 ( .A(n_676), .B(n_635), .C(n_671), .D(n_696), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_644), .A2(n_647), .B1(n_560), .B2(n_661), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_810), .B(n_812), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_807), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_762), .B(n_742), .Y(n_817) );
INVx1_ASAP7_75t_SL g818 ( .A(n_749), .Y(n_818) );
INVx2_ASAP7_75t_SL g819 ( .A(n_809), .Y(n_819) );
XNOR2xp5_ASAP7_75t_L g820 ( .A(n_811), .B(n_754), .Y(n_820) );
CKINVDCx16_ASAP7_75t_R g821 ( .A(n_805), .Y(n_821) );
NOR3xp33_ASAP7_75t_L g822 ( .A(n_808), .B(n_774), .C(n_756), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_772), .B(n_778), .Y(n_823) );
AND4x1_ASAP7_75t_L g824 ( .A(n_740), .B(n_814), .C(n_806), .D(n_804), .Y(n_824) );
NAND2xp5_ASAP7_75t_SL g825 ( .A(n_777), .B(n_740), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_805), .B(n_744), .Y(n_826) );
INVx3_ASAP7_75t_L g827 ( .A(n_785), .Y(n_827) );
INVx3_ASAP7_75t_L g828 ( .A(n_785), .Y(n_828) );
OR2x2_ASAP7_75t_L g829 ( .A(n_779), .B(n_783), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_773), .Y(n_830) );
NAND4xp75_ASAP7_75t_L g831 ( .A(n_771), .B(n_781), .C(n_780), .D(n_794), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_773), .Y(n_832) );
NOR3xp33_ASAP7_75t_L g833 ( .A(n_750), .B(n_813), .C(n_804), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_805), .Y(n_834) );
NOR3xp33_ASAP7_75t_SL g835 ( .A(n_784), .B(n_741), .C(n_802), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_747), .B(n_741), .Y(n_836) );
NAND4xp75_ASAP7_75t_SL g837 ( .A(n_777), .B(n_791), .C(n_803), .D(n_768), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_785), .Y(n_838) );
NOR3xp33_ASAP7_75t_L g839 ( .A(n_775), .B(n_786), .C(n_764), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_775), .B(n_782), .Y(n_840) );
XNOR2xp5_ASAP7_75t_L g841 ( .A(n_787), .B(n_814), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_745), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_760), .B(n_755), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_789), .Y(n_844) );
NAND4xp75_ASAP7_75t_SL g845 ( .A(n_791), .B(n_803), .C(n_763), .D(n_757), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_748), .Y(n_846) );
OR2x2_ASAP7_75t_L g847 ( .A(n_788), .B(n_790), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_790), .B(n_795), .Y(n_848) );
XOR2x2_ASAP7_75t_L g849 ( .A(n_806), .B(n_769), .Y(n_849) );
NAND2xp5_ASAP7_75t_SL g850 ( .A(n_789), .B(n_797), .Y(n_850) );
NAND4xp75_ASAP7_75t_SL g851 ( .A(n_770), .B(n_797), .C(n_761), .D(n_767), .Y(n_851) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_776), .Y(n_852) );
BUFx3_ASAP7_75t_L g853 ( .A(n_766), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_800), .B(n_798), .Y(n_854) );
NAND3xp33_ASAP7_75t_L g855 ( .A(n_770), .B(n_776), .C(n_765), .Y(n_855) );
NOR2x1_ASAP7_75t_L g856 ( .A(n_793), .B(n_796), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_793), .Y(n_857) );
INVx1_ASAP7_75t_SL g858 ( .A(n_818), .Y(n_858) );
NOR2x1_ASAP7_75t_L g859 ( .A(n_856), .B(n_801), .Y(n_859) );
XNOR2xp5_ASAP7_75t_L g860 ( .A(n_820), .B(n_800), .Y(n_860) );
XOR2x2_ASAP7_75t_L g861 ( .A(n_820), .B(n_799), .Y(n_861) );
XOR2x2_ASAP7_75t_L g862 ( .A(n_824), .B(n_743), .Y(n_862) );
NOR2x1_ASAP7_75t_L g863 ( .A(n_856), .B(n_746), .Y(n_863) );
INVx2_ASAP7_75t_SL g864 ( .A(n_819), .Y(n_864) );
XOR2x2_ASAP7_75t_L g865 ( .A(n_824), .B(n_765), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_829), .Y(n_866) );
INVx2_ASAP7_75t_SL g867 ( .A(n_819), .Y(n_867) );
INVxp33_ASAP7_75t_L g868 ( .A(n_833), .Y(n_868) );
NOR2x1_ASAP7_75t_L g869 ( .A(n_837), .B(n_753), .Y(n_869) );
XNOR2x1_ASAP7_75t_L g870 ( .A(n_849), .B(n_758), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_829), .Y(n_871) );
INVx1_ASAP7_75t_SL g872 ( .A(n_844), .Y(n_872) );
XNOR2xp5_ASAP7_75t_L g873 ( .A(n_849), .B(n_798), .Y(n_873) );
OA22x2_ASAP7_75t_L g874 ( .A1(n_825), .A2(n_751), .B1(n_752), .B2(n_767), .Y(n_874) );
OA22x2_ASAP7_75t_L g875 ( .A1(n_834), .A2(n_759), .B1(n_792), .B2(n_841), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_815), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_815), .Y(n_877) );
CKINVDCx8_ASAP7_75t_R g878 ( .A(n_821), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_842), .Y(n_879) );
INVxp67_ASAP7_75t_L g880 ( .A(n_852), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_842), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_840), .Y(n_882) );
XNOR2xp5_ASAP7_75t_L g883 ( .A(n_841), .B(n_759), .Y(n_883) );
XNOR2x1_ASAP7_75t_L g884 ( .A(n_831), .B(n_851), .Y(n_884) );
XNOR2xp5_ASAP7_75t_L g885 ( .A(n_831), .B(n_835), .Y(n_885) );
XOR2xp5_ASAP7_75t_L g886 ( .A(n_845), .B(n_821), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_878), .A2(n_834), .B1(n_850), .B2(n_855), .Y(n_887) );
OA22x2_ASAP7_75t_SL g888 ( .A1(n_875), .A2(n_857), .B1(n_838), .B2(n_844), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_875), .A2(n_822), .B1(n_854), .B2(n_839), .Y(n_889) );
XNOR2xp5_ASAP7_75t_L g890 ( .A(n_884), .B(n_885), .Y(n_890) );
OA22x2_ASAP7_75t_L g891 ( .A1(n_873), .A2(n_854), .B1(n_836), .B2(n_826), .Y(n_891) );
AO22x2_ASAP7_75t_L g892 ( .A1(n_858), .A2(n_857), .B1(n_827), .B2(n_828), .Y(n_892) );
INVx2_ASAP7_75t_L g893 ( .A(n_858), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_866), .Y(n_894) );
AO22x2_ASAP7_75t_L g895 ( .A1(n_870), .A2(n_828), .B1(n_827), .B2(n_855), .Y(n_895) );
XOR2x2_ASAP7_75t_L g896 ( .A(n_862), .B(n_823), .Y(n_896) );
BUFx3_ASAP7_75t_L g897 ( .A(n_864), .Y(n_897) );
XOR2x2_ASAP7_75t_L g898 ( .A(n_861), .B(n_817), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_871), .Y(n_899) );
AO22x1_ASAP7_75t_L g900 ( .A1(n_859), .A2(n_828), .B1(n_827), .B2(n_838), .Y(n_900) );
INVx2_ASAP7_75t_L g901 ( .A(n_872), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_876), .Y(n_902) );
HB1xp67_ASAP7_75t_L g903 ( .A(n_893), .Y(n_903) );
INVx2_ASAP7_75t_SL g904 ( .A(n_897), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_901), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_890), .B(n_868), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_901), .Y(n_907) );
OAI322xp33_ASAP7_75t_L g908 ( .A1(n_888), .A2(n_860), .A3(n_880), .B1(n_882), .B2(n_886), .C1(n_883), .C2(n_874), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_889), .A2(n_863), .B1(n_868), .B2(n_880), .Y(n_909) );
AOI322xp5_ASAP7_75t_L g910 ( .A1(n_888), .A2(n_817), .A3(n_869), .B1(n_848), .B2(n_877), .C1(n_867), .C2(n_846), .Y(n_910) );
INVx2_ASAP7_75t_SL g911 ( .A(n_897), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_903), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_903), .Y(n_913) );
OAI22x1_ASAP7_75t_L g914 ( .A1(n_904), .A2(n_895), .B1(n_891), .B2(n_887), .Y(n_914) );
OA22x2_ASAP7_75t_L g915 ( .A1(n_911), .A2(n_887), .B1(n_891), .B2(n_895), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_905), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_915), .A2(n_895), .B1(n_906), .B2(n_909), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_913), .A2(n_906), .B1(n_907), .B2(n_892), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_912), .A2(n_892), .B1(n_874), .B2(n_894), .Y(n_919) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_917), .A2(n_914), .B1(n_865), .B2(n_919), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_918), .Y(n_921) );
AO22x1_ASAP7_75t_L g922 ( .A1(n_917), .A2(n_912), .B1(n_916), .B2(n_908), .Y(n_922) );
INVx2_ASAP7_75t_L g923 ( .A(n_921), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_922), .A2(n_896), .B1(n_898), .B2(n_892), .Y(n_924) );
NAND5xp2_ASAP7_75t_L g925 ( .A(n_924), .B(n_920), .C(n_910), .D(n_843), .E(n_900), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_923), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_926), .B(n_872), .Y(n_927) );
NOR2x1_ASAP7_75t_L g928 ( .A(n_926), .B(n_899), .Y(n_928) );
OAI22xp5_ASAP7_75t_SL g929 ( .A1(n_927), .A2(n_925), .B1(n_828), .B2(n_827), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_929), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g931 ( .A1(n_930), .A2(n_928), .B1(n_902), .B2(n_846), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_931), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_932), .A2(n_830), .B1(n_853), .B2(n_832), .Y(n_933) );
XNOR2xp5_ASAP7_75t_L g934 ( .A(n_933), .B(n_847), .Y(n_934) );
AOI221xp5_ASAP7_75t_L g935 ( .A1(n_934), .A2(n_830), .B1(n_881), .B2(n_879), .C(n_853), .Y(n_935) );
AOI211xp5_ASAP7_75t_L g936 ( .A1(n_935), .A2(n_847), .B(n_816), .C(n_832), .Y(n_936) );
endmodule