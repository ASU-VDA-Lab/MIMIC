module fake_netlist_5_752_n_2067 (n_137, n_294, n_431, n_318, n_380, n_419, n_611, n_444, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_620, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_600, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_489, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2067);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_611;
input n_444;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_600;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2067;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_785;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_1007;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2001;
wire n_1494;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_1939;
wire n_1806;
wire n_933;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_1230;
wire n_668;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2058;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_1078;
wire n_1670;
wire n_775;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_1948;
wire n_1984;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_926;
wire n_1218;
wire n_1931;
wire n_1070;
wire n_777;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_889;
wire n_973;
wire n_1700;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_1403;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_1819;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_857;
wire n_832;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_809;
wire n_870;
wire n_931;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2009;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_1308;
wire n_1767;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_1121;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_959;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_1609;
wire n_1989;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_662;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_700;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_1823;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_860;
wire n_1805;
wire n_1816;
wire n_948;
wire n_1217;
wire n_628;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_1435;
wire n_879;
wire n_824;
wire n_1645;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_815;
wire n_1795;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_803;
wire n_1092;
wire n_1776;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_1958;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_1346;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_912;
wire n_968;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_885;
wire n_1432;
wire n_1357;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_1179;
wire n_753;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_896;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_1174;
wire n_1371;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_679;
wire n_710;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_676;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_1999;
wire n_2065;
wire n_1372;
wire n_1273;
wire n_1822;
wire n_643;
wire n_916;
wire n_1081;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_812;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_1341;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_1842;
wire n_871;
wire n_685;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_1589;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_1937;
wire n_1739;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2027;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1996;
wire n_1879;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_2044;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_1542;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_587),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_379),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_419),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_497),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_518),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_551),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_29),
.Y(n_632)
);

BUFx10_ASAP7_75t_L g633 ( 
.A(n_562),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_31),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_613),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_514),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_327),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_495),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_407),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_147),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_344),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_570),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_325),
.Y(n_643)
);

BUFx10_ASAP7_75t_L g644 ( 
.A(n_383),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_275),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_545),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_395),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_598),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_537),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_136),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_168),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_529),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_585),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_137),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_581),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_285),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_549),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_597),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_600),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_359),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_92),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_566),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_14),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_274),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_313),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_599),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_540),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_575),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_84),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_425),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_611),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_224),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_595),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_197),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_606),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_572),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_618),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_596),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_496),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_42),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_617),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_542),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_356),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_588),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_283),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_165),
.Y(n_686)
);

BUFx5_ASAP7_75t_L g687 ( 
.A(n_458),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_393),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_168),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_57),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_49),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_214),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_141),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_329),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_70),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_557),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_352),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_464),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_412),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_550),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_152),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_126),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_479),
.Y(n_703)
);

CKINVDCx14_ASAP7_75t_R g704 ( 
.A(n_185),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_556),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_213),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_564),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_601),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_589),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_592),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_157),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_81),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_248),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_394),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_355),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_226),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_87),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_610),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_292),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_38),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_420),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_457),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_603),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_530),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_619),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_531),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_415),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_579),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_342),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_424),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_546),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_462),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_280),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_455),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_485),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_594),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_125),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_305),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_243),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_565),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_118),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_605),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_547),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_439),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_364),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_385),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_83),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_405),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_609),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_30),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_474),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_314),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_607),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_471),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_586),
.Y(n_755)
);

CKINVDCx6p67_ASAP7_75t_R g756 ( 
.A(n_590),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_476),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_475),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_442),
.Y(n_759)
);

BUFx2_ASAP7_75t_SL g760 ( 
.A(n_131),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_604),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_558),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_561),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_437),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_583),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_145),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_582),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_130),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_555),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_559),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_573),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_567),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_271),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_608),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_231),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_267),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_602),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_53),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_388),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_59),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_389),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_574),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_54),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_554),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_552),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_332),
.Y(n_786)
);

BUFx8_ASAP7_75t_SL g787 ( 
.A(n_538),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_456),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_568),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_536),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_370),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_463),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_516),
.Y(n_793)
);

CKINVDCx16_ASAP7_75t_R g794 ( 
.A(n_197),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_431),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_204),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_24),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_519),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_539),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_3),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_520),
.Y(n_801)
);

CKINVDCx16_ASAP7_75t_R g802 ( 
.A(n_584),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_491),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_48),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_409),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_226),
.Y(n_806)
);

BUFx5_ASAP7_75t_L g807 ( 
.A(n_505),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_91),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_449),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_612),
.Y(n_810)
);

CKINVDCx16_ASAP7_75t_R g811 ( 
.A(n_367),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_167),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_577),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_19),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_593),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_548),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_371),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_578),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_571),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_500),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_304),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_397),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_157),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_133),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_132),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_184),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_544),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_362),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_553),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_484),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_576),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_102),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_297),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_193),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_396),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_72),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_560),
.Y(n_837)
);

CKINVDCx14_ASAP7_75t_R g838 ( 
.A(n_427),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_398),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_481),
.Y(n_840)
);

CKINVDCx14_ASAP7_75t_R g841 ( 
.A(n_591),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_541),
.Y(n_842)
);

INVxp33_ASAP7_75t_L g843 ( 
.A(n_543),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_151),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_569),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_78),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_369),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_563),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_4),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_580),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_515),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_87),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_402),
.Y(n_853)
);

CKINVDCx16_ASAP7_75t_R g854 ( 
.A(n_794),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_843),
.B(n_1),
.Y(n_855)
);

INVxp33_ASAP7_75t_SL g856 ( 
.A(n_669),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_787),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_773),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_704),
.B(n_0),
.Y(n_859)
);

CKINVDCx16_ASAP7_75t_R g860 ( 
.A(n_802),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_675),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_773),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_665),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_626),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_627),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_628),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_629),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_773),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_636),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_639),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_641),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_747),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_632),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_760),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_630),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_660),
.B(n_1),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_642),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_712),
.B(n_0),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_656),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_875),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_860),
.B(n_811),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_854),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_858),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_862),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_868),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_875),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_864),
.B(n_838),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_865),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_856),
.B(n_730),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_875),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_863),
.B(n_874),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_866),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_867),
.B(n_841),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_869),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_873),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_879),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_870),
.B(n_871),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_878),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_855),
.Y(n_899)
);

OAI21x1_ASAP7_75t_L g900 ( 
.A1(n_859),
.A2(n_637),
.B(n_631),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_877),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_876),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_872),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_857),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_861),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_858),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_891),
.B(n_829),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_901),
.B(n_851),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_880),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_880),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_896),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_899),
.A2(n_739),
.B1(n_741),
.B2(n_713),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_880),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_887),
.B(n_638),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_902),
.A2(n_654),
.B1(n_732),
.B2(n_697),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_890),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_883),
.Y(n_917)
);

INVx4_ASAP7_75t_L g918 ( 
.A(n_894),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_893),
.B(n_897),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_888),
.Y(n_920)
);

NOR3xp33_ASAP7_75t_L g921 ( 
.A(n_889),
.B(n_680),
.C(n_640),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_898),
.B(n_701),
.Y(n_922)
);

INVx4_ASAP7_75t_L g923 ( 
.A(n_905),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_884),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_895),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_885),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_906),
.B(n_647),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_900),
.B(n_655),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_892),
.B(n_822),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_905),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_881),
.B(n_649),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_903),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_904),
.Y(n_933)
);

NAND3x1_ASAP7_75t_L g934 ( 
.A(n_882),
.B(n_674),
.C(n_661),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_905),
.A2(n_825),
.B1(n_852),
.B2(n_768),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_899),
.B(n_758),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_896),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_894),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_886),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_882),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_896),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_891),
.B(n_717),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_896),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_896),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_917),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_944),
.Y(n_946)
);

AO22x2_ASAP7_75t_L g947 ( 
.A1(n_915),
.A2(n_691),
.B1(n_750),
.B2(n_706),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_931),
.A2(n_646),
.B(n_648),
.C(n_643),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_944),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_926),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_926),
.Y(n_951)
);

AO22x2_ASAP7_75t_L g952 ( 
.A1(n_921),
.A2(n_832),
.B1(n_844),
.B2(n_823),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_911),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_920),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_937),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_914),
.A2(n_761),
.B1(n_791),
.B2(n_784),
.Y(n_956)
);

AND2x6_ASAP7_75t_L g957 ( 
.A(n_933),
.B(n_653),
.Y(n_957)
);

OR2x6_ASAP7_75t_L g958 ( 
.A(n_923),
.B(n_693),
.Y(n_958)
);

AO22x2_ASAP7_75t_L g959 ( 
.A1(n_922),
.A2(n_766),
.B1(n_737),
.B2(n_775),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_942),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_907),
.B(n_799),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_941),
.Y(n_962)
);

CKINVDCx16_ASAP7_75t_R g963 ( 
.A(n_940),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_924),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_932),
.B(n_778),
.Y(n_965)
);

OAI221xp5_ASAP7_75t_L g966 ( 
.A1(n_912),
.A2(n_826),
.B1(n_834),
.B2(n_808),
.C(n_800),
.Y(n_966)
);

OAI221xp5_ASAP7_75t_L g967 ( 
.A1(n_936),
.A2(n_752),
.B1(n_762),
.B2(n_731),
.C(n_723),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_943),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_925),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_939),
.Y(n_970)
);

AO22x2_ASAP7_75t_L g971 ( 
.A1(n_934),
.A2(n_681),
.B1(n_694),
.B2(n_670),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_927),
.B(n_916),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_929),
.A2(n_827),
.B1(n_830),
.B2(n_819),
.Y(n_973)
);

AO22x2_ASAP7_75t_L g974 ( 
.A1(n_918),
.A2(n_698),
.B1(n_718),
.B2(n_699),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_938),
.Y(n_975)
);

AO22x2_ASAP7_75t_L g976 ( 
.A1(n_927),
.A2(n_722),
.B1(n_735),
.B2(n_721),
.Y(n_976)
);

NOR2xp67_ASAP7_75t_L g977 ( 
.A(n_909),
.B(n_652),
.Y(n_977)
);

OAI221xp5_ASAP7_75t_L g978 ( 
.A1(n_935),
.A2(n_771),
.B1(n_815),
.B2(n_764),
.C(n_755),
.Y(n_978)
);

INVxp33_ASAP7_75t_L g979 ( 
.A(n_910),
.Y(n_979)
);

OR2x2_ASAP7_75t_SL g980 ( 
.A(n_910),
.B(n_702),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_928),
.A2(n_831),
.B1(n_658),
.B2(n_659),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_928),
.B(n_913),
.Y(n_982)
);

AO22x2_ASAP7_75t_L g983 ( 
.A1(n_913),
.A2(n_740),
.B1(n_744),
.B2(n_736),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_944),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_919),
.A2(n_754),
.B1(n_840),
.B2(n_746),
.Y(n_985)
);

AO22x2_ASAP7_75t_L g986 ( 
.A1(n_915),
.A2(n_749),
.B1(n_753),
.B2(n_748),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_914),
.B(n_769),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_944),
.Y(n_988)
);

OAI221xp5_ASAP7_75t_L g989 ( 
.A1(n_912),
.A2(n_850),
.B1(n_839),
.B2(n_774),
.C(n_779),
.Y(n_989)
);

AO22x2_ASAP7_75t_L g990 ( 
.A1(n_915),
.A2(n_781),
.B1(n_786),
.B2(n_777),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_942),
.B(n_719),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_920),
.Y(n_992)
);

AO22x2_ASAP7_75t_L g993 ( 
.A1(n_915),
.A2(n_793),
.B1(n_805),
.B2(n_792),
.Y(n_993)
);

OAI221xp5_ASAP7_75t_L g994 ( 
.A1(n_912),
.A2(n_842),
.B1(n_820),
.B2(n_817),
.C(n_816),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_944),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_944),
.Y(n_996)
);

OAI221xp5_ASAP7_75t_L g997 ( 
.A1(n_912),
.A2(n_634),
.B1(n_651),
.B2(n_650),
.C(n_645),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_914),
.B(n_662),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_944),
.Y(n_999)
);

BUFx8_ASAP7_75t_L g1000 ( 
.A(n_930),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_944),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_908),
.B(n_848),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_944),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_944),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_920),
.Y(n_1005)
);

INVxp33_ASAP7_75t_SL g1006 ( 
.A(n_920),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_944),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_914),
.B(n_666),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_944),
.Y(n_1009)
);

AO22x2_ASAP7_75t_L g1010 ( 
.A1(n_915),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_944),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_944),
.Y(n_1012)
);

OAI221xp5_ASAP7_75t_L g1013 ( 
.A1(n_912),
.A2(n_672),
.B1(n_685),
.B2(n_664),
.C(n_663),
.Y(n_1013)
);

AO22x2_ASAP7_75t_L g1014 ( 
.A1(n_915),
.A2(n_6),
.B1(n_2),
.B2(n_5),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_914),
.B(n_667),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_914),
.B(n_668),
.Y(n_1016)
);

OAI221xp5_ASAP7_75t_L g1017 ( 
.A1(n_912),
.A2(n_690),
.B1(n_692),
.B2(n_689),
.C(n_686),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_942),
.B(n_695),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_919),
.A2(n_673),
.B1(n_676),
.B2(n_671),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_944),
.Y(n_1020)
);

INVxp33_ASAP7_75t_SL g1021 ( 
.A(n_920),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_942),
.B(n_711),
.Y(n_1022)
);

NAND2x1p5_ASAP7_75t_L g1023 ( 
.A(n_918),
.B(n_630),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_960),
.B(n_716),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_SL g1025 ( 
.A(n_975),
.B(n_677),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_998),
.B(n_678),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_1008),
.B(n_679),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_1015),
.B(n_682),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_1016),
.B(n_981),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_961),
.B(n_683),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_946),
.B(n_684),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_956),
.B(n_688),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_949),
.B(n_950),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_1018),
.B(n_1022),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_951),
.B(n_696),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_984),
.B(n_700),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_988),
.B(n_703),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_995),
.B(n_705),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_996),
.B(n_707),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_999),
.B(n_708),
.Y(n_1040)
);

NAND2xp33_ASAP7_75t_SL g1041 ( 
.A(n_954),
.B(n_709),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_1001),
.B(n_710),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_1003),
.B(n_714),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_1004),
.B(n_715),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_991),
.B(n_720),
.Y(n_1045)
);

NAND2xp33_ASAP7_75t_SL g1046 ( 
.A(n_992),
.B(n_724),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_1007),
.B(n_725),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_1009),
.B(n_726),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_1011),
.B(n_727),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_1012),
.B(n_728),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_1020),
.B(n_729),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_953),
.B(n_734),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_955),
.B(n_962),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_SL g1054 ( 
.A(n_1005),
.B(n_738),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_973),
.B(n_742),
.Y(n_1055)
);

NAND2xp33_ASAP7_75t_SL g1056 ( 
.A(n_979),
.B(n_743),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_968),
.B(n_745),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_1006),
.B(n_751),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_1021),
.B(n_1019),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_972),
.B(n_294),
.Y(n_1060)
);

NAND2xp33_ASAP7_75t_SL g1061 ( 
.A(n_982),
.B(n_757),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_945),
.B(n_964),
.Y(n_1062)
);

NAND2xp33_ASAP7_75t_SL g1063 ( 
.A(n_1002),
.B(n_763),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_969),
.B(n_765),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_970),
.B(n_772),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_985),
.B(n_785),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_977),
.B(n_789),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_948),
.B(n_790),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_965),
.B(n_798),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_1023),
.B(n_803),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_963),
.B(n_1000),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_986),
.B(n_809),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_SL g1073 ( 
.A(n_990),
.B(n_810),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_993),
.B(n_813),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_959),
.B(n_818),
.Y(n_1075)
);

NAND2xp33_ASAP7_75t_SL g1076 ( 
.A(n_1010),
.B(n_821),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_SL g1077 ( 
.A(n_1014),
.B(n_828),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_976),
.B(n_833),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_947),
.B(n_835),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_958),
.B(n_733),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_958),
.B(n_837),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_957),
.B(n_295),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_974),
.B(n_845),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_980),
.B(n_847),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_952),
.B(n_776),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_983),
.B(n_853),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_997),
.B(n_687),
.Y(n_1087)
);

NAND2xp33_ASAP7_75t_SL g1088 ( 
.A(n_971),
.B(n_780),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_SL g1089 ( 
.A(n_967),
.B(n_783),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_1013),
.B(n_633),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_1017),
.B(n_633),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_989),
.B(n_644),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_994),
.B(n_644),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_978),
.B(n_657),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_966),
.B(n_657),
.Y(n_1095)
);

NAND2xp33_ASAP7_75t_SL g1096 ( 
.A(n_975),
.B(n_796),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_972),
.B(n_296),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_960),
.B(n_759),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_SL g1099 ( 
.A(n_975),
.B(n_797),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_960),
.B(n_759),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_960),
.B(n_767),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_960),
.B(n_767),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_960),
.B(n_804),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_960),
.B(n_770),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_960),
.B(n_770),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_987),
.B(n_687),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_960),
.B(n_770),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_960),
.B(n_806),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_972),
.B(n_298),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_987),
.B(n_687),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_960),
.B(n_788),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_960),
.B(n_788),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_SL g1113 ( 
.A(n_975),
.B(n_812),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_987),
.B(n_687),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_960),
.B(n_795),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_L g1116 ( 
.A(n_987),
.B(n_687),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_960),
.B(n_801),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_960),
.B(n_801),
.Y(n_1118)
);

NAND2xp33_ASAP7_75t_SL g1119 ( 
.A(n_975),
.B(n_814),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_987),
.B(n_807),
.Y(n_1120)
);

NAND2xp33_ASAP7_75t_SL g1121 ( 
.A(n_975),
.B(n_824),
.Y(n_1121)
);

NAND2xp33_ASAP7_75t_L g1122 ( 
.A(n_987),
.B(n_807),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_960),
.B(n_635),
.Y(n_1123)
);

NAND2xp33_ASAP7_75t_SL g1124 ( 
.A(n_975),
.B(n_836),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_SL g1125 ( 
.A(n_1006),
.B(n_756),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_960),
.B(n_635),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_960),
.B(n_782),
.Y(n_1127)
);

NAND2xp33_ASAP7_75t_R g1128 ( 
.A(n_954),
.B(n_846),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_960),
.B(n_782),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_987),
.B(n_807),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_960),
.B(n_782),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_987),
.B(n_807),
.Y(n_1132)
);

NAND2xp33_ASAP7_75t_SL g1133 ( 
.A(n_975),
.B(n_849),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_960),
.B(n_795),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_960),
.B(n_801),
.Y(n_1135)
);

NAND2xp33_ASAP7_75t_SL g1136 ( 
.A(n_975),
.B(n_6),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_960),
.B(n_807),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_960),
.B(n_299),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_960),
.B(n_300),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_960),
.B(n_301),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_960),
.B(n_302),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1033),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1024),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_1029),
.A2(n_306),
.B(n_307),
.C(n_303),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1106),
.A2(n_309),
.B(n_308),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1110),
.A2(n_311),
.B(n_310),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1114),
.A2(n_315),
.B(n_312),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1060),
.Y(n_1148)
);

OR2x6_ASAP7_75t_L g1149 ( 
.A(n_1071),
.B(n_7),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_1087),
.A2(n_625),
.A3(n_624),
.B(n_317),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1053),
.A2(n_318),
.B(n_316),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1062),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1026),
.A2(n_1028),
.B(n_1027),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1034),
.B(n_8),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_SL g1155 ( 
.A(n_1125),
.B(n_9),
.C(n_10),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1120),
.A2(n_320),
.B(n_319),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_SL g1157 ( 
.A1(n_1138),
.A2(n_322),
.B(n_323),
.C(n_321),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1130),
.A2(n_326),
.B(n_324),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_1103),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1031),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_1132),
.A2(n_622),
.A3(n_623),
.B(n_621),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1137),
.A2(n_330),
.B(n_328),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1108),
.B(n_11),
.Y(n_1163)
);

BUFx12f_ASAP7_75t_L g1164 ( 
.A(n_1082),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1045),
.B(n_12),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1060),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1059),
.B(n_13),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1035),
.A2(n_1037),
.B(n_1036),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1052),
.A2(n_333),
.B1(n_334),
.B2(n_331),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1097),
.A2(n_336),
.B(n_335),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1038),
.A2(n_338),
.B(n_337),
.Y(n_1171)
);

NAND2x1p5_ASAP7_75t_L g1172 ( 
.A(n_1097),
.B(n_339),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1039),
.A2(n_341),
.B(n_340),
.Y(n_1173)
);

BUFx12f_ASAP7_75t_L g1174 ( 
.A(n_1082),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1057),
.B(n_15),
.Y(n_1175)
);

OAI22x1_ASAP7_75t_L g1176 ( 
.A1(n_1075),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1065),
.A2(n_345),
.B(n_343),
.Y(n_1177)
);

AOI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1040),
.A2(n_347),
.B(n_346),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_1128),
.B(n_16),
.C(n_17),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1032),
.A2(n_349),
.B1(n_350),
.B2(n_348),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1109),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1116),
.A2(n_615),
.A3(n_616),
.B(n_614),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_1058),
.B(n_18),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1042),
.A2(n_353),
.B1(n_354),
.B2(n_351),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1043),
.A2(n_1047),
.B(n_1044),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1098),
.B(n_18),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1100),
.Y(n_1187)
);

BUFx10_ASAP7_75t_L g1188 ( 
.A(n_1041),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1048),
.A2(n_358),
.B(n_357),
.Y(n_1189)
);

OAI22x1_ASAP7_75t_L g1190 ( 
.A1(n_1079),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1101),
.B(n_21),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1049),
.A2(n_361),
.B(n_360),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1050),
.A2(n_365),
.B(n_363),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1102),
.B(n_22),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1051),
.A2(n_368),
.B(n_366),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1064),
.A2(n_373),
.B(n_372),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1104),
.B(n_23),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1080),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1122),
.A2(n_620),
.A3(n_375),
.B(n_376),
.Y(n_1199)
);

NAND3x1_ASAP7_75t_L g1200 ( 
.A(n_1085),
.B(n_25),
.C(n_26),
.Y(n_1200)
);

INVx4_ASAP7_75t_L g1201 ( 
.A(n_1046),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_SL g1202 ( 
.A(n_1054),
.B(n_374),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1055),
.A2(n_378),
.B1(n_380),
.B2(n_377),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1105),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1073),
.B(n_381),
.Y(n_1205)
);

AOI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1030),
.A2(n_384),
.B(n_382),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1139),
.A2(n_387),
.B(n_386),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1140),
.Y(n_1208)
);

AO32x2_ASAP7_75t_L g1209 ( 
.A1(n_1076),
.A2(n_1077),
.A3(n_1074),
.B1(n_1072),
.B2(n_1086),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1107),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1141),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1084),
.B(n_25),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1111),
.B(n_26),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1081),
.B(n_390),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_1136),
.Y(n_1215)
);

AO21x2_ASAP7_75t_L g1216 ( 
.A1(n_1067),
.A2(n_392),
.B(n_391),
.Y(n_1216)
);

INVxp67_ASAP7_75t_L g1217 ( 
.A(n_1056),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1112),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1115),
.B(n_27),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1117),
.Y(n_1220)
);

CKINVDCx8_ASAP7_75t_R g1221 ( 
.A(n_1096),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1090),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_1222)
);

BUFx12f_ASAP7_75t_L g1223 ( 
.A(n_1088),
.Y(n_1223)
);

OR2x6_ASAP7_75t_L g1224 ( 
.A(n_1078),
.B(n_28),
.Y(n_1224)
);

NAND3x1_ASAP7_75t_L g1225 ( 
.A(n_1099),
.B(n_31),
.C(n_32),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1118),
.B(n_32),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1123),
.A2(n_400),
.B(n_399),
.Y(n_1227)
);

AOI221x1_ASAP7_75t_L g1228 ( 
.A1(n_1089),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.C(n_36),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1126),
.A2(n_403),
.B(n_401),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1127),
.B(n_33),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1129),
.B(n_34),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1131),
.B(n_35),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1159),
.B(n_1134),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1143),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1145),
.A2(n_1066),
.B(n_1135),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1146),
.A2(n_1070),
.B(n_1068),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1142),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1152),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1147),
.A2(n_1158),
.B(n_1156),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1160),
.B(n_1091),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1181),
.A2(n_1069),
.B1(n_1093),
.B2(n_1092),
.Y(n_1241)
);

BUFx12f_ASAP7_75t_L g1242 ( 
.A(n_1164),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1174),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1153),
.A2(n_1061),
.B(n_1063),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1148),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_SL g1246 ( 
.A(n_1221),
.B(n_1025),
.Y(n_1246)
);

INVxp67_ASAP7_75t_L g1247 ( 
.A(n_1198),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1167),
.A2(n_1094),
.B1(n_1095),
.B2(n_1083),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1215),
.A2(n_1113),
.B1(n_1121),
.B2(n_1119),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1166),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1162),
.A2(n_1133),
.B(n_1124),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1154),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1189),
.A2(n_406),
.B(n_404),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1187),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1223),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1163),
.B(n_37),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1217),
.B(n_408),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1165),
.B(n_1208),
.Y(n_1258)
);

AOI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1168),
.A2(n_1185),
.B(n_1205),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1183),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1188),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1175),
.B(n_1211),
.Y(n_1262)
);

AOI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1206),
.A2(n_411),
.B(n_410),
.Y(n_1263)
);

AO21x1_ASAP7_75t_L g1264 ( 
.A1(n_1222),
.A2(n_40),
.B(n_39),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1192),
.A2(n_1195),
.B(n_1193),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1204),
.A2(n_1210),
.B1(n_1220),
.B2(n_1218),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_SL g1267 ( 
.A1(n_1178),
.A2(n_414),
.B(n_413),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1209),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1201),
.B(n_416),
.Y(n_1269)
);

OR2x6_ASAP7_75t_L g1270 ( 
.A(n_1172),
.B(n_417),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1207),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1219),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1149),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1212),
.B(n_44),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1227),
.A2(n_421),
.B(n_418),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1214),
.B(n_45),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1151),
.A2(n_423),
.B(n_422),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_SL g1278 ( 
.A1(n_1229),
.A2(n_428),
.B(n_426),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1213),
.B(n_46),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1224),
.A2(n_1155),
.B1(n_1190),
.B2(n_1176),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1224),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1186),
.B(n_46),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1191),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1194),
.A2(n_430),
.B(n_429),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1197),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1180),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1149),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1202),
.A2(n_433),
.B(n_432),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1226),
.A2(n_1232),
.B(n_1231),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1171),
.A2(n_435),
.B(n_434),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1230),
.B(n_47),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_1200),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1173),
.A2(n_438),
.B(n_436),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1196),
.A2(n_441),
.B(n_440),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1179),
.B(n_443),
.Y(n_1295)
);

INVx8_ASAP7_75t_L g1296 ( 
.A(n_1170),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1184),
.Y(n_1297)
);

AOI21xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1169),
.A2(n_50),
.B(n_51),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1228),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1216),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1182),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1150),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1203),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1177),
.A2(n_445),
.B(n_444),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1225),
.A2(n_447),
.B(n_446),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1150),
.A2(n_450),
.B(n_448),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1144),
.A2(n_452),
.B(n_451),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1157),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1182),
.B(n_453),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1199),
.B(n_454),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1161),
.Y(n_1311)
);

NAND2x1p5_ASAP7_75t_L g1312 ( 
.A(n_1159),
.B(n_468),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1145),
.A2(n_460),
.B(n_459),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1143),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1142),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1142),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1142),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1145),
.A2(n_465),
.B(n_461),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1228),
.A2(n_467),
.A3(n_469),
.B(n_466),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1145),
.A2(n_472),
.B(n_470),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1145),
.A2(n_477),
.B(n_473),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1164),
.Y(n_1322)
);

OR2x6_ASAP7_75t_L g1323 ( 
.A(n_1164),
.B(n_478),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1142),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1159),
.B(n_488),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1145),
.A2(n_482),
.B(n_480),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1164),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1153),
.A2(n_486),
.B(n_483),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1167),
.A2(n_55),
.B1(n_52),
.B2(n_54),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1237),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1315),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1316),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1317),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1324),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1243),
.B(n_487),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1238),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1322),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1254),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1266),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1265),
.A2(n_490),
.B(n_489),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1252),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1283),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1297),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1343)
);

AO31x2_ASAP7_75t_L g1344 ( 
.A1(n_1311),
.A2(n_493),
.A3(n_494),
.B(n_492),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1285),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1245),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1250),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1322),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1262),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1242),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1327),
.Y(n_1351)
);

AOI21xp33_ASAP7_75t_L g1352 ( 
.A1(n_1248),
.A2(n_56),
.B(n_58),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1314),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1260),
.B(n_59),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1327),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1240),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1291),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1268),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1239),
.A2(n_1236),
.B(n_1259),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1258),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1247),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1234),
.Y(n_1362)
);

OR2x6_ASAP7_75t_L g1363 ( 
.A(n_1270),
.B(n_498),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1302),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1271),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1244),
.A2(n_501),
.B(n_499),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1299),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1255),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1261),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1255),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1263),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1309),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1279),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1289),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1264),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1286),
.A2(n_60),
.B(n_61),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1267),
.Y(n_1377)
);

AOI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1301),
.A2(n_503),
.B(n_502),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1319),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1233),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1278),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1274),
.B(n_61),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1319),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1257),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1273),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1292),
.B(n_504),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1241),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1313),
.A2(n_507),
.B(n_506),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1310),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1290),
.Y(n_1390)
);

AOI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1235),
.A2(n_509),
.B(n_508),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1256),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1282),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1361),
.Y(n_1394)
);

XNOR2xp5_ASAP7_75t_L g1395 ( 
.A(n_1384),
.B(n_1287),
.Y(n_1395)
);

NAND2xp33_ASAP7_75t_SL g1396 ( 
.A(n_1393),
.B(n_1281),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1349),
.B(n_1280),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1392),
.B(n_1249),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1367),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1330),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1337),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1353),
.B(n_1270),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1337),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_R g1404 ( 
.A(n_1350),
.B(n_1246),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1360),
.B(n_1295),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1331),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1370),
.Y(n_1407)
);

NAND2xp33_ASAP7_75t_R g1408 ( 
.A(n_1363),
.B(n_1323),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_R g1409 ( 
.A(n_1355),
.B(n_1369),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1355),
.Y(n_1410)
);

NAND2xp33_ASAP7_75t_R g1411 ( 
.A(n_1363),
.B(n_1269),
.Y(n_1411)
);

INVxp67_ASAP7_75t_L g1412 ( 
.A(n_1380),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1362),
.Y(n_1413)
);

XNOR2xp5_ASAP7_75t_L g1414 ( 
.A(n_1385),
.B(n_1312),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1334),
.Y(n_1415)
);

OR2x6_ASAP7_75t_L g1416 ( 
.A(n_1389),
.B(n_1296),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1348),
.B(n_1281),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1351),
.B(n_1372),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1356),
.B(n_1276),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1373),
.B(n_1329),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1332),
.Y(n_1421)
);

NAND2xp33_ASAP7_75t_R g1422 ( 
.A(n_1335),
.B(n_1308),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1333),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1346),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1336),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1347),
.B(n_1305),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1382),
.B(n_1272),
.Y(n_1427)
);

CKINVDCx16_ASAP7_75t_R g1428 ( 
.A(n_1368),
.Y(n_1428)
);

NAND2xp33_ASAP7_75t_R g1429 ( 
.A(n_1386),
.B(n_1306),
.Y(n_1429)
);

BUFx10_ASAP7_75t_L g1430 ( 
.A(n_1357),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1338),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1341),
.B(n_1288),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1398),
.A2(n_1376),
.B1(n_1352),
.B2(n_1303),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1423),
.B(n_1387),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1431),
.B(n_1374),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1424),
.B(n_1358),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1415),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1412),
.B(n_1342),
.Y(n_1438)
);

INVxp67_ASAP7_75t_SL g1439 ( 
.A(n_1399),
.Y(n_1439)
);

AND2x4_ASAP7_75t_SL g1440 ( 
.A(n_1430),
.B(n_1345),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1400),
.B(n_1364),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1406),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1419),
.B(n_1354),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1421),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1425),
.B(n_1379),
.Y(n_1445)
);

NAND2x1_ASAP7_75t_L g1446 ( 
.A(n_1416),
.B(n_1339),
.Y(n_1446)
);

AOI21xp33_ASAP7_75t_L g1447 ( 
.A1(n_1429),
.A2(n_1375),
.B(n_1420),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1426),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1413),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1394),
.B(n_1343),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1397),
.B(n_1383),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1405),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1427),
.B(n_1377),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1416),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1402),
.B(n_1381),
.Y(n_1455)
);

AND2x4_ASAP7_75t_SL g1456 ( 
.A(n_1418),
.B(n_1365),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1432),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1414),
.B(n_1344),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1401),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1395),
.B(n_1344),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1403),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1409),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1396),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1428),
.B(n_1371),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1417),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1404),
.B(n_1325),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1407),
.B(n_1359),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1410),
.B(n_1298),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1422),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1408),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1411),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1433),
.A2(n_1277),
.B1(n_1284),
.B2(n_1366),
.Y(n_1472)
);

OAI31xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1447),
.A2(n_1251),
.A3(n_1340),
.B(n_1388),
.Y(n_1473)
);

INVx5_ASAP7_75t_L g1474 ( 
.A(n_1459),
.Y(n_1474)
);

INVxp67_ASAP7_75t_SL g1475 ( 
.A(n_1445),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1442),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1459),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_R g1478 ( 
.A(n_1469),
.B(n_62),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1444),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1441),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1470),
.B(n_1390),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1459),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1454),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1471),
.B(n_1328),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1437),
.Y(n_1485)
);

INVx5_ASAP7_75t_L g1486 ( 
.A(n_1462),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1440),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1436),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1461),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1460),
.B(n_1300),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1435),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1453),
.B(n_1391),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1457),
.B(n_1378),
.Y(n_1493)
);

INVx4_ASAP7_75t_L g1494 ( 
.A(n_1456),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1451),
.B(n_1391),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1434),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1449),
.B(n_1318),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1452),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1455),
.B(n_1320),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1448),
.B(n_1321),
.Y(n_1500)
);

NAND3xp33_ASAP7_75t_L g1501 ( 
.A(n_1443),
.B(n_1275),
.C(n_1378),
.Y(n_1501)
);

OAI33xp33_ASAP7_75t_L g1502 ( 
.A1(n_1438),
.A2(n_65),
.A3(n_67),
.B1(n_63),
.B2(n_64),
.B3(n_66),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1467),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1464),
.B(n_68),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1465),
.B(n_1463),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1466),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1458),
.B(n_1326),
.Y(n_1507)
);

INVx5_ASAP7_75t_L g1508 ( 
.A(n_1446),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1463),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1450),
.B(n_68),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1446),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1468),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1442),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1452),
.B(n_69),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1470),
.B(n_1304),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1470),
.B(n_1253),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1470),
.B(n_1293),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1439),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1439),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1433),
.A2(n_1294),
.B1(n_1307),
.B2(n_71),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1459),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1469),
.A2(n_511),
.B(n_510),
.Y(n_1522)
);

INVx4_ASAP7_75t_L g1523 ( 
.A(n_1459),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1452),
.B(n_69),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1469),
.B(n_70),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1442),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1439),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1449),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1442),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1488),
.B(n_71),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1483),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1476),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1474),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1503),
.B(n_72),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1479),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1486),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1486),
.B(n_73),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1513),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1486),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1475),
.B(n_74),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1505),
.B(n_74),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1526),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1529),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1496),
.B(n_75),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1518),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1480),
.B(n_1498),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1491),
.B(n_75),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1511),
.B(n_76),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1519),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1512),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1527),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1528),
.B(n_77),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1509),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1490),
.B(n_77),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1485),
.B(n_78),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1481),
.B(n_79),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1504),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1506),
.B(n_80),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1495),
.B(n_81),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1489),
.B(n_82),
.Y(n_1560)
);

NOR2x1_ASAP7_75t_L g1561 ( 
.A(n_1487),
.B(n_82),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1523),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1477),
.B(n_84),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1492),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1484),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1497),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1507),
.B(n_85),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_L g1568 ( 
.A(n_1472),
.B(n_85),
.C(n_86),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1493),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1515),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1500),
.Y(n_1571)
);

INVx6_ASAP7_75t_L g1572 ( 
.A(n_1474),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1508),
.B(n_88),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1517),
.B(n_88),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1482),
.B(n_1521),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1516),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1522),
.A2(n_513),
.B(n_512),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1508),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1510),
.B(n_89),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1514),
.B(n_89),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1494),
.B(n_1499),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1508),
.B(n_90),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1525),
.B(n_90),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1524),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1473),
.B(n_91),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1501),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1520),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1478),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1502),
.B(n_92),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_R g1590 ( 
.A(n_1487),
.B(n_93),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1483),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1488),
.B(n_94),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1483),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1498),
.B(n_94),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1483),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1498),
.B(n_95),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1498),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1498),
.B(n_95),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1476),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1503),
.B(n_96),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1498),
.B(n_97),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1503),
.B(n_97),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1476),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1483),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1557),
.B(n_98),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1587),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1606)
);

CKINVDCx8_ASAP7_75t_R g1607 ( 
.A(n_1573),
.Y(n_1607)
);

OAI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1585),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.C(n_104),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1586),
.B(n_103),
.Y(n_1609)
);

OAI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1536),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1553),
.B(n_105),
.Y(n_1611)
);

INVxp33_ASAP7_75t_SL g1612 ( 
.A(n_1590),
.Y(n_1612)
);

INVx3_ASAP7_75t_SL g1613 ( 
.A(n_1548),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1532),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1562),
.B(n_107),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1564),
.B(n_108),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1597),
.B(n_109),
.Y(n_1617)
);

AO221x2_ASAP7_75t_L g1618 ( 
.A1(n_1588),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.C(n_112),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1579),
.B(n_110),
.Y(n_1619)
);

INVxp33_ASAP7_75t_SL g1620 ( 
.A(n_1561),
.Y(n_1620)
);

NAND2xp33_ASAP7_75t_R g1621 ( 
.A(n_1573),
.B(n_111),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1545),
.B(n_112),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1549),
.B(n_113),
.Y(n_1623)
);

NAND2xp33_ASAP7_75t_SL g1624 ( 
.A(n_1537),
.B(n_113),
.Y(n_1624)
);

NOR2xp67_ASAP7_75t_L g1625 ( 
.A(n_1578),
.B(n_114),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1539),
.B(n_115),
.Y(n_1626)
);

OAI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1559),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_1627)
);

NOR2x1_ASAP7_75t_L g1628 ( 
.A(n_1582),
.B(n_116),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1572),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1569),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1551),
.B(n_1546),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1589),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1580),
.B(n_119),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1535),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1600),
.B(n_120),
.Y(n_1635)
);

NOR2xp67_ASAP7_75t_L g1636 ( 
.A(n_1533),
.B(n_121),
.Y(n_1636)
);

OAI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1577),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.C(n_125),
.Y(n_1637)
);

AO221x1_ASAP7_75t_L g1638 ( 
.A1(n_1570),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.C(n_126),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1576),
.B(n_127),
.Y(n_1639)
);

NAND2xp33_ASAP7_75t_SL g1640 ( 
.A(n_1602),
.B(n_128),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1565),
.B(n_129),
.Y(n_1641)
);

AO221x2_ASAP7_75t_L g1642 ( 
.A1(n_1531),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.C(n_133),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1567),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_1643)
);

NAND2xp33_ASAP7_75t_SL g1644 ( 
.A(n_1534),
.B(n_135),
.Y(n_1644)
);

OAI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1556),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.C(n_141),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1581),
.A2(n_1548),
.B1(n_1572),
.B2(n_1541),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1552),
.B(n_140),
.Y(n_1647)
);

AO221x2_ASAP7_75t_L g1648 ( 
.A1(n_1594),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.C(n_145),
.Y(n_1648)
);

AO221x2_ASAP7_75t_L g1649 ( 
.A1(n_1596),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.C(n_149),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1598),
.B(n_150),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1571),
.Y(n_1651)
);

AO221x2_ASAP7_75t_L g1652 ( 
.A1(n_1591),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.C(n_153),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1566),
.B(n_153),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1575),
.B(n_154),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1601),
.B(n_154),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1599),
.B(n_155),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1563),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1583),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1603),
.Y(n_1659)
);

AND2x4_ASAP7_75t_SL g1660 ( 
.A(n_1593),
.B(n_155),
.Y(n_1660)
);

AO221x2_ASAP7_75t_L g1661 ( 
.A1(n_1595),
.A2(n_159),
.B1(n_156),
.B2(n_158),
.C(n_160),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1604),
.B(n_156),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1538),
.B(n_158),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1554),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_1664)
);

AO221x2_ASAP7_75t_L g1665 ( 
.A1(n_1542),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.C(n_164),
.Y(n_1665)
);

NAND2xp33_ASAP7_75t_SL g1666 ( 
.A(n_1540),
.B(n_162),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1558),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_1667)
);

AO221x2_ASAP7_75t_L g1668 ( 
.A1(n_1543),
.A2(n_169),
.B1(n_166),
.B2(n_167),
.C(n_170),
.Y(n_1668)
);

AO221x2_ASAP7_75t_L g1669 ( 
.A1(n_1530),
.A2(n_170),
.B1(n_166),
.B2(n_169),
.C(n_171),
.Y(n_1669)
);

NAND2xp33_ASAP7_75t_SL g1670 ( 
.A(n_1592),
.B(n_171),
.Y(n_1670)
);

NOR2xp67_ASAP7_75t_L g1671 ( 
.A(n_1574),
.B(n_172),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_L g1672 ( 
.A(n_1560),
.B(n_173),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1555),
.B(n_174),
.Y(n_1673)
);

CKINVDCx20_ASAP7_75t_R g1674 ( 
.A(n_1544),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1547),
.B(n_174),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1575),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1557),
.B(n_175),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1536),
.B(n_175),
.Y(n_1678)
);

INVx4_ASAP7_75t_L g1679 ( 
.A(n_1573),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1597),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1590),
.Y(n_1681)
);

OAI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1585),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1550),
.B(n_177),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1568),
.A2(n_181),
.B(n_179),
.C(n_180),
.Y(n_1684)
);

OAI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1585),
.A2(n_182),
.B1(n_179),
.B2(n_181),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1532),
.Y(n_1686)
);

OAI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1585),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1584),
.B(n_183),
.Y(n_1688)
);

NAND2xp33_ASAP7_75t_SL g1689 ( 
.A(n_1590),
.B(n_186),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1584),
.B(n_186),
.Y(n_1690)
);

OAI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1585),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1584),
.B(n_187),
.Y(n_1692)
);

CKINVDCx14_ASAP7_75t_R g1693 ( 
.A(n_1590),
.Y(n_1693)
);

AO221x2_ASAP7_75t_L g1694 ( 
.A1(n_1588),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_191),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1620),
.B(n_191),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1680),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1609),
.B(n_192),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1679),
.B(n_1629),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1612),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1659),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1614),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1634),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1681),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1676),
.B(n_194),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1613),
.B(n_195),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1646),
.B(n_1651),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1663),
.B(n_195),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1686),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1656),
.B(n_196),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1616),
.B(n_196),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1662),
.B(n_198),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1654),
.B(n_198),
.Y(n_1712)
);

NOR2x1_ASAP7_75t_L g1713 ( 
.A(n_1678),
.B(n_199),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1621),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1628),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1641),
.B(n_199),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1636),
.B(n_200),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1639),
.B(n_200),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1617),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1607),
.B(n_1657),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1653),
.B(n_201),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1683),
.B(n_202),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1671),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1658),
.B(n_202),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1608),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1684),
.B(n_203),
.C(n_205),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1622),
.B(n_206),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1672),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1615),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1688),
.B(n_206),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1689),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1623),
.B(n_207),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1690),
.B(n_207),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1626),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1692),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1673),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1660),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1635),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1625),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1611),
.B(n_208),
.Y(n_1740)
);

CKINVDCx16_ASAP7_75t_R g1741 ( 
.A(n_1693),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1644),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1674),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1647),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1675),
.B(n_209),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1666),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1638),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1605),
.B(n_209),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1665),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1665),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1661),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1668),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1668),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1661),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1648),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1648),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1633),
.B(n_210),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1677),
.B(n_210),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1650),
.B(n_1655),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1619),
.B(n_211),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1632),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1682),
.B(n_211),
.Y(n_1762)
);

AOI22x1_ASAP7_75t_L g1763 ( 
.A1(n_1649),
.A2(n_215),
.B1(n_212),
.B2(n_213),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1669),
.B(n_212),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1649),
.Y(n_1765)
);

INVx1_ASAP7_75t_SL g1766 ( 
.A(n_1670),
.Y(n_1766)
);

BUFx3_ASAP7_75t_L g1767 ( 
.A(n_1618),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1640),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1669),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1685),
.B(n_215),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1687),
.B(n_216),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1694),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1694),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1642),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1624),
.Y(n_1775)
);

BUFx3_ASAP7_75t_L g1776 ( 
.A(n_1652),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1667),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1691),
.A2(n_216),
.B(n_217),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1645),
.A2(n_217),
.B(n_218),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1627),
.Y(n_1780)
);

INVx4_ASAP7_75t_L g1781 ( 
.A(n_1610),
.Y(n_1781)
);

AND2x4_ASAP7_75t_SL g1782 ( 
.A(n_1664),
.B(n_219),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1643),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1637),
.B(n_220),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1606),
.B(n_220),
.Y(n_1785)
);

INVx3_ASAP7_75t_SL g1786 ( 
.A(n_1681),
.Y(n_1786)
);

AND2x4_ASAP7_75t_SL g1787 ( 
.A(n_1679),
.B(n_221),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1608),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1620),
.B(n_223),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1680),
.B(n_225),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1679),
.B(n_225),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1620),
.B(n_227),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1680),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1607),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1630),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1612),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1631),
.B(n_227),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1629),
.B(n_228),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1614),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1629),
.B(n_228),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1680),
.B(n_229),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1620),
.B(n_229),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1631),
.B(n_230),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1614),
.Y(n_1804)
);

AND3x1_ASAP7_75t_L g1805 ( 
.A(n_1678),
.B(n_231),
.C(n_232),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1629),
.B(n_232),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1629),
.B(n_233),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1630),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1614),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_SL g1810 ( 
.A(n_1620),
.B(n_234),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1608),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_1811)
);

INVxp67_ASAP7_75t_L g1812 ( 
.A(n_1678),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_SL g1813 ( 
.A(n_1620),
.B(n_235),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1614),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1614),
.Y(n_1815)
);

BUFx3_ASAP7_75t_L g1816 ( 
.A(n_1681),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1680),
.B(n_237),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1614),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1680),
.B(n_237),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1608),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1629),
.B(n_238),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1629),
.B(n_239),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1629),
.B(n_240),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1629),
.B(n_241),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1680),
.Y(n_1825)
);

NAND2x1p5_ASAP7_75t_L g1826 ( 
.A(n_1679),
.B(n_241),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1631),
.B(n_242),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1680),
.B(n_242),
.Y(n_1828)
);

INVx2_ASAP7_75t_SL g1829 ( 
.A(n_1613),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1701),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1741),
.B(n_243),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1708),
.Y(n_1832)
);

OAI33xp33_ASAP7_75t_L g1833 ( 
.A1(n_1765),
.A2(n_246),
.A3(n_248),
.B1(n_244),
.B2(n_245),
.B3(n_247),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1702),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1715),
.B(n_244),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1699),
.B(n_1796),
.Y(n_1836)
);

O2A1O1Ixp5_ASAP7_75t_L g1837 ( 
.A1(n_1781),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1772),
.A2(n_1755),
.B1(n_1751),
.B2(n_1769),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1774),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1754),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1749),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1799),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1804),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1786),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1809),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1738),
.B(n_252),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1714),
.B(n_253),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1814),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1779),
.A2(n_254),
.B(n_255),
.Y(n_1849)
);

INVx2_ASAP7_75t_SL g1850 ( 
.A(n_1816),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1696),
.B(n_255),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1728),
.B(n_256),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1731),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1794),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1747),
.B(n_256),
.Y(n_1855)
);

INVx1_ASAP7_75t_SL g1856 ( 
.A(n_1743),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1829),
.B(n_1746),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1815),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1723),
.B(n_257),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1698),
.B(n_258),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1818),
.Y(n_1861)
);

OAI21xp33_ASAP7_75t_L g1862 ( 
.A1(n_1725),
.A2(n_258),
.B(n_259),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1750),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_1863)
);

INVx2_ASAP7_75t_SL g1864 ( 
.A(n_1734),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1812),
.B(n_1752),
.Y(n_1865)
);

INVx2_ASAP7_75t_SL g1866 ( 
.A(n_1739),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_SL g1867 ( 
.A1(n_1805),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1720),
.Y(n_1868)
);

NAND4xp25_ASAP7_75t_L g1869 ( 
.A(n_1767),
.B(n_264),
.C(n_262),
.D(n_263),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1736),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1793),
.B(n_264),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_SL g1872 ( 
.A(n_1768),
.B(n_265),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1825),
.Y(n_1873)
);

OAI31xp33_ASAP7_75t_L g1874 ( 
.A1(n_1775),
.A2(n_1776),
.A3(n_1742),
.B(n_1766),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1706),
.B(n_266),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1700),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1719),
.Y(n_1877)
);

AOI211xp5_ASAP7_75t_L g1878 ( 
.A1(n_1771),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1735),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1753),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.C(n_273),
.Y(n_1880)
);

NOR2x1p5_ASAP7_75t_L g1881 ( 
.A(n_1756),
.B(n_273),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1703),
.Y(n_1882)
);

NOR2xp67_ASAP7_75t_L g1883 ( 
.A(n_1717),
.B(n_274),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1729),
.B(n_276),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1761),
.B(n_277),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1795),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1808),
.Y(n_1887)
);

OAI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1773),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1737),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1744),
.B(n_278),
.Y(n_1890)
);

INVxp67_ASAP7_75t_L g1891 ( 
.A(n_1713),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1777),
.B(n_279),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1791),
.Y(n_1893)
);

AO21x1_ASAP7_75t_L g1894 ( 
.A1(n_1810),
.A2(n_281),
.B(n_282),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1763),
.A2(n_1811),
.B1(n_1820),
.B2(n_1788),
.Y(n_1895)
);

AOI21xp33_ASAP7_75t_L g1896 ( 
.A1(n_1784),
.A2(n_281),
.B(n_282),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1780),
.Y(n_1897)
);

AOI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1726),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1783),
.A2(n_287),
.B1(n_284),
.B2(n_286),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1762),
.A2(n_1770),
.B(n_1792),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1705),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1695),
.Y(n_1902)
);

OAI21xp33_ASAP7_75t_L g1903 ( 
.A1(n_1778),
.A2(n_287),
.B(n_288),
.Y(n_1903)
);

AOI221x1_ASAP7_75t_L g1904 ( 
.A1(n_1764),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.C(n_291),
.Y(n_1904)
);

NAND4xp25_ASAP7_75t_SL g1905 ( 
.A(n_1785),
.B(n_292),
.C(n_290),
.D(n_291),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1717),
.B(n_293),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1790),
.Y(n_1907)
);

OAI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1789),
.A2(n_1802),
.B1(n_1813),
.B2(n_1759),
.C(n_1826),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1797),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1828),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1801),
.Y(n_1911)
);

O2A1O1Ixp33_ASAP7_75t_L g1912 ( 
.A1(n_1817),
.A2(n_1819),
.B(n_1748),
.C(n_1697),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1803),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1827),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1722),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1787),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1798),
.Y(n_1917)
);

XOR2xp5_ASAP7_75t_L g1918 ( 
.A(n_1745),
.B(n_517),
.Y(n_1918)
);

BUFx3_ASAP7_75t_L g1919 ( 
.A(n_1740),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1800),
.B(n_1806),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1710),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1704),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1807),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1900),
.A2(n_1709),
.B(n_1730),
.Y(n_1924)
);

INVx2_ASAP7_75t_SL g1925 ( 
.A(n_1919),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1891),
.B(n_1732),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1854),
.B(n_1821),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1838),
.B(n_1822),
.Y(n_1928)
);

INVxp67_ASAP7_75t_L g1929 ( 
.A(n_1836),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1866),
.B(n_1853),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1917),
.B(n_1823),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1889),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1857),
.B(n_1824),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1844),
.B(n_1716),
.Y(n_1934)
);

HB1xp67_ASAP7_75t_L g1935 ( 
.A(n_1864),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1901),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1915),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1850),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1882),
.B(n_1718),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1923),
.B(n_1727),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1856),
.B(n_1721),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1921),
.Y(n_1942)
);

INVx1_ASAP7_75t_SL g1943 ( 
.A(n_1916),
.Y(n_1943)
);

NAND2xp33_ASAP7_75t_SL g1944 ( 
.A(n_1867),
.B(n_1724),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1868),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1875),
.B(n_1757),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1922),
.B(n_1760),
.Y(n_1947)
);

OAI21xp5_ASAP7_75t_SL g1948 ( 
.A1(n_1874),
.A2(n_1782),
.B(n_1758),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1873),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1834),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1913),
.B(n_1712),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1902),
.B(n_1707),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1894),
.B(n_1712),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1914),
.B(n_1711),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1842),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1906),
.Y(n_1956)
);

AOI22xp33_ASAP7_75t_L g1957 ( 
.A1(n_1895),
.A2(n_1745),
.B1(n_1740),
.B2(n_1733),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1843),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1865),
.B(n_521),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1909),
.B(n_522),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1845),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1920),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1893),
.B(n_1897),
.Y(n_1963)
);

NOR2x1_ASAP7_75t_L g1964 ( 
.A(n_1872),
.B(n_523),
.Y(n_1964)
);

INVx2_ASAP7_75t_SL g1965 ( 
.A(n_1881),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1908),
.B(n_524),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1886),
.Y(n_1967)
);

AND2x4_ASAP7_75t_L g1968 ( 
.A(n_1883),
.B(n_525),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1885),
.B(n_526),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1830),
.B(n_527),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1884),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1887),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1848),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1859),
.B(n_528),
.Y(n_1974)
);

INVxp67_ASAP7_75t_L g1975 ( 
.A(n_1831),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1858),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1899),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1907),
.B(n_1910),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1911),
.B(n_532),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1862),
.A2(n_535),
.B1(n_533),
.B2(n_534),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1861),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1927),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1936),
.Y(n_1983)
);

BUFx2_ASAP7_75t_L g1984 ( 
.A(n_1965),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1954),
.Y(n_1985)
);

INVxp67_ASAP7_75t_SL g1986 ( 
.A(n_1953),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1944),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1978),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1949),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1950),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1955),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1958),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1961),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1973),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1976),
.Y(n_1995)
);

BUFx4f_ASAP7_75t_SL g1996 ( 
.A(n_1943),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1925),
.Y(n_1997)
);

CKINVDCx20_ASAP7_75t_R g1998 ( 
.A(n_1975),
.Y(n_1998)
);

INVx5_ASAP7_75t_L g1999 ( 
.A(n_1968),
.Y(n_1999)
);

INVx5_ASAP7_75t_L g2000 ( 
.A(n_1970),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1981),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1963),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1935),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1929),
.B(n_1956),
.Y(n_2004)
);

INVx1_ASAP7_75t_SL g2005 ( 
.A(n_1933),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1930),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1937),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1942),
.Y(n_2008)
);

BUFx2_ASAP7_75t_L g2009 ( 
.A(n_1938),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1951),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1932),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1947),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1948),
.B(n_1946),
.Y(n_2013)
);

NOR3xp33_ASAP7_75t_L g2014 ( 
.A(n_1987),
.B(n_1926),
.C(n_1934),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1996),
.B(n_1977),
.Y(n_2015)
);

INVxp67_ASAP7_75t_SL g2016 ( 
.A(n_1984),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1986),
.B(n_2005),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1983),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_2003),
.B(n_1931),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1985),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_SL g2021 ( 
.A(n_1998),
.B(n_1964),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_2000),
.B(n_1939),
.Y(n_2022)
);

NAND4xp25_ASAP7_75t_L g2023 ( 
.A(n_2013),
.B(n_1962),
.C(n_1957),
.D(n_1928),
.Y(n_2023)
);

OAI221xp5_ASAP7_75t_L g2024 ( 
.A1(n_2004),
.A2(n_1839),
.B1(n_1878),
.B2(n_1837),
.C(n_1849),
.Y(n_2024)
);

NOR4xp25_ASAP7_75t_SL g2025 ( 
.A(n_2009),
.B(n_1835),
.C(n_1860),
.D(n_1832),
.Y(n_2025)
);

NAND3xp33_ASAP7_75t_L g2026 ( 
.A(n_2006),
.B(n_1904),
.C(n_1880),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1997),
.B(n_1971),
.Y(n_2027)
);

NOR3xp33_ASAP7_75t_L g2028 ( 
.A(n_2002),
.B(n_1896),
.C(n_1945),
.Y(n_2028)
);

NOR3x1_ASAP7_75t_SL g2029 ( 
.A(n_1999),
.B(n_1905),
.C(n_1966),
.Y(n_2029)
);

NOR2xp67_ASAP7_75t_L g2030 ( 
.A(n_2000),
.B(n_1941),
.Y(n_2030)
);

OAI211xp5_ASAP7_75t_SL g2031 ( 
.A1(n_2012),
.A2(n_1924),
.B(n_1912),
.C(n_1940),
.Y(n_2031)
);

A2O1A1Ixp33_ASAP7_75t_L g2032 ( 
.A1(n_2026),
.A2(n_1903),
.B(n_1869),
.C(n_1898),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2016),
.Y(n_2033)
);

AOI221xp5_ASAP7_75t_L g2034 ( 
.A1(n_2023),
.A2(n_1988),
.B1(n_2010),
.B2(n_1989),
.C(n_2008),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_2015),
.Y(n_2035)
);

AOI211xp5_ASAP7_75t_L g2036 ( 
.A1(n_2031),
.A2(n_1888),
.B(n_1840),
.C(n_1863),
.Y(n_2036)
);

CKINVDCx16_ASAP7_75t_R g2037 ( 
.A(n_2021),
.Y(n_2037)
);

OAI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_2024),
.A2(n_1982),
.B1(n_1870),
.B2(n_2011),
.C(n_1999),
.Y(n_2038)
);

AND4x1_ASAP7_75t_L g2039 ( 
.A(n_2014),
.B(n_1952),
.C(n_1847),
.D(n_1855),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_2019),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2033),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2040),
.Y(n_2042)
);

NAND3x1_ASAP7_75t_L g2043 ( 
.A(n_2039),
.B(n_2017),
.C(n_2027),
.Y(n_2043)
);

AOI22xp33_ASAP7_75t_SL g2044 ( 
.A1(n_2037),
.A2(n_2029),
.B1(n_2025),
.B2(n_2018),
.Y(n_2044)
);

XNOR2x1_ASAP7_75t_L g2045 ( 
.A(n_2035),
.B(n_2030),
.Y(n_2045)
);

NAND4xp75_ASAP7_75t_L g2046 ( 
.A(n_2034),
.B(n_2022),
.C(n_2020),
.D(n_2007),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2032),
.B(n_2028),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2038),
.Y(n_2048)
);

NAND2xp33_ASAP7_75t_SL g2049 ( 
.A(n_2045),
.B(n_1851),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_R g2050 ( 
.A(n_2042),
.B(n_1846),
.Y(n_2050)
);

XNOR2xp5_ASAP7_75t_L g2051 ( 
.A(n_2043),
.B(n_2036),
.Y(n_2051)
);

XOR2xp5_ASAP7_75t_L g2052 ( 
.A(n_2044),
.B(n_1918),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_R g2053 ( 
.A(n_2048),
.B(n_1852),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2051),
.Y(n_2054)
);

AOI221xp5_ASAP7_75t_SL g2055 ( 
.A1(n_2052),
.A2(n_2047),
.B1(n_2041),
.B2(n_1991),
.C(n_1993),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2054),
.Y(n_2056)
);

O2A1O1Ixp33_ASAP7_75t_SL g2057 ( 
.A1(n_2056),
.A2(n_1992),
.B(n_1994),
.C(n_1990),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_2057),
.A2(n_2049),
.B1(n_2053),
.B2(n_2050),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_2057),
.A2(n_2001),
.B1(n_1995),
.B2(n_1967),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2058),
.B(n_2046),
.Y(n_2060)
);

OAI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_2059),
.A2(n_1972),
.B1(n_1877),
.B2(n_1879),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_2060),
.A2(n_1833),
.B1(n_1841),
.B2(n_1876),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_2061),
.A2(n_2055),
.B1(n_1892),
.B2(n_1974),
.Y(n_2063)
);

XNOR2xp5_ASAP7_75t_L g2064 ( 
.A(n_2063),
.B(n_1890),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2062),
.Y(n_2065)
);

OAI221xp5_ASAP7_75t_R g2066 ( 
.A1(n_2064),
.A2(n_1980),
.B1(n_1960),
.B2(n_1959),
.C(n_1871),
.Y(n_2066)
);

AOI211xp5_ASAP7_75t_L g2067 ( 
.A1(n_2066),
.A2(n_2065),
.B(n_1969),
.C(n_1979),
.Y(n_2067)
);


endmodule