module real_jpeg_23955_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_53),
.B1(n_54),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_1),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_1),
.A2(n_32),
.B1(n_40),
.B2(n_71),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_71),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_5),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_5),
.A2(n_67),
.B1(n_68),
.B2(n_146),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_146),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_146),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_6),
.A2(n_43),
.B1(n_149),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_6),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_154),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_154),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_6),
.A2(n_67),
.B1(n_68),
.B2(n_154),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_8),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_8),
.B(n_105),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_8),
.B(n_63),
.C(n_67),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_150),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_8),
.B(n_59),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_8),
.A2(n_90),
.B1(n_92),
.B2(n_221),
.Y(n_220)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_10),
.A2(n_37),
.B1(n_67),
.B2(n_68),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_11),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_48),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_11),
.A2(n_48),
.B1(n_67),
.B2(n_68),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_13),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_144),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_144),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_13),
.A2(n_67),
.B1(n_68),
.B2(n_144),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_14),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_14),
.A2(n_34),
.B1(n_53),
.B2(n_54),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_14),
.A2(n_34),
.B1(n_67),
.B2(n_68),
.Y(n_166)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_15),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_122),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_19),
.B(n_106),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.C(n_86),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_20),
.A2(n_74),
.B1(n_75),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_20),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_44),
.B2(n_73),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_21),
.A2(n_22),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_22),
.B(n_45),
.C(n_72),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B(n_35),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_23),
.A2(n_101),
.B1(n_153),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_24),
.A2(n_27),
.B(n_151),
.C(n_168),
.Y(n_167)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_25),
.B(n_26),
.C(n_38),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_26),
.A2(n_27),
.B1(n_52),
.B2(n_55),
.Y(n_56)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

HAxp5_ASAP7_75t_SL g239 ( 
.A(n_27),
.B(n_150),
.CON(n_239),
.SN(n_239)
);

NAND3xp33_ASAP7_75t_L g240 ( 
.A(n_27),
.B(n_53),
.C(n_55),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_29),
.Y(n_117)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_30),
.Y(n_149)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_41),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_36),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_38),
.B(n_150),
.Y(n_151)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_41),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_41),
.A2(n_105),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_41),
.A2(n_105),
.B1(n_148),
.B2(n_152),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_41),
.A2(n_105),
.B1(n_160),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_60),
.B2(n_72),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B(n_57),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_49),
.A2(n_113),
.B(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_49),
.A2(n_51),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_49),
.A2(n_57),
.B(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_59),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_58),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_50),
.A2(n_59),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_50),
.A2(n_59),
.B1(n_178),
.B2(n_239),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_51),
.A2(n_78),
.B(n_115),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_52),
.A2(n_54),
.B(n_239),
.C(n_240),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_54),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_59),
.B(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_60),
.A2(n_72),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B(n_69),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_61),
.A2(n_69),
.B(n_98),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_61),
.A2(n_66),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_61),
.A2(n_66),
.B1(n_198),
.B2(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_61),
.A2(n_81),
.B(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_61),
.A2(n_66),
.B1(n_97),
.B2(n_137),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_66),
.A2(n_83),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_66),
.B(n_150),
.Y(n_228)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_68),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_75),
.A2(n_76),
.B(n_80),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_84),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_82),
.A2(n_85),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_86),
.B(n_327),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_99),
.B(n_100),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_87),
.A2(n_88),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_89),
.A2(n_96),
.B1(n_99),
.B2(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_89),
.A2(n_99),
.B1(n_100),
.B2(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B(n_94),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_90),
.A2(n_92),
.B1(n_132),
.B2(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_90),
.B(n_135),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_90),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_90),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_90),
.A2(n_214),
.B1(n_221),
.B2(n_230),
.Y(n_229)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g184 ( 
.A(n_91),
.Y(n_184)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_91),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_93),
.B(n_95),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_95),
.A2(n_134),
.B(n_212),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_96),
.Y(n_299)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_100),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B(n_104),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_101),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_103),
.B(n_105),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_119),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_116),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_114),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_324),
.B(n_329),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_311),
.B(n_323),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_294),
.B(n_310),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_186),
.B(n_271),
.C(n_293),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_170),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_127),
.B(n_170),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_155),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_138),
.B2(n_139),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_129),
.B(n_139),
.C(n_155),
.Y(n_272)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_136),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_131),
.B(n_136),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_147),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_143),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_172),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B(n_151),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_150),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_163),
.B2(n_169),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_158),
.B(n_161),
.C(n_169),
.Y(n_292)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_163),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_167),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_166),
.A2(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.C(n_175),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_171),
.B(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_174),
.B(n_175),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.C(n_182),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_176),
.B(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_256)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_185),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_270),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_265),
.B(n_269),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_251),
.B(n_264),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_235),
.B(n_250),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_209),
.B(n_234),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_199),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_193),
.A2(n_195),
.B1(n_196),
.B2(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_206),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_204),
.C(n_206),
.Y(n_249)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_207),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_208),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_218),
.B(n_233),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_216),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_227),
.B(n_232),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_228),
.B(n_229),
.Y(n_232)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_249),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_249),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_244),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_245),
.C(n_248),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_238),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_243),
.Y(n_259)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_247),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_253),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_260),
.C(n_262),
.Y(n_268)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_259),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_268),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_273),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_292),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_284),
.B1(n_290),
.B2(n_291),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_280),
.Y(n_304)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_290),
.C(n_292),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_295),
.B(n_296),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_309),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_300),
.C(n_309),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_307),
.B2(n_308),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_306),
.C(n_308),
.Y(n_322)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_313),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_322),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_320),
.B2(n_321),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_320),
.C(n_322),
.Y(n_325)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);


endmodule