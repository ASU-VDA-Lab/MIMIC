module fake_jpeg_15896_n_265 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_14),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_0),
.A2(n_11),
.B(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_42),
.B(n_45),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_0),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_19),
.B(n_1),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_67),
.B(n_22),
.C(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_30),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_53),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_19),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_93)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_55),
.Y(n_81)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_59),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_4),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_5),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_5),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_27),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_27),
.Y(n_68)
);

AO21x1_ASAP7_75t_L g142 ( 
.A1(n_68),
.A2(n_74),
.B(n_77),
.Y(n_142)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_66),
.C(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_105),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_19),
.B1(n_36),
.B2(n_32),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_76),
.A2(n_88),
.B1(n_64),
.B2(n_14),
.Y(n_122)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_40),
.A2(n_36),
.B1(n_39),
.B2(n_37),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_80),
.A2(n_86),
.B(n_72),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_87),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_40),
.A2(n_26),
.B1(n_37),
.B2(n_35),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_38),
.B1(n_30),
.B2(n_22),
.Y(n_88)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_104),
.B1(n_69),
.B2(n_70),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_34),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_6),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_67),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_56),
.A2(n_30),
.B1(n_10),
.B2(n_12),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_8),
.B1(n_10),
.B2(n_14),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_115),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_8),
.B(n_10),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_112),
.B(n_118),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_63),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_15),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_119),
.A2(n_120),
.B1(n_127),
.B2(n_128),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_69),
.A2(n_55),
.B1(n_63),
.B2(n_62),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_43),
.C(n_41),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_125),
.C(n_141),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_123),
.B1(n_136),
.B2(n_141),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_78),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_131),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_73),
.C(n_68),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_135),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_79),
.A2(n_104),
.B1(n_99),
.B2(n_89),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_82),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_87),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_133),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_85),
.Y(n_135)
);

AO22x2_ASAP7_75t_L g136 ( 
.A1(n_85),
.A2(n_72),
.B1(n_90),
.B2(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_111),
.Y(n_148)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_75),
.B(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_138),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_102),
.B(n_76),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_164),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_130),
.B1(n_123),
.B2(n_128),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_160),
.B1(n_113),
.B2(n_129),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_122),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_159),
.C(n_166),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_136),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_174),
.B(n_129),
.Y(n_183)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_110),
.B(n_107),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_113),
.B(n_117),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_146),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_161),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_125),
.B(n_141),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_112),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_177),
.C(n_185),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_119),
.Y(n_177)
);

NAND2x1_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_134),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_183),
.B(n_187),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_193),
.B1(n_169),
.B2(n_165),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_174),
.B(n_163),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_188),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_147),
.C(n_148),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_191),
.C(n_198),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_166),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_147),
.A2(n_171),
.B1(n_150),
.B2(n_160),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_194),
.A2(n_199),
.B1(n_157),
.B2(n_170),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_158),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_153),
.C(n_149),
.Y(n_198)
);

AO22x1_ASAP7_75t_SL g199 ( 
.A1(n_161),
.A2(n_153),
.B1(n_163),
.B2(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_201),
.B(n_212),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_205),
.A2(n_211),
.B1(n_220),
.B2(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_156),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_180),
.A2(n_168),
.B(n_156),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_197),
.B(n_212),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_189),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_210),
.B(n_214),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_179),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_144),
.B1(n_193),
.B2(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_144),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_182),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_176),
.B(n_177),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_218),
.B(n_220),
.Y(n_225)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_175),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_190),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_224),
.C(n_228),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_185),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_198),
.C(n_192),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_229),
.A2(n_225),
.B(n_233),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_215),
.C(n_206),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_222),
.C(n_228),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_231),
.B(n_202),
.Y(n_237)
);

OAI22x1_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_205),
.B1(n_216),
.B2(n_201),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_225),
.B1(n_233),
.B2(n_227),
.Y(n_245)
);

AOI321xp33_ASAP7_75t_L g236 ( 
.A1(n_235),
.A2(n_214),
.A3(n_211),
.B1(n_216),
.B2(n_207),
.C(n_213),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_246),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_238),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_213),
.CI(n_204),
.CON(n_238),
.SN(n_238)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_218),
.B(n_200),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_229),
.A2(n_208),
.B(n_209),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_231),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_232),
.B1(n_226),
.B2(n_223),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_224),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_252),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_253),
.A2(n_244),
.B(n_241),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_240),
.B(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_247),
.C(n_249),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_257),
.Y(n_258)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_246),
.C(n_239),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_250),
.B(n_236),
.C(n_249),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_260),
.A2(n_256),
.B(n_242),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_251),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_258),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_264),
.Y(n_265)
);


endmodule