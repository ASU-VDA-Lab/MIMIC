module fake_jpeg_3583_n_395 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_4),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_56),
.Y(n_169)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g121 ( 
.A(n_57),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_8),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_58),
.B(n_100),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_8),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_98),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_28),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_68),
.A2(n_38),
.B(n_0),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

CKINVDCx6p67_ASAP7_75t_R g129 ( 
.A(n_69),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_70),
.Y(n_175)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_23),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_88),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_77),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_91),
.C(n_96),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_86),
.B(n_93),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

NAND2x1_ASAP7_75t_SL g91 ( 
.A(n_22),
.B(n_0),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_30),
.Y(n_92)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_94),
.B(n_95),
.Y(n_163)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_29),
.B(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_104),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_101),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_18),
.B(n_2),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_18),
.B(n_7),
.Y(n_102)
);

HAxp5_ASAP7_75t_SL g171 ( 
.A(n_102),
.B(n_100),
.CON(n_171),
.SN(n_171)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_20),
.B(n_9),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_19),
.C(n_49),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_105),
.B(n_106),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_107),
.B(n_98),
.Y(n_166)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_109),
.Y(n_118)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_32),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_51),
.B1(n_37),
.B2(n_53),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_112),
.A2(n_123),
.B1(n_126),
.B2(n_153),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_58),
.B(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_114),
.B(n_141),
.Y(n_208)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_32),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_115),
.B(n_171),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_116),
.B(n_159),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_119),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_65),
.A2(n_51),
.B1(n_53),
.B2(n_39),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_59),
.A2(n_27),
.B1(n_47),
.B2(n_46),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_124),
.A2(n_156),
.B1(n_164),
.B2(n_153),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_63),
.A2(n_39),
.B1(n_34),
.B2(n_25),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_34),
.C(n_25),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_138),
.B(n_121),
.C(n_129),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_73),
.A2(n_26),
.B1(n_47),
.B2(n_46),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_140),
.A2(n_162),
.B1(n_174),
.B2(n_129),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_21),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_92),
.B(n_21),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_157),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_67),
.A2(n_26),
.B1(n_38),
.B2(n_49),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_70),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_86),
.B(n_13),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_93),
.A2(n_94),
.B1(n_90),
.B2(n_78),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_104),
.A2(n_107),
.B1(n_106),
.B2(n_105),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_74),
.A2(n_87),
.B1(n_89),
.B2(n_79),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_163),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_101),
.B(n_57),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_68),
.B(n_69),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_62),
.B(n_58),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_140),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_73),
.A2(n_43),
.B1(n_104),
.B2(n_92),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_176),
.Y(n_251)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_177),
.Y(n_268)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_135),
.B(n_127),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_181),
.B(n_184),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_183),
.A2(n_190),
.B1(n_215),
.B2(n_208),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_117),
.B(n_115),
.Y(n_184)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_113),
.B(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_187),
.B(n_194),
.Y(n_243)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_188),
.Y(n_237)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_192),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_132),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_196),
.Y(n_258)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_197),
.Y(n_267)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_206),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_121),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_199),
.B(n_217),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_204),
.Y(n_246)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_120),
.B(n_155),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_202),
.B(n_205),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_203),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_129),
.B(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_207),
.B(n_226),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_124),
.B(n_145),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_209),
.B(n_211),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_213),
.B1(n_224),
.B2(n_216),
.Y(n_240)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_212),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_143),
.A2(n_163),
.B1(n_162),
.B2(n_165),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_147),
.B(n_122),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_219),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_147),
.B(n_170),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_225),
.Y(n_250)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_111),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_216),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_150),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_137),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_221),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_160),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_222),
.B(n_223),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_175),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_156),
.A2(n_123),
.B(n_112),
.C(n_174),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_210),
.Y(n_241)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_136),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_228),
.Y(n_264)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_229),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_142),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_238),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_164),
.B1(n_142),
.B2(n_158),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_231),
.A2(n_254),
.B1(n_267),
.B2(n_258),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_218),
.A2(n_158),
.B1(n_195),
.B2(n_213),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_235),
.A2(n_241),
.B1(n_253),
.B2(n_265),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_182),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_240),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_185),
.B(n_204),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_260),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_180),
.B(n_183),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_190),
.A2(n_196),
.B1(n_197),
.B2(n_191),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_178),
.B(n_177),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_270),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_188),
.B(n_186),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_192),
.B1(n_207),
.B2(n_229),
.Y(n_271)
);

INVxp33_ASAP7_75t_SL g303 ( 
.A(n_271),
.Y(n_303)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_260),
.A2(n_212),
.B1(n_221),
.B2(n_189),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_277),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_251),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_276),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_203),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_275),
.B(n_279),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_255),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_253),
.A2(n_227),
.B1(n_238),
.B2(n_246),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_255),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_268),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_280),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_236),
.B(n_252),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_291),
.B(n_299),
.Y(n_313)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_245),
.B(n_230),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_286),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_246),
.A2(n_240),
.B1(n_241),
.B2(n_235),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_287),
.B(n_264),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_234),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_289),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_246),
.B(n_242),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_264),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_233),
.B(n_263),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_250),
.Y(n_293)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_265),
.A2(n_247),
.B1(n_250),
.B2(n_269),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_294),
.A2(n_262),
.B1(n_264),
.B2(n_267),
.Y(n_319)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_295),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_248),
.A2(n_249),
.B(n_233),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_296),
.A2(n_297),
.B(n_232),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_259),
.A2(n_262),
.B(n_237),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_244),
.Y(n_298)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_239),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_237),
.B1(n_257),
.B2(n_239),
.Y(n_304)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_304),
.A2(n_322),
.B1(n_294),
.B2(n_297),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_272),
.B(n_283),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_307),
.B(n_310),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_284),
.A2(n_262),
.B(n_257),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_314),
.A2(n_275),
.B(n_291),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_295),
.Y(n_316)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_319),
.A2(n_301),
.B1(n_298),
.B2(n_299),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_323),
.B(n_278),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_322),
.A2(n_284),
.B1(n_281),
.B2(n_288),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_324),
.A2(n_329),
.B1(n_337),
.B2(n_308),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_296),
.Y(n_325)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_325),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_285),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_327),
.B(n_328),
.C(n_329),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_290),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_277),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_330),
.A2(n_317),
.B1(n_302),
.B2(n_316),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_306),
.B(n_282),
.Y(n_331)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_333),
.B(n_309),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_313),
.A2(n_293),
.B1(n_281),
.B2(n_278),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_334),
.A2(n_338),
.B1(n_341),
.B2(n_311),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_287),
.C(n_292),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_337),
.C(n_339),
.Y(n_355)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_312),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_336),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_292),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_273),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_274),
.Y(n_340)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_340),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_353),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_309),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_345),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_338),
.A2(n_305),
.B(n_302),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_344),
.A2(n_339),
.B(n_328),
.Y(n_362)
);

XNOR2x1_ASAP7_75t_L g345 ( 
.A(n_335),
.B(n_319),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_332),
.A2(n_308),
.B1(n_311),
.B2(n_303),
.Y(n_350)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_350),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_352),
.B(n_324),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_354),
.Y(n_360)
);

OAI21x1_ASAP7_75t_L g356 ( 
.A1(n_351),
.A2(n_305),
.B(n_341),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_356),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_352),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_344),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_359),
.B(n_366),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_362),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_333),
.C(n_326),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_348),
.C(n_355),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_349),
.B(n_261),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_365),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_347),
.B(n_346),
.Y(n_366)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_368),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_362),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_369),
.B(n_370),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_350),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_371),
.B(n_364),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_374),
.A2(n_360),
.B(n_358),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_375),
.A2(n_370),
.B(n_372),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_380),
.C(n_361),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_363),
.C(n_345),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_379),
.B(n_381),
.Y(n_382)
);

AOI31xp33_ASAP7_75t_L g380 ( 
.A1(n_373),
.A2(n_348),
.A3(n_357),
.B(n_342),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_363),
.C(n_372),
.Y(n_381)
);

AOI21x1_ASAP7_75t_L g388 ( 
.A1(n_383),
.A2(n_385),
.B(n_386),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_378),
.B(n_367),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_384),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_376),
.A2(n_357),
.B1(n_361),
.B2(n_343),
.Y(n_385)
);

NOR3x1_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_381),
.C(n_317),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_389),
.B(n_321),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_387),
.B(n_379),
.C(n_315),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_390),
.B(n_388),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_315),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_392),
.B(n_393),
.C(n_316),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_320),
.Y(n_395)
);


endmodule