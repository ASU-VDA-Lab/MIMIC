module fake_jpeg_28483_n_451 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_451);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_451;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_48),
.Y(n_128)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g109 ( 
.A(n_50),
.Y(n_109)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_57),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_17),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_20),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_26),
.A2(n_10),
.B(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_81),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_78),
.Y(n_108)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_36),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_22),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_83),
.B(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_22),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_36),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_44),
.Y(n_112)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_91),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_95),
.B(n_101),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_112),
.B(n_116),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_114),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_53),
.B(n_33),
.Y(n_116)
);

CKINVDCx12_ASAP7_75t_R g120 ( 
.A(n_85),
.Y(n_120)
);

CKINVDCx12_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_52),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_91),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_55),
.B(n_33),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_35),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_79),
.B1(n_62),
.B2(n_88),
.Y(n_143)
);

AO22x2_ASAP7_75t_L g195 ( 
.A1(n_143),
.A2(n_130),
.B1(n_131),
.B2(n_139),
.Y(n_195)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_161),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_113),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_151),
.B(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_117),
.B(n_129),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_152),
.B(n_177),
.C(n_41),
.Y(n_206)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_41),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_80),
.B1(n_51),
.B2(n_77),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_166),
.B1(n_81),
.B2(n_99),
.Y(n_192)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_118),
.A2(n_89),
.B1(n_86),
.B2(n_82),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_94),
.B(n_30),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_167),
.B(n_93),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_168),
.B(n_174),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_78),
.B1(n_45),
.B2(n_48),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_169),
.A2(n_175),
.B1(n_179),
.B2(n_108),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_173),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_172),
.A2(n_176),
.B1(n_178),
.B2(n_140),
.Y(n_201)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_54),
.B1(n_65),
.B2(n_47),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_96),
.B(n_35),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_63),
.B1(n_56),
.B2(n_73),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_206),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_183),
.A2(n_192),
.B1(n_199),
.B2(n_97),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_116),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_193),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_143),
.A2(n_93),
.B(n_30),
.C(n_31),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_190),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_41),
.C(n_33),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_171),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_183),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_102),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_173),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_131),
.B1(n_141),
.B2(n_140),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

OAI22x1_ASAP7_75t_SL g207 ( 
.A1(n_162),
.A2(n_75),
.B1(n_109),
.B2(n_105),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_109),
.B(n_107),
.Y(n_233)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_210),
.Y(n_236)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_193),
.A2(n_179),
.B1(n_169),
.B2(n_157),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_187),
.Y(n_261)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_222),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_153),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_185),
.B(n_154),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_223),
.B(n_224),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_184),
.B(n_30),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_142),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_230),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_233),
.B1(n_134),
.B2(n_195),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_147),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_191),
.B(n_35),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_29),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_235),
.A2(n_216),
.B1(n_233),
.B2(n_211),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_190),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_258),
.C(n_229),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_182),
.B(n_195),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_240),
.A2(n_220),
.B(n_215),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_245),
.B(n_29),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_182),
.B(n_188),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_247),
.B(n_212),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_195),
.B1(n_199),
.B2(n_205),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_250),
.B1(n_260),
.B2(n_219),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_197),
.B1(n_198),
.B2(n_205),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_261),
.B1(n_230),
.B2(n_212),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_160),
.B1(n_158),
.B2(n_172),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_202),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_257),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_221),
.B(n_196),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_224),
.A2(n_142),
.B(n_149),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_SL g290 ( 
.A(n_259),
.B(n_163),
.C(n_149),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_230),
.A2(n_178),
.B1(n_145),
.B2(n_146),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_238),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_265),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_239),
.Y(n_264)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_264),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_209),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_267),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_239),
.B(n_218),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_268),
.A2(n_273),
.B1(n_275),
.B2(n_282),
.Y(n_316)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_270),
.Y(n_303)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_272),
.A2(n_291),
.B1(n_202),
.B2(n_176),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_255),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_216),
.B1(n_211),
.B2(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_276),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_277),
.A2(n_279),
.B1(n_289),
.B2(n_164),
.Y(n_318)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_261),
.A2(n_233),
.B1(n_213),
.B2(n_231),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_233),
.B(n_210),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_280),
.A2(n_284),
.B(n_290),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_258),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_247),
.A2(n_214),
.B1(n_225),
.B2(n_194),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_210),
.Y(n_284)
);

NOR2x1_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_220),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_285),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_137),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_244),
.B(n_232),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_253),
.Y(n_293)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_248),
.A2(n_225),
.B1(n_194),
.B2(n_189),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_245),
.A2(n_42),
.B1(n_31),
.B2(n_44),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_300),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_277),
.A2(n_242),
.B1(n_250),
.B2(n_246),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_312),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_244),
.Y(n_297)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_297),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_272),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_314),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_237),
.C(n_236),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_271),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_255),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_315),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_262),
.C(n_279),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_278),
.C(n_276),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_313),
.A2(n_268),
.B1(n_290),
.B2(n_283),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_269),
.B(n_42),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_215),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_318),
.A2(n_289),
.B1(n_292),
.B2(n_115),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_286),
.A2(n_44),
.B1(n_28),
.B2(n_97),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_312),
.Y(n_342)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

OA21x2_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_285),
.B(n_284),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_323),
.A2(n_332),
.B(n_344),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_288),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_307),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_318),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_334),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_330),
.A2(n_320),
.B1(n_298),
.B2(n_296),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_300),
.C(n_305),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_331),
.B(n_338),
.C(n_346),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_295),
.A2(n_31),
.B(n_42),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_294),
.B(n_163),
.Y(n_334)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_337),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_123),
.C(n_126),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_303),
.Y(n_339)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_339),
.Y(n_352)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_302),
.Y(n_340)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_308),
.Y(n_341)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_341),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_342),
.A2(n_28),
.B1(n_44),
.B2(n_49),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_299),
.A2(n_103),
.B(n_106),
.Y(n_343)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_343),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_295),
.A2(n_165),
.B(n_132),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_309),
.Y(n_345)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_345),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_165),
.C(n_46),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_333),
.A2(n_316),
.B(n_307),
.Y(n_348)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_348),
.Y(n_377)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_354),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_311),
.Y(n_354)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_355),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_310),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_364),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_319),
.Y(n_359)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_359),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_360),
.A2(n_27),
.B1(n_32),
.B2(n_43),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_100),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_363),
.B(n_365),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_335),
.A2(n_66),
.B1(n_76),
.B2(n_4),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_27),
.C(n_100),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_114),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_330),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_27),
.C(n_29),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_369),
.Y(n_388)
);

OAI322xp33_ASAP7_75t_L g372 ( 
.A1(n_363),
.A2(n_323),
.A3(n_334),
.B1(n_344),
.B2(n_328),
.C1(n_338),
.C2(n_346),
.Y(n_372)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_372),
.Y(n_389)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_353),
.Y(n_373)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_347),
.A2(n_323),
.B(n_335),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_374),
.B(n_375),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_356),
.A2(n_335),
.B(n_332),
.Y(n_375)
);

XNOR2x1_ASAP7_75t_SL g379 ( 
.A(n_361),
.B(n_328),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_382),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_384),
.Y(n_393)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_357),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_368),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_352),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_367),
.A2(n_43),
.B1(n_32),
.B2(n_134),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_387),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_356),
.A2(n_43),
.B(n_32),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_377),
.A2(n_362),
.B(n_349),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_390),
.A2(n_387),
.B(n_386),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_362),
.C(n_351),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_394),
.B(n_397),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_400),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_354),
.C(n_366),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_380),
.C(n_381),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_388),
.B(n_369),
.C(n_361),
.Y(n_397)
);

INVxp33_ASAP7_75t_SL g399 ( 
.A(n_375),
.Y(n_399)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_399),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_365),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_364),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_383),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_350),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_403),
.B(n_370),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_410),
.C(n_416),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_407),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_403),
.B(n_370),
.C(n_371),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_399),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_412),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_389),
.A2(n_392),
.B1(n_398),
.B2(n_391),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_393),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_396),
.B(n_371),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_415),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_414),
.A2(n_58),
.B(n_37),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_392),
.B(n_373),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_SL g419 ( 
.A(n_409),
.B(n_401),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_419),
.B(n_9),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_401),
.C(n_13),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_423),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_12),
.C(n_17),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_425),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_11),
.C(n_15),
.Y(n_425)
);

AO21x1_ASAP7_75t_L g426 ( 
.A1(n_411),
.A2(n_11),
.B(n_15),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_426),
.B(n_8),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_408),
.C(n_12),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_427),
.B(n_9),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_9),
.C(n_14),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_428),
.B(n_430),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_429),
.Y(n_441)
);

OAI321xp33_ASAP7_75t_L g439 ( 
.A1(n_431),
.A2(n_5),
.A3(n_2),
.B1(n_0),
.B2(n_39),
.C(n_37),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_14),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_432),
.B(n_433),
.C(n_436),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_7),
.C(n_4),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_16),
.C(n_5),
.Y(n_436)
);

OAI21x1_ASAP7_75t_SL g437 ( 
.A1(n_434),
.A2(n_417),
.B(n_7),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_L g445 ( 
.A1(n_437),
.A2(n_439),
.B(n_442),
.C(n_0),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_431),
.A2(n_37),
.B(n_38),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_441),
.B(n_435),
.C(n_38),
.Y(n_443)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_443),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_438),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_444),
.A2(n_445),
.B(n_440),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_447),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_446),
.Y(n_449)
);

AND2x4_ASAP7_75t_SL g450 ( 
.A(n_449),
.B(n_2),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_2),
.Y(n_451)
);


endmodule