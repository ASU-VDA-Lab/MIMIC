module real_aes_7641_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g463 ( .A1(n_0), .A2(n_141), .B(n_464), .C(n_467), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_1), .B(n_458), .Y(n_469) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_2), .B(n_88), .C(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g432 ( .A(n_2), .Y(n_432) );
INVx1_ASAP7_75t_L g179 ( .A(n_3), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_4), .B(n_142), .Y(n_541) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_5), .A2(n_120), .B1(n_121), .B2(n_427), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g427 ( .A(n_5), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_5), .A2(n_95), .B1(n_427), .B2(n_736), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_6), .A2(n_443), .B(n_490), .Y(n_489) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_7), .A2(n_148), .B(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_8), .A2(n_37), .B1(n_145), .B2(n_197), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_9), .A2(n_103), .B1(n_112), .B2(n_745), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_10), .B(n_148), .Y(n_165) );
AND2x6_ASAP7_75t_L g150 ( .A(n_11), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_12), .A2(n_150), .B(n_446), .C(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_13), .B(n_39), .Y(n_106) );
INVx1_ASAP7_75t_L g132 ( .A(n_14), .Y(n_132) );
INVx1_ASAP7_75t_L g171 ( .A(n_15), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_16), .B(n_138), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_17), .B(n_142), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_18), .B(n_128), .Y(n_127) );
AO32x2_ASAP7_75t_L g208 ( .A1(n_19), .A2(n_148), .A3(n_149), .B1(n_168), .B2(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_20), .B(n_145), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_21), .B(n_128), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_22), .A2(n_55), .B1(n_145), .B2(n_197), .Y(n_211) );
AOI22xp33_ASAP7_75t_SL g205 ( .A1(n_23), .A2(n_80), .B1(n_138), .B2(n_145), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_24), .B(n_145), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_25), .A2(n_149), .B(n_446), .C(n_448), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_26), .A2(n_149), .B(n_446), .C(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_27), .Y(n_136) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_28), .A2(n_96), .B1(n_115), .B2(n_116), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_28), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_29), .B(n_187), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_30), .A2(n_443), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_31), .B(n_187), .Y(n_224) );
INVx2_ASAP7_75t_L g140 ( .A(n_32), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_33), .A2(n_478), .B(n_479), .C(n_483), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_34), .B(n_145), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_35), .B(n_187), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_36), .B(n_193), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_38), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_40), .B(n_442), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_41), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_42), .B(n_142), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_43), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_44), .B(n_443), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_45), .A2(n_478), .B(n_483), .C(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_46), .B(n_145), .Y(n_158) );
INVx1_ASAP7_75t_L g465 ( .A(n_47), .Y(n_465) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_48), .A2(n_734), .B1(n_737), .B2(n_738), .Y(n_733) );
INVx1_ASAP7_75t_L g738 ( .A(n_48), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_49), .A2(n_89), .B1(n_197), .B2(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g504 ( .A(n_50), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_51), .B(n_145), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_52), .B(n_145), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_53), .B(n_443), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_54), .B(n_163), .Y(n_162) );
AOI22xp33_ASAP7_75t_SL g144 ( .A1(n_56), .A2(n_60), .B1(n_138), .B2(n_145), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_57), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_58), .B(n_145), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_59), .B(n_145), .Y(n_244) );
INVx1_ASAP7_75t_L g151 ( .A(n_61), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_62), .B(n_443), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_63), .B(n_458), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_64), .A2(n_163), .B(n_174), .C(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_65), .B(n_145), .Y(n_180) );
INVx1_ASAP7_75t_L g131 ( .A(n_66), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_67), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_68), .B(n_142), .Y(n_481) );
AO32x2_ASAP7_75t_L g201 ( .A1(n_69), .A2(n_148), .A3(n_149), .B1(n_202), .B2(n_206), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_70), .B(n_143), .Y(n_515) );
INVx1_ASAP7_75t_L g243 ( .A(n_71), .Y(n_243) );
INVx1_ASAP7_75t_L g219 ( .A(n_72), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_73), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_74), .B(n_450), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_75), .A2(n_446), .B(n_483), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_76), .B(n_138), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_77), .Y(n_491) );
INVx1_ASAP7_75t_L g111 ( .A(n_78), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_79), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_81), .B(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_82), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_83), .B(n_138), .Y(n_223) );
INVx2_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_85), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_86), .B(n_135), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_87), .B(n_138), .Y(n_159) );
OR2x2_ASAP7_75t_L g430 ( .A(n_88), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g718 ( .A(n_88), .Y(n_718) );
OR2x2_ASAP7_75t_L g732 ( .A(n_88), .B(n_726), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g137 ( .A1(n_90), .A2(n_101), .B1(n_138), .B2(n_139), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_91), .B(n_443), .Y(n_476) );
INVx1_ASAP7_75t_L g480 ( .A(n_92), .Y(n_480) );
INVxp67_ASAP7_75t_L g494 ( .A(n_93), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_94), .B(n_138), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_95), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_96), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_97), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g511 ( .A(n_98), .Y(n_511) );
INVx1_ASAP7_75t_L g540 ( .A(n_99), .Y(n_540) );
AND2x2_ASAP7_75t_L g506 ( .A(n_100), .B(n_187), .Y(n_506) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g745 ( .A(n_105), .Y(n_745) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
AND2x2_ASAP7_75t_L g431 ( .A(n_106), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AO221x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_727), .B1(n_730), .B2(n_739), .C(n_741), .Y(n_112) );
OAI222xp33_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_117), .B1(n_719), .B2(n_720), .C1(n_723), .C2(n_724), .Y(n_113) );
INVx1_ASAP7_75t_L g719 ( .A(n_114), .Y(n_719) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_428), .B1(n_433), .B2(n_715), .Y(n_118) );
INVx1_ASAP7_75t_L g722 ( .A(n_119), .Y(n_722) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
XNOR2xp5_ASAP7_75t_L g734 ( .A(n_121), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_SL g121 ( .A(n_122), .B(n_361), .Y(n_121) );
NOR5xp2_ASAP7_75t_L g122 ( .A(n_123), .B(n_274), .C(n_320), .D(n_333), .E(n_345), .Y(n_122) );
OAI211xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_182), .B(n_228), .C(n_255), .Y(n_123) );
INVx1_ASAP7_75t_SL g356 ( .A(n_124), .Y(n_356) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_152), .Y(n_124) );
AND2x2_ASAP7_75t_L g280 ( .A(n_125), .B(n_153), .Y(n_280) );
AND2x2_ASAP7_75t_L g308 ( .A(n_125), .B(n_254), .Y(n_308) );
AND2x2_ASAP7_75t_L g316 ( .A(n_125), .B(n_259), .Y(n_316) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g246 ( .A(n_126), .B(n_154), .Y(n_246) );
INVx2_ASAP7_75t_L g258 ( .A(n_126), .Y(n_258) );
AND2x2_ASAP7_75t_L g383 ( .A(n_126), .B(n_325), .Y(n_383) );
OR2x2_ASAP7_75t_L g385 ( .A(n_126), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_133), .Y(n_126) );
INVx1_ASAP7_75t_L g252 ( .A(n_127), .Y(n_252) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_128), .Y(n_148) );
INVx1_ASAP7_75t_L g168 ( .A(n_128), .Y(n_168) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_129), .B(n_130), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
NAND3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_147), .C(n_149), .Y(n_133) );
AO21x1_ASAP7_75t_L g251 ( .A1(n_134), .A2(n_147), .B(n_252), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_137), .B1(n_141), .B2(n_144), .Y(n_134) );
INVx2_ASAP7_75t_L g198 ( .A(n_135), .Y(n_198) );
OAI22xp5_ASAP7_75t_SL g202 ( .A1(n_135), .A2(n_143), .B1(n_203), .B2(n_205), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_135), .A2(n_141), .B1(n_210), .B2(n_211), .Y(n_209) );
INVx4_ASAP7_75t_L g466 ( .A(n_135), .Y(n_466) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx3_ASAP7_75t_L g143 ( .A(n_136), .Y(n_143) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
INVx1_ASAP7_75t_L g193 ( .A(n_136), .Y(n_193) );
AND2x2_ASAP7_75t_L g444 ( .A(n_136), .B(n_164), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_136), .Y(n_447) );
INVx2_ASAP7_75t_L g172 ( .A(n_138), .Y(n_172) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
INVx1_ASAP7_75t_L g164 ( .A(n_140), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_141), .A2(n_161), .B(n_162), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_141), .A2(n_178), .B(n_179), .C(n_180), .Y(n_177) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_142), .A2(n_158), .B(n_159), .Y(n_157) );
O2A1O1Ixp5_ASAP7_75t_SL g217 ( .A1(n_142), .A2(n_218), .B(n_219), .C(n_220), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_142), .A2(n_240), .B(n_241), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_142), .B(n_494), .Y(n_493) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx3_ASAP7_75t_L g218 ( .A(n_145), .Y(n_218) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_145), .Y(n_542) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g197 ( .A(n_146), .Y(n_197) );
BUFx3_ASAP7_75t_L g204 ( .A(n_146), .Y(n_204) );
AND2x6_ASAP7_75t_L g446 ( .A(n_146), .B(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g458 ( .A(n_147), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_147), .B(n_485), .Y(n_484) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_147), .A2(n_510), .B(n_517), .Y(n_509) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_147), .A2(n_537), .B(n_544), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_147), .B(n_545), .Y(n_544) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_148), .A2(n_156), .B(n_165), .Y(n_155) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_148), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_148), .A2(n_522), .B(n_523), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_149), .A2(n_239), .B(n_242), .Y(n_238) );
BUFx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI21xp5_ASAP7_75t_L g156 ( .A1(n_150), .A2(n_157), .B(n_160), .Y(n_156) );
OAI21xp5_ASAP7_75t_L g169 ( .A1(n_150), .A2(n_170), .B(n_177), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_150), .A2(n_189), .B(n_194), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_150), .A2(n_217), .B(n_221), .Y(n_216) );
AND2x4_ASAP7_75t_L g443 ( .A(n_150), .B(n_444), .Y(n_443) );
INVx4_ASAP7_75t_SL g468 ( .A(n_150), .Y(n_468) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_150), .B(n_444), .Y(n_512) );
INVx2_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g296 ( .A(n_153), .B(n_268), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_153), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g410 ( .A(n_153), .B(n_250), .Y(n_410) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_166), .Y(n_153) );
AND2x2_ASAP7_75t_L g253 ( .A(n_154), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g300 ( .A(n_154), .Y(n_300) );
AND2x2_ASAP7_75t_L g325 ( .A(n_154), .B(n_237), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_154), .B(n_358), .Y(n_395) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_L g259 ( .A(n_155), .B(n_237), .Y(n_259) );
AND2x2_ASAP7_75t_L g273 ( .A(n_155), .B(n_236), .Y(n_273) );
AND2x2_ASAP7_75t_L g290 ( .A(n_155), .B(n_166), .Y(n_290) );
AND2x2_ASAP7_75t_L g347 ( .A(n_155), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_155), .B(n_254), .Y(n_360) );
AND2x2_ASAP7_75t_L g412 ( .A(n_155), .B(n_337), .Y(n_412) );
INVx2_ASAP7_75t_L g178 ( .A(n_163), .Y(n_178) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g235 ( .A(n_166), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g254 ( .A(n_166), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_166), .B(n_237), .Y(n_331) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B(n_181), .Y(n_166) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_167), .A2(n_238), .B(n_245), .Y(n_237) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_168), .B(n_518), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_173), .C(n_174), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_172), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_172), .A2(n_525), .B(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_174), .A2(n_540), .B(n_541), .C(n_542), .Y(n_539) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_175), .A2(n_222), .B(n_223), .Y(n_221) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g450 ( .A(n_176), .Y(n_450) );
O2A1O1Ixp5_ASAP7_75t_L g242 ( .A1(n_178), .A2(n_198), .B(n_243), .C(n_244), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_178), .A2(n_449), .B(n_451), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_212), .B(n_225), .Y(n_182) );
INVx1_ASAP7_75t_SL g344 ( .A(n_183), .Y(n_344) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_200), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_SL g232 ( .A(n_185), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g227 ( .A(n_186), .Y(n_227) );
INVx1_ASAP7_75t_L g264 ( .A(n_186), .Y(n_264) );
AND2x2_ASAP7_75t_L g285 ( .A(n_186), .B(n_207), .Y(n_285) );
AND2x2_ASAP7_75t_L g319 ( .A(n_186), .B(n_208), .Y(n_319) );
OR2x2_ASAP7_75t_L g338 ( .A(n_186), .B(n_214), .Y(n_338) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_186), .Y(n_352) );
AND2x2_ASAP7_75t_L g365 ( .A(n_186), .B(n_366), .Y(n_365) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_199), .Y(n_186) );
INVx2_ASAP7_75t_L g206 ( .A(n_187), .Y(n_206) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_187), .A2(n_216), .B(n_224), .Y(n_215) );
INVx1_ASAP7_75t_L g456 ( .A(n_187), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_187), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_187), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_192), .Y(n_189) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_198), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_200), .A2(n_287), .B1(n_288), .B2(n_297), .Y(n_286) );
AND2x2_ASAP7_75t_L g370 ( .A(n_200), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_207), .Y(n_200) );
INVx1_ASAP7_75t_L g231 ( .A(n_201), .Y(n_231) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_201), .Y(n_268) );
INVx1_ASAP7_75t_L g279 ( .A(n_201), .Y(n_279) );
AND2x2_ASAP7_75t_L g294 ( .A(n_201), .B(n_208), .Y(n_294) );
INVx2_ASAP7_75t_L g467 ( .A(n_204), .Y(n_467) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_204), .Y(n_482) );
INVx1_ASAP7_75t_L g453 ( .A(n_206), .Y(n_453) );
OR2x2_ASAP7_75t_L g248 ( .A(n_207), .B(n_233), .Y(n_248) );
AND2x2_ASAP7_75t_L g278 ( .A(n_207), .B(n_279), .Y(n_278) );
NOR2xp67_ASAP7_75t_L g366 ( .A(n_207), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g226 ( .A(n_208), .B(n_227), .Y(n_226) );
BUFx2_ASAP7_75t_L g335 ( .A(n_208), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_212), .B(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g313 ( .A(n_213), .B(n_279), .Y(n_313) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g225 ( .A(n_214), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g284 ( .A(n_214), .Y(n_284) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g233 ( .A(n_215), .Y(n_233) );
OR2x2_ASAP7_75t_L g263 ( .A(n_215), .B(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_215), .Y(n_318) );
AOI32xp33_ASAP7_75t_L g355 ( .A1(n_225), .A2(n_285), .A3(n_356), .B1(n_357), .B2(n_359), .Y(n_355) );
AND2x2_ASAP7_75t_L g281 ( .A(n_226), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_226), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_226), .B(n_313), .Y(n_399) );
INVx1_ASAP7_75t_L g404 ( .A(n_226), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_234), .B1(n_247), .B2(n_249), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
AND2x2_ASAP7_75t_L g334 ( .A(n_230), .B(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_231), .B(n_233), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_232), .A2(n_256), .B1(n_260), .B2(n_270), .Y(n_255) );
AND2x2_ASAP7_75t_L g277 ( .A(n_232), .B(n_278), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g328 ( .A1(n_232), .A2(n_246), .B(n_294), .C(n_329), .Y(n_328) );
OAI332xp33_ASAP7_75t_L g333 ( .A1(n_232), .A2(n_334), .A3(n_336), .B1(n_338), .B2(n_339), .B3(n_341), .C1(n_342), .C2(n_344), .Y(n_333) );
INVx2_ASAP7_75t_L g374 ( .A(n_232), .Y(n_374) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_233), .Y(n_292) );
INVx1_ASAP7_75t_L g367 ( .A(n_233), .Y(n_367) );
AND2x2_ASAP7_75t_L g421 ( .A(n_233), .B(n_285), .Y(n_421) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_246), .Y(n_234) );
AND2x2_ASAP7_75t_L g301 ( .A(n_236), .B(n_251), .Y(n_301) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g250 ( .A(n_237), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g349 ( .A(n_237), .B(n_251), .Y(n_349) );
INVx1_ASAP7_75t_L g358 ( .A(n_237), .Y(n_358) );
INVx1_ASAP7_75t_L g332 ( .A(n_246), .Y(n_332) );
INVxp67_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g416 ( .A(n_248), .B(n_268), .Y(n_416) );
INVx1_ASAP7_75t_SL g327 ( .A(n_249), .Y(n_327) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_253), .Y(n_249) );
AND2x2_ASAP7_75t_L g354 ( .A(n_250), .B(n_312), .Y(n_354) );
INVx1_ASAP7_75t_L g373 ( .A(n_250), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_250), .B(n_340), .Y(n_375) );
INVx1_ASAP7_75t_L g272 ( .A(n_251), .Y(n_272) );
AND2x2_ASAP7_75t_L g276 ( .A(n_253), .B(n_257), .Y(n_276) );
AND2x2_ASAP7_75t_L g343 ( .A(n_253), .B(n_301), .Y(n_343) );
INVx2_ASAP7_75t_L g386 ( .A(n_253), .Y(n_386) );
INVx2_ASAP7_75t_L g269 ( .A(n_254), .Y(n_269) );
AND2x2_ASAP7_75t_L g271 ( .A(n_254), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
INVx1_ASAP7_75t_L g287 ( .A(n_257), .Y(n_287) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_258), .B(n_331), .Y(n_337) );
OR2x2_ASAP7_75t_L g401 ( .A(n_258), .B(n_360), .Y(n_401) );
INVx1_ASAP7_75t_L g425 ( .A(n_258), .Y(n_425) );
INVx1_ASAP7_75t_L g381 ( .A(n_259), .Y(n_381) );
AND2x2_ASAP7_75t_L g426 ( .A(n_259), .B(n_269), .Y(n_426) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_263), .A2(n_289), .B1(n_291), .B2(n_295), .Y(n_288) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI322xp33_ASAP7_75t_SL g372 ( .A1(n_266), .A2(n_373), .A3(n_374), .B1(n_375), .B2(n_376), .C1(n_379), .C2(n_381), .Y(n_372) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
AND2x2_ASAP7_75t_L g369 ( .A(n_267), .B(n_285), .Y(n_369) );
OR2x2_ASAP7_75t_L g403 ( .A(n_267), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g406 ( .A(n_267), .B(n_338), .Y(n_406) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g351 ( .A(n_268), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g407 ( .A(n_268), .B(n_338), .Y(n_407) );
INVx3_ASAP7_75t_L g340 ( .A(n_269), .Y(n_340) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g396 ( .A(n_271), .Y(n_396) );
AOI222xp33_ASAP7_75t_L g275 ( .A1(n_273), .A2(n_276), .B1(n_277), .B2(n_280), .C1(n_281), .C2(n_283), .Y(n_275) );
INVx1_ASAP7_75t_L g306 ( .A(n_273), .Y(n_306) );
NAND3xp33_ASAP7_75t_SL g274 ( .A(n_275), .B(n_286), .C(n_303), .Y(n_274) );
AND2x2_ASAP7_75t_L g391 ( .A(n_278), .B(n_292), .Y(n_391) );
BUFx2_ASAP7_75t_L g282 ( .A(n_279), .Y(n_282) );
INVx1_ASAP7_75t_L g323 ( .A(n_279), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_280), .A2(n_316), .B1(n_369), .B2(n_370), .C(n_372), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_282), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_285), .Y(n_309) );
AND2x2_ASAP7_75t_L g322 ( .A(n_285), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_290), .B(n_301), .Y(n_302) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
OAI21xp33_ASAP7_75t_L g297 ( .A1(n_292), .A2(n_298), .B(n_302), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_292), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g389 ( .A(n_294), .B(n_371), .Y(n_389) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g312 ( .A(n_300), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_301), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g418 ( .A(n_301), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_309), .B1(n_310), .B2(n_313), .C(n_314), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_305), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g414 ( .A(n_313), .B(n_319), .Y(n_414) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
OAI31xp33_ASAP7_75t_SL g382 ( .A1(n_317), .A2(n_356), .A3(n_383), .B(n_384), .Y(n_382) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g371 ( .A(n_318), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_319), .B(n_323), .Y(n_422) );
OAI221xp5_ASAP7_75t_SL g320 ( .A1(n_321), .A2(n_324), .B1(n_326), .B2(n_327), .C(n_328), .Y(n_320) );
INVx1_ASAP7_75t_L g326 ( .A(n_322), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_325), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g341 ( .A(n_334), .Y(n_341) );
INVx2_ASAP7_75t_L g377 ( .A(n_335), .Y(n_377) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g363 ( .A(n_340), .B(n_349), .Y(n_363) );
A2O1A1Ixp33_ASAP7_75t_L g413 ( .A1(n_340), .A2(n_357), .B(n_414), .C(n_415), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g345 ( .A1(n_341), .A2(n_346), .B1(n_350), .B2(n_353), .C(n_355), .Y(n_345) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
A2O1A1Ixp33_ASAP7_75t_L g408 ( .A1(n_344), .A2(n_409), .B(n_411), .C(n_413), .Y(n_408) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_347), .A2(n_398), .B1(n_400), .B2(n_402), .C(n_405), .Y(n_397) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
NOR4xp25_ASAP7_75t_L g361 ( .A(n_362), .B(n_387), .C(n_408), .D(n_419), .Y(n_361) );
OAI211xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_364), .B(n_368), .C(n_382), .Y(n_362) );
INVx1_ASAP7_75t_SL g417 ( .A(n_369), .Y(n_417) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_SL g380 ( .A(n_378), .Y(n_380) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_385), .A2(n_394), .B1(n_406), .B2(n_407), .Y(n_405) );
A2O1A1Ixp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B(n_392), .C(n_397), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI31xp33_ASAP7_75t_L g419 ( .A1(n_390), .A2(n_420), .A3(n_422), .B(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_417), .B(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_430), .A2(n_434), .B1(n_717), .B2(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g717 ( .A(n_431), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g726 ( .A(n_431), .Y(n_726) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_SL g434 ( .A(n_435), .B(n_651), .Y(n_434) );
NOR5xp2_ASAP7_75t_L g435 ( .A(n_436), .B(n_582), .C(n_611), .D(n_631), .E(n_638), .Y(n_435) );
OAI211xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_470), .B(n_527), .C(n_569), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_438), .A2(n_654), .B1(n_656), .B2(n_657), .Y(n_653) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_457), .Y(n_438) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_439), .Y(n_530) );
AND2x4_ASAP7_75t_L g562 ( .A(n_439), .B(n_563), .Y(n_562) );
INVx5_ASAP7_75t_L g580 ( .A(n_439), .Y(n_580) );
AND2x2_ASAP7_75t_L g589 ( .A(n_439), .B(n_581), .Y(n_589) );
AND2x2_ASAP7_75t_L g601 ( .A(n_439), .B(n_474), .Y(n_601) );
AND2x2_ASAP7_75t_L g697 ( .A(n_439), .B(n_565), .Y(n_697) );
OR2x6_ASAP7_75t_L g439 ( .A(n_440), .B(n_454), .Y(n_439) );
AOI21xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_445), .B(n_453), .Y(n_440) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx5_ASAP7_75t_L g462 ( .A(n_446), .Y(n_462) );
INVx2_ASAP7_75t_L g452 ( .A(n_450), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_452), .A2(n_480), .B(n_481), .C(n_482), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_452), .A2(n_482), .B(n_504), .C(n_505), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx2_ASAP7_75t_L g563 ( .A(n_457), .Y(n_563) );
AND2x2_ASAP7_75t_L g581 ( .A(n_457), .B(n_536), .Y(n_581) );
AND2x2_ASAP7_75t_L g600 ( .A(n_457), .B(n_535), .Y(n_600) );
AND2x2_ASAP7_75t_L g640 ( .A(n_457), .B(n_580), .Y(n_640) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_469), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_462), .B(n_463), .C(n_468), .Y(n_460) );
INVx2_ASAP7_75t_L g478 ( .A(n_462), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_462), .A2(n_468), .B(n_491), .C(n_492), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g483 ( .A(n_468), .Y(n_483) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_496), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AOI322xp5_ASAP7_75t_L g699 ( .A1(n_473), .A2(n_507), .A3(n_554), .B1(n_562), .B2(n_616), .C1(n_700), .C2(n_703), .Y(n_699) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_486), .Y(n_473) );
INVx5_ASAP7_75t_L g532 ( .A(n_474), .Y(n_532) );
AND2x2_ASAP7_75t_L g548 ( .A(n_474), .B(n_534), .Y(n_548) );
BUFx2_ASAP7_75t_L g626 ( .A(n_474), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_474), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g703 ( .A(n_474), .B(n_610), .Y(n_703) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_486), .B(n_498), .Y(n_557) );
INVx1_ASAP7_75t_L g584 ( .A(n_486), .Y(n_584) );
AND2x2_ASAP7_75t_L g597 ( .A(n_486), .B(n_519), .Y(n_597) );
AND2x2_ASAP7_75t_L g698 ( .A(n_486), .B(n_616), .Y(n_698) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g552 ( .A(n_487), .B(n_498), .Y(n_552) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_487), .Y(n_560) );
OR2x2_ASAP7_75t_L g567 ( .A(n_487), .B(n_519), .Y(n_567) );
AND2x2_ASAP7_75t_L g577 ( .A(n_487), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_487), .B(n_509), .Y(n_606) );
INVxp67_ASAP7_75t_L g630 ( .A(n_487), .Y(n_630) );
AND2x2_ASAP7_75t_L g637 ( .A(n_487), .B(n_507), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_487), .B(n_519), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_487), .B(n_508), .Y(n_663) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B(n_495), .Y(n_487) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_498), .B(n_520), .Y(n_607) );
OR2x2_ASAP7_75t_L g629 ( .A(n_498), .B(n_508), .Y(n_629) );
AND2x2_ASAP7_75t_L g642 ( .A(n_498), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_498), .B(n_597), .Y(n_648) );
OAI211xp5_ASAP7_75t_SL g652 ( .A1(n_498), .A2(n_653), .B(n_658), .C(n_667), .Y(n_652) );
AND2x2_ASAP7_75t_L g713 ( .A(n_498), .B(n_519), .Y(n_713) );
INVx5_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g566 ( .A(n_499), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_499), .B(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_499), .B(n_561), .Y(n_573) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_499), .Y(n_575) );
OR2x2_ASAP7_75t_L g586 ( .A(n_499), .B(n_508), .Y(n_586) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_499), .B(n_577), .Y(n_591) );
AND2x2_ASAP7_75t_L g616 ( .A(n_499), .B(n_508), .Y(n_616) );
AND2x2_ASAP7_75t_L g636 ( .A(n_499), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g674 ( .A(n_499), .B(n_507), .Y(n_674) );
OR2x2_ASAP7_75t_L g677 ( .A(n_499), .B(n_663), .Y(n_677) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_506), .Y(n_499) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_519), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g620 ( .A1(n_508), .A2(n_621), .B(n_624), .C(n_630), .Y(n_620) );
INVx5_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_509), .B(n_519), .Y(n_551) );
AND2x2_ASAP7_75t_L g555 ( .A(n_509), .B(n_520), .Y(n_555) );
OR2x2_ASAP7_75t_L g561 ( .A(n_509), .B(n_519), .Y(n_561) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_513), .Y(n_510) );
INVx1_ASAP7_75t_SL g578 ( .A(n_519), .Y(n_578) );
OR2x2_ASAP7_75t_L g706 ( .A(n_519), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_546), .B(n_549), .C(n_558), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AOI31xp33_ASAP7_75t_L g631 ( .A1(n_529), .A2(n_632), .A3(n_634), .B(n_635), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_530), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_531), .B(n_562), .Y(n_568) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_532), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g588 ( .A(n_532), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g593 ( .A(n_532), .B(n_563), .Y(n_593) );
AND2x2_ASAP7_75t_L g603 ( .A(n_532), .B(n_562), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_532), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g623 ( .A(n_532), .B(n_580), .Y(n_623) );
AND2x2_ASAP7_75t_L g628 ( .A(n_532), .B(n_600), .Y(n_628) );
OR2x2_ASAP7_75t_L g647 ( .A(n_532), .B(n_534), .Y(n_647) );
OR2x2_ASAP7_75t_L g649 ( .A(n_532), .B(n_650), .Y(n_649) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_532), .Y(n_696) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g596 ( .A(n_534), .B(n_563), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_534), .B(n_580), .Y(n_619) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g565 ( .A(n_536), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_543), .Y(n_537) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g656 ( .A(n_548), .B(n_580), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g658 ( .A1(n_548), .A2(n_562), .A3(n_600), .B1(n_659), .B2(n_660), .C1(n_661), .C2(n_664), .Y(n_658) );
INVx1_ASAP7_75t_L g666 ( .A(n_548), .Y(n_666) );
NAND2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx1_ASAP7_75t_SL g660 ( .A(n_550), .Y(n_660) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
OR2x2_ASAP7_75t_L g612 ( .A(n_551), .B(n_557), .Y(n_612) );
INVx1_ASAP7_75t_L g643 ( .A(n_551), .Y(n_643) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI32xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .A3(n_564), .B1(n_566), .B2(n_568), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AOI21xp33_ASAP7_75t_SL g598 ( .A1(n_561), .A2(n_576), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_SL g613 ( .A(n_562), .Y(n_613) );
AND2x4_ASAP7_75t_L g610 ( .A(n_563), .B(n_580), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_563), .B(n_646), .Y(n_645) );
AOI322xp5_ASAP7_75t_L g675 ( .A1(n_564), .A2(n_591), .A3(n_610), .B1(n_643), .B2(n_676), .C1(n_678), .C2(n_679), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_564), .A2(n_641), .B1(n_705), .B2(n_706), .C(n_708), .Y(n_704) );
AND2x2_ASAP7_75t_L g592 ( .A(n_565), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_SL g572 ( .A(n_567), .Y(n_572) );
OR2x2_ASAP7_75t_L g644 ( .A(n_567), .B(n_629), .Y(n_644) );
OAI31xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_573), .A3(n_574), .B(n_579), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_570), .A2(n_603), .B1(n_604), .B2(n_608), .Y(n_602) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g615 ( .A(n_572), .B(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_574), .A2(n_615), .B1(n_668), .B2(n_671), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g657 ( .A(n_577), .B(n_626), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_577), .B(n_616), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_578), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g691 ( .A(n_578), .B(n_629), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_579), .A2(n_674), .B1(n_687), .B2(n_690), .Y(n_686) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx2_ASAP7_75t_L g595 ( .A(n_580), .Y(n_595) );
AND2x2_ASAP7_75t_L g678 ( .A(n_580), .B(n_600), .Y(n_678) );
OR2x2_ASAP7_75t_L g680 ( .A(n_580), .B(n_647), .Y(n_680) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_580), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_581), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_581), .B(n_626), .Y(n_634) );
OAI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_587), .B(n_590), .C(n_602), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_594), .B2(n_597), .C(n_598), .Y(n_590) );
INVxp67_ASAP7_75t_L g702 ( .A(n_593), .Y(n_702) );
INVx1_ASAP7_75t_L g669 ( .A(n_594), .Y(n_669) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AND2x2_ASAP7_75t_L g633 ( .A(n_595), .B(n_600), .Y(n_633) );
INVx1_ASAP7_75t_L g650 ( .A(n_596), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_596), .B(n_623), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g665 ( .A(n_600), .Y(n_665) );
AND2x2_ASAP7_75t_L g671 ( .A(n_600), .B(n_626), .Y(n_671) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_SL g659 ( .A(n_607), .Y(n_659) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_610), .B(n_646), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B1(n_614), .B2(n_617), .C(n_620), .Y(n_611) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g707 ( .A(n_616), .Y(n_707) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g625 ( .A(n_619), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_623), .B(n_682), .Y(n_681) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B(n_629), .Y(n_624) );
OAI211xp5_ASAP7_75t_SL g672 ( .A1(n_627), .A2(n_673), .B(n_675), .C(n_681), .Y(n_672) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g684 ( .A(n_629), .Y(n_684) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI222xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B1(n_644), .B2(n_645), .C1(n_648), .C2(n_649), .Y(n_638) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g714 ( .A(n_645), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_646), .B(n_689), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_646), .A2(n_693), .B1(n_695), .B2(n_698), .Y(n_692) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
NOR4xp25_ASAP7_75t_L g651 ( .A(n_652), .B(n_672), .C(n_685), .D(n_704), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_654), .B(n_684), .Y(n_694) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g661 ( .A(n_659), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_662), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_692), .C(n_699), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx2_ASAP7_75t_L g701 ( .A(n_697), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
OAI21xp5_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_711), .B(n_714), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NOR2x2_ASAP7_75t_L g725 ( .A(n_718), .B(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
BUFx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_SL g740 ( .A(n_728), .Y(n_740) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g744 ( .A(n_732), .Y(n_744) );
INVx1_ASAP7_75t_L g737 ( .A(n_734), .Y(n_737) );
BUFx3_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
endmodule