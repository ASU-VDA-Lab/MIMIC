module fake_netlist_6_3622_n_2141 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2141);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2141;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_90),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_63),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_155),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_127),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_136),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_98),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_28),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_118),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_34),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_199),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_187),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_179),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_83),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_128),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_46),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_124),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_75),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_76),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_103),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_7),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_157),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_125),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_146),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_193),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_22),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_64),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_5),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_75),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_154),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_7),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_121),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_107),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_67),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_76),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_167),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_202),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_86),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_184),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_109),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_45),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_117),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_5),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_181),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_15),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_190),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_6),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_168),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_100),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_93),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_71),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_96),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_78),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_137),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_34),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_22),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_60),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_55),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_51),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_205),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_139),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_82),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_0),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_0),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_91),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_79),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_108),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_68),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_64),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_158),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_70),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_106),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_26),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_11),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_122),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_66),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_12),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_6),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_148),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_182),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_88),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_101),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_85),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_4),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_12),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_131),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_63),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_185),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_57),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_134),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_57),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_175),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_188),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_49),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_56),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_142),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_49),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_169),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_166),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_16),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_35),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_11),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_73),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_84),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_2),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_39),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_52),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_113),
.Y(n_323)
);

BUFx8_ASAP7_75t_SL g324 ( 
.A(n_114),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_162),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_80),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_132),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_42),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_204),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_8),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_195),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_145),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_51),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_27),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_165),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_197),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_66),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_89),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_52),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_8),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_111),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_140),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_126),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_104),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_156),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_152),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_21),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_24),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_25),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_129),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_40),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_25),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_200),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_186),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_24),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_44),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_62),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_194),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_27),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_37),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_26),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_21),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_72),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_54),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_3),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_32),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_172),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_178),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_36),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_56),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_177),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_81),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_170),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_70),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_9),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_77),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_38),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_198),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_19),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_133),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_65),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_40),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_9),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_58),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_46),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_67),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_102),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_50),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_163),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_60),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_116),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_17),
.Y(n_392)
);

INVxp33_ASAP7_75t_SL g393 ( 
.A(n_14),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_29),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_130),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_196),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_2),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_1),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_13),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_31),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_10),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_3),
.Y(n_402)
);

BUFx4f_ASAP7_75t_SL g403 ( 
.A(n_18),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_30),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_97),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_324),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_260),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_210),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_244),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_244),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_213),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_244),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_215),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_232),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_244),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_244),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_217),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_244),
.Y(n_418)
);

NAND2xp33_ASAP7_75t_R g419 ( 
.A(n_393),
.B(n_1),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_244),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_216),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_218),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_222),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_244),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_244),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_232),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_232),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_232),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_232),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_223),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_251),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_225),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_287),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_258),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_346),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_258),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_391),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_258),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_258),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_258),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_249),
.B(n_4),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_226),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_264),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_227),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_229),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_290),
.B(n_319),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_278),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_236),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_260),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_264),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_268),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_278),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_239),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_278),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_278),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_240),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_245),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_278),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_288),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_369),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_247),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_248),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_349),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_253),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_366),
.B(n_10),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_255),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_257),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_261),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_265),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_379),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_288),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_267),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_269),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_369),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_275),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_276),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_212),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_369),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_369),
.Y(n_479)
);

INVxp33_ASAP7_75t_SL g480 ( 
.A(n_230),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_369),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_361),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_280),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_361),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_361),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_270),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g487 ( 
.A(n_224),
.B(n_13),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_281),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_285),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_270),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_296),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_221),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_318),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_297),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_303),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_313),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_268),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_373),
.B(n_14),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_314),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_323),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_325),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_373),
.B(n_15),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_327),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_332),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_336),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_277),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_318),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_342),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_334),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_208),
.B(n_16),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_334),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_426),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_414),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_409),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_441),
.B(n_259),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_414),
.B(n_405),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_426),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_410),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_427),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_414),
.B(n_277),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_497),
.B(n_344),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_412),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_482),
.B(n_208),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_427),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_428),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_506),
.B(n_345),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_482),
.B(n_238),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_465),
.B(n_366),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_465),
.B(n_209),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_428),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_498),
.B(n_350),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_412),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_429),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_443),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_429),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_477),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_434),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_511),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_449),
.B(n_224),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_434),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_436),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_450),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_408),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_415),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_451),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_438),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_415),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_484),
.B(n_211),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_446),
.B(n_259),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_416),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_438),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_416),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_418),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_411),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_418),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_439),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_502),
.B(n_353),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_420),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_439),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_420),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_424),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_440),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_440),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_424),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_407),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_447),
.B(n_354),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_484),
.B(n_211),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_487),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_425),
.Y(n_572)
);

AND2x6_ASAP7_75t_L g573 ( 
.A(n_425),
.B(n_228),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_451),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_419),
.A2(n_360),
.B1(n_272),
.B2(n_400),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_485),
.B(n_238),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_447),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_452),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_452),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_454),
.B(n_358),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_454),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_413),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_485),
.B(n_254),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_455),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_455),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_458),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_458),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_460),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_460),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_474),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_474),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_SL g593 ( 
.A(n_510),
.B(n_256),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_480),
.B(n_237),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_478),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_478),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_479),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_417),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_479),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_514),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_524),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_594),
.B(n_422),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_523),
.B(n_423),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_524),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_573),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_548),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_524),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_514),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_534),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_531),
.B(n_511),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_534),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_523),
.B(n_430),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_514),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_594),
.B(n_432),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_531),
.B(n_254),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_548),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_522),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_536),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_534),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_516),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_589),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_522),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_552),
.B(n_442),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_522),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_552),
.B(n_444),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_515),
.A2(n_348),
.B1(n_256),
.B2(n_337),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_546),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_589),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_589),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_546),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_548),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_515),
.A2(n_274),
.B1(n_306),
.B2(n_300),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_584),
.B(n_459),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_584),
.B(n_471),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_528),
.B(n_445),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_545),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_519),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_528),
.B(n_448),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_519),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_557),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_516),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_551),
.B(n_509),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_546),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_533),
.A2(n_348),
.B1(n_388),
.B2(n_337),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_574),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_533),
.B(n_453),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_556),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_560),
.A2(n_402),
.B1(n_388),
.B2(n_463),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_571),
.B(n_456),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_550),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_556),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_SL g652 ( 
.A(n_582),
.B(n_406),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_519),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_573),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_556),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_519),
.Y(n_656)
);

AND2x6_ASAP7_75t_L g657 ( 
.A(n_564),
.B(n_380),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_558),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_574),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_558),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_558),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_520),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_516),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_560),
.B(n_457),
.Y(n_664)
);

AND2x6_ASAP7_75t_L g665 ( 
.A(n_564),
.B(n_380),
.Y(n_665)
);

INVxp33_ASAP7_75t_L g666 ( 
.A(n_568),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_561),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_516),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_517),
.B(n_461),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_571),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_516),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_520),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_593),
.A2(n_402),
.B1(n_470),
.B2(n_241),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_561),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_561),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_593),
.A2(n_241),
.B1(n_243),
.B2(n_221),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_520),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_551),
.B(n_509),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_598),
.B(n_462),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_598),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_550),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_530),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_520),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_569),
.B(n_468),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_567),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_569),
.B(n_469),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_530),
.A2(n_271),
.B1(n_273),
.B2(n_243),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_553),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_530),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_553),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_567),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_538),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_567),
.Y(n_693)
);

INVx6_ASAP7_75t_L g694 ( 
.A(n_513),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_516),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_516),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_580),
.B(n_473),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_553),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_553),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_564),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_598),
.B(n_476),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_541),
.B(n_483),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_522),
.B(n_214),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_555),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_538),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_522),
.B(n_214),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_580),
.B(n_488),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_555),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_564),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_555),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_564),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_555),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_541),
.B(n_491),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_550),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_572),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_536),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_572),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_513),
.B(n_496),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_572),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_572),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_579),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_516),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_536),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_537),
.Y(n_724)
);

AOI21x1_ASAP7_75t_L g725 ( 
.A1(n_512),
.A2(n_481),
.B(n_231),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_579),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_537),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_579),
.Y(n_728)
);

INVx5_ASAP7_75t_L g729 ( 
.A(n_573),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_550),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_544),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_537),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_541),
.B(n_499),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_537),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_SL g735 ( 
.A(n_568),
.B(n_464),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_579),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_544),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_586),
.Y(n_738)
);

NOR2x1p5_ASAP7_75t_L g739 ( 
.A(n_551),
.B(n_271),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_513),
.B(n_501),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_570),
.B(n_220),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_570),
.B(n_220),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_550),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_575),
.B(n_505),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_513),
.B(n_508),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_512),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_570),
.B(n_507),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_575),
.B(n_466),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_518),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_576),
.B(n_467),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_518),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_623),
.B(n_475),
.C(n_472),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_600),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_646),
.B(n_550),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_602),
.B(n_489),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_610),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_610),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_640),
.Y(n_758)
);

INVx8_ASAP7_75t_L g759 ( 
.A(n_615),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_684),
.B(n_513),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_686),
.B(n_550),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_600),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_600),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_697),
.B(n_550),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_617),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_606),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_608),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_707),
.A2(n_495),
.B1(n_500),
.B2(n_494),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_682),
.A2(n_492),
.B(n_481),
.C(n_576),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_664),
.B(n_563),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_670),
.B(n_421),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_645),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_617),
.B(n_563),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_617),
.B(n_563),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_615),
.B(n_228),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_603),
.B(n_563),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_608),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_622),
.B(n_563),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_612),
.B(n_563),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_622),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_608),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_613),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_622),
.B(n_563),
.Y(n_783)
);

BUFx6f_ASAP7_75t_SL g784 ( 
.A(n_692),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_624),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_633),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_624),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_624),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_682),
.B(n_563),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_635),
.B(n_540),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_724),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_614),
.B(n_503),
.Y(n_792)
);

NOR2x1p5_ASAP7_75t_L g793 ( 
.A(n_633),
.B(n_233),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_638),
.B(n_504),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_613),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_689),
.B(n_228),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_670),
.B(n_606),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_SL g798 ( 
.A1(n_680),
.A2(n_433),
.B1(n_435),
.B2(n_431),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_740),
.B(n_540),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_689),
.B(n_437),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_669),
.B(n_540),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_634),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_615),
.A2(n_525),
.B1(n_529),
.B2(n_576),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_616),
.B(n_544),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_631),
.B(n_228),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_634),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_645),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_724),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_631),
.B(n_228),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_727),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_741),
.B(n_540),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_615),
.A2(n_525),
.B1(n_529),
.B2(n_576),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_659),
.B(n_262),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_666),
.B(n_403),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_702),
.B(n_252),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_727),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_718),
.B(n_540),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_613),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_741),
.B(n_525),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_713),
.B(n_305),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_741),
.B(n_525),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_733),
.B(n_284),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_659),
.B(n_288),
.Y(n_823)
);

NOR2xp67_ASAP7_75t_L g824 ( 
.A(n_745),
.B(n_521),
.Y(n_824)
);

O2A1O1Ixp5_ASAP7_75t_L g825 ( 
.A1(n_703),
.A2(n_583),
.B(n_576),
.C(n_525),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_703),
.B(n_294),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_732),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_734),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_746),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_732),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_741),
.B(n_703),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_636),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_703),
.B(n_529),
.Y(n_833)
);

BUFx5_ASAP7_75t_L g834 ( 
.A(n_657),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_744),
.B(n_235),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_625),
.B(n_242),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_706),
.B(n_529),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_739),
.B(n_231),
.Y(n_838)
);

AND2x2_ASAP7_75t_SL g839 ( 
.A(n_626),
.B(n_395),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_746),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_739),
.Y(n_841)
);

O2A1O1Ixp5_ASAP7_75t_L g842 ( 
.A1(n_706),
.A2(n_709),
.B(n_711),
.C(n_700),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_642),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_SL g844 ( 
.A(n_632),
.B(n_250),
.C(n_246),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_692),
.B(n_288),
.Y(n_845)
);

INVxp33_ASAP7_75t_SL g846 ( 
.A(n_652),
.Y(n_846)
);

INVx8_ASAP7_75t_L g847 ( 
.A(n_615),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_749),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_706),
.B(n_294),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_700),
.B(n_294),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_709),
.B(n_294),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_711),
.B(n_294),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_642),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_678),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_615),
.A2(n_750),
.B1(n_742),
.B2(n_649),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_615),
.A2(n_583),
.B1(n_395),
.B2(n_234),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_749),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_751),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_679),
.B(n_266),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_751),
.B(n_583),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_678),
.B(n_583),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_692),
.B(n_583),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_701),
.B(n_279),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_748),
.B(n_286),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_605),
.B(n_329),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_747),
.B(n_521),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_747),
.B(n_526),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_605),
.B(n_329),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_621),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_618),
.B(n_291),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_632),
.B(n_692),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_694),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_621),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_734),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_L g875 ( 
.A(n_657),
.B(n_329),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_734),
.B(n_526),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_742),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_742),
.B(n_694),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_605),
.B(n_329),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_605),
.B(n_329),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_605),
.B(n_368),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_742),
.B(n_527),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_605),
.B(n_371),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_628),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_601),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_742),
.B(n_527),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_694),
.B(n_532),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_735),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_SL g889 ( 
.A(n_705),
.B(n_259),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_629),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_694),
.B(n_532),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_663),
.B(n_535),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_657),
.A2(n_378),
.B1(n_387),
.B2(n_376),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_663),
.B(n_535),
.Y(n_894)
);

INVx3_ASAP7_75t_R g895 ( 
.A(n_716),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_629),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_663),
.B(n_539),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_R g898 ( 
.A(n_723),
.B(n_293),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_654),
.B(n_729),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_705),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_663),
.B(n_539),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_653),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_668),
.B(n_542),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_668),
.B(n_542),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_668),
.B(n_543),
.Y(n_905)
);

NOR3xp33_ASAP7_75t_L g906 ( 
.A(n_731),
.B(n_304),
.C(n_299),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_620),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_668),
.B(n_543),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_671),
.B(n_547),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_648),
.A2(n_392),
.B(n_283),
.C(n_289),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_601),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_653),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_705),
.B(n_309),
.Y(n_913)
);

INVxp67_ASAP7_75t_SL g914 ( 
.A(n_620),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_705),
.B(n_486),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_654),
.B(n_234),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_653),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_656),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_854),
.B(n_644),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_872),
.A2(n_681),
.B(n_650),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_854),
.B(n_604),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_872),
.A2(n_681),
.B(n_650),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_843),
.B(n_853),
.Y(n_923)
);

AO21x1_ASAP7_75t_L g924 ( 
.A1(n_796),
.A2(n_764),
.B(n_761),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_842),
.A2(n_607),
.B(n_604),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_828),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_915),
.B(n_737),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_872),
.B(n_654),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_811),
.A2(n_681),
.B(n_650),
.Y(n_929)
);

AO21x1_ASAP7_75t_L g930 ( 
.A1(n_796),
.A2(n_282),
.B(n_263),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_815),
.A2(n_282),
.B(n_298),
.C(n_263),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_760),
.B(n_609),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_829),
.B(n_840),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_828),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_825),
.A2(n_619),
.B(n_611),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_766),
.B(n_687),
.Y(n_936)
);

BUFx8_ASAP7_75t_L g937 ( 
.A(n_784),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_776),
.A2(n_681),
.B(n_650),
.Y(n_938)
);

INVx1_ASAP7_75t_SL g939 ( 
.A(n_772),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_794),
.B(n_755),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_819),
.A2(n_619),
.B(n_611),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_792),
.B(n_730),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_786),
.B(n_730),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_800),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_829),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_756),
.A2(n_757),
.B(n_867),
.C(n_866),
.Y(n_946)
);

INVx4_ASAP7_75t_L g947 ( 
.A(n_828),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_802),
.B(n_730),
.Y(n_948)
);

BUFx4f_ASAP7_75t_L g949 ( 
.A(n_807),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_806),
.B(n_766),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_779),
.A2(n_770),
.B(n_887),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_828),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_844),
.B(n_730),
.Y(n_953)
);

NOR2xp67_ASAP7_75t_SL g954 ( 
.A(n_780),
.B(n_654),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_797),
.B(n_654),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_780),
.Y(n_956)
);

AO21x1_ASAP7_75t_L g957 ( 
.A1(n_754),
.A2(n_301),
.B(n_298),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_L g958 ( 
.A(n_820),
.B(n_676),
.C(n_673),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_840),
.B(n_848),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_891),
.A2(n_714),
.B(n_641),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_821),
.A2(n_630),
.B(n_627),
.Y(n_961)
);

BUFx8_ASAP7_75t_SL g962 ( 
.A(n_758),
.Y(n_962)
);

NAND3xp33_ASAP7_75t_SL g963 ( 
.A(n_835),
.B(n_307),
.C(n_301),
.Y(n_963)
);

NOR2xp67_ASAP7_75t_L g964 ( 
.A(n_752),
.B(n_627),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_871),
.B(n_822),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_813),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_848),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_823),
.B(n_845),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_771),
.B(n_804),
.Y(n_969)
);

CKINVDCx6p67_ASAP7_75t_R g970 ( 
.A(n_784),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_857),
.Y(n_971)
);

OAI22xp33_ASAP7_75t_L g972 ( 
.A1(n_855),
.A2(n_308),
.B1(n_311),
.B2(n_307),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_857),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_831),
.A2(n_714),
.B(n_641),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_754),
.A2(n_714),
.B(n_641),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_841),
.A2(n_665),
.B1(n_657),
.B2(n_671),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_858),
.B(n_630),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_799),
.A2(n_714),
.B(n_641),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_878),
.A2(n_641),
.B(n_620),
.Y(n_979)
);

NAND2x1_ASAP7_75t_L g980 ( 
.A(n_780),
.B(n_671),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_833),
.A2(n_620),
.B(n_743),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_837),
.A2(n_620),
.B(n_743),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_858),
.B(n_861),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_790),
.B(n_643),
.Y(n_984)
);

INVxp67_ASAP7_75t_R g985 ( 
.A(n_862),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_834),
.B(n_654),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_870),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_801),
.B(n_643),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_791),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_838),
.B(n_647),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_787),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_805),
.A2(n_651),
.B(n_655),
.C(n_647),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_753),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_787),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_805),
.A2(n_809),
.B(n_886),
.C(n_882),
.Y(n_995)
);

NOR2xp67_ASAP7_75t_L g996 ( 
.A(n_768),
.B(n_651),
.Y(n_996)
);

OAI22x1_ASAP7_75t_L g997 ( 
.A1(n_864),
.A2(n_312),
.B1(n_317),
.B2(n_310),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_877),
.A2(n_311),
.B1(n_326),
.B2(n_308),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_762),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_762),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_763),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_SL g1002 ( 
.A(n_846),
.B(n_259),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_841),
.A2(n_665),
.B1(n_657),
.B2(n_695),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_914),
.A2(n_743),
.B(n_696),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_838),
.B(n_655),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_838),
.B(n_808),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_789),
.A2(n_660),
.B(n_658),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_775),
.A2(n_743),
.B(n_696),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_877),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_810),
.B(n_816),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_827),
.B(n_658),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_832),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_765),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_785),
.A2(n_396),
.B1(n_389),
.B2(n_343),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_839),
.A2(n_657),
.B1(n_665),
.B2(n_385),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_830),
.B(n_660),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_788),
.A2(n_326),
.B1(n_331),
.B2(n_335),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_SL g1018 ( 
.A(n_846),
.B(n_219),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_874),
.B(n_661),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_759),
.A2(n_396),
.B1(n_389),
.B2(n_343),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_773),
.A2(n_667),
.B(n_661),
.Y(n_1021)
);

AO21x1_ASAP7_75t_L g1022 ( 
.A1(n_809),
.A2(n_335),
.B(n_331),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_775),
.A2(n_696),
.B(n_695),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_900),
.B(n_729),
.Y(n_1024)
);

AO21x2_ASAP7_75t_L g1025 ( 
.A1(n_824),
.A2(n_725),
.B(n_674),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_773),
.A2(n_696),
.B(n_695),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_885),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_774),
.A2(n_722),
.B(n_729),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_888),
.B(n_667),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_900),
.Y(n_1030)
);

AO21x1_ASAP7_75t_L g1031 ( 
.A1(n_836),
.A2(n_341),
.B(n_338),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_860),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_889),
.B(n_674),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_839),
.B(n_675),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_911),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_793),
.B(n_338),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_774),
.A2(n_783),
.B(n_778),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_876),
.B(n_675),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_778),
.A2(n_722),
.B(n_729),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_783),
.A2(n_722),
.B(n_729),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_859),
.A2(n_372),
.B(n_367),
.C(n_341),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_869),
.B(n_685),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_869),
.B(n_873),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_884),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_910),
.A2(n_691),
.B(n_693),
.C(n_662),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_890),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_863),
.B(n_693),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_817),
.A2(n_722),
.B(n_729),
.Y(n_1048)
);

AND2x6_ASAP7_75t_L g1049 ( 
.A(n_907),
.B(n_656),
.Y(n_1049)
);

AOI21x1_ASAP7_75t_L g1050 ( 
.A1(n_881),
.A2(n_639),
.B(n_637),
.Y(n_1050)
);

BUFx8_ASAP7_75t_L g1051 ( 
.A(n_784),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_763),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_834),
.B(n_637),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_759),
.A2(n_672),
.B(n_639),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_767),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_890),
.B(n_672),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_767),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_896),
.B(n_677),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_896),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_759),
.A2(n_683),
.B(n_677),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_826),
.A2(n_662),
.B(n_656),
.C(n_683),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_759),
.A2(n_690),
.B(n_688),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_902),
.B(n_688),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_902),
.B(n_690),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_777),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_912),
.B(n_698),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_895),
.Y(n_1067)
);

AO21x1_ASAP7_75t_L g1068 ( 
.A1(n_826),
.A2(n_372),
.B(n_725),
.Y(n_1068)
);

INVx5_ASAP7_75t_L g1069 ( 
.A(n_847),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_847),
.A2(n_699),
.B(n_698),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_777),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_847),
.A2(n_704),
.B(n_699),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_814),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_781),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_834),
.B(n_704),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_913),
.B(n_708),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_881),
.A2(n_710),
.B(n_708),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_907),
.B(n_662),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_781),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_906),
.B(n_273),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_847),
.A2(n_712),
.B(n_710),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_803),
.A2(n_715),
.B(n_712),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_812),
.A2(n_717),
.B(n_715),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_907),
.B(n_283),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_899),
.A2(n_719),
.B(n_717),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_782),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_912),
.B(n_719),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_898),
.Y(n_1088)
);

AO21x1_ASAP7_75t_L g1089 ( 
.A1(n_849),
.A2(n_292),
.B(n_289),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_782),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_795),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_917),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_849),
.A2(n_720),
.B(n_547),
.C(n_549),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_917),
.B(n_720),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_883),
.A2(n_856),
.B1(n_893),
.B2(n_916),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_918),
.B(n_657),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_918),
.B(n_892),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_894),
.A2(n_738),
.B(n_728),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_899),
.A2(n_721),
.B(n_726),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_795),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_818),
.B(n_665),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_L g1102 ( 
.A1(n_850),
.A2(n_721),
.B(n_736),
.C(n_728),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_951),
.A2(n_875),
.B(n_883),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_934),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_965),
.A2(n_769),
.B(n_909),
.C(n_908),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_934),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_983),
.A2(n_875),
.B(n_897),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_984),
.A2(n_903),
.B(n_901),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_SL g1109 ( 
.A1(n_965),
.A2(n_818),
.B(n_905),
.C(n_904),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1090),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_927),
.B(n_798),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_988),
.A2(n_834),
.B(n_916),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_940),
.A2(n_852),
.B(n_851),
.C(n_850),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_940),
.A2(n_665),
.B1(n_852),
.B2(n_851),
.Y(n_1114)
);

O2A1O1Ixp5_ASAP7_75t_L g1115 ( 
.A1(n_924),
.A2(n_880),
.B(n_879),
.C(n_868),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1082),
.A2(n_665),
.B(n_865),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_978),
.A2(n_834),
.B(n_880),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1032),
.B(n_665),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_939),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_920),
.A2(n_922),
.B(n_932),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_967),
.Y(n_1121)
);

AO22x1_ASAP7_75t_L g1122 ( 
.A1(n_968),
.A2(n_321),
.B1(n_320),
.B2(n_322),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_987),
.B(n_328),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_969),
.B(n_486),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1090),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_963),
.A2(n_316),
.B(n_398),
.C(n_397),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1069),
.A2(n_834),
.B(n_865),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_966),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1069),
.A2(n_834),
.B(n_879),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_963),
.A2(n_302),
.B(n_398),
.C(n_397),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_996),
.B(n_219),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_962),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_991),
.Y(n_1133)
);

AO32x2_ASAP7_75t_L g1134 ( 
.A1(n_998),
.A2(n_302),
.A3(n_392),
.B1(n_386),
.B2(n_385),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1032),
.B(n_726),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_973),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1091),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1091),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_993),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_944),
.B(n_923),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1069),
.A2(n_868),
.B(n_728),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_931),
.A2(n_292),
.B(n_315),
.C(n_316),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1041),
.A2(n_362),
.B(n_386),
.C(n_359),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_947),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_945),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1069),
.A2(n_938),
.B(n_929),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_974),
.A2(n_738),
.B(n_736),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_991),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_923),
.B(n_490),
.Y(n_1149)
);

XOR2xp5_ASAP7_75t_L g1150 ( 
.A(n_1067),
.B(n_87),
.Y(n_1150)
);

AO21x2_ASAP7_75t_L g1151 ( 
.A1(n_941),
.A2(n_562),
.B(n_549),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_947),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1073),
.B(n_330),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_971),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_952),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_958),
.A2(n_362),
.B(n_315),
.C(n_359),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_950),
.B(n_490),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_949),
.Y(n_1158)
);

NOR3xp33_ASAP7_75t_SL g1159 ( 
.A(n_1088),
.B(n_370),
.C(n_365),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_949),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_961),
.A2(n_738),
.B(n_736),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_1012),
.B(n_333),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_972),
.A2(n_333),
.B1(n_340),
.B2(n_351),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_928),
.A2(n_726),
.B(n_595),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_991),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_972),
.A2(n_1015),
.B1(n_1047),
.B2(n_919),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1047),
.B(n_554),
.Y(n_1167)
);

CKINVDCx8_ASAP7_75t_R g1168 ( 
.A(n_1036),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1083),
.A2(n_573),
.B(n_599),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_989),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_946),
.A2(n_355),
.B(n_352),
.C(n_351),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_991),
.B(n_340),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1030),
.B(n_493),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_928),
.A2(n_595),
.B(n_590),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1027),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_1006),
.B(n_493),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_994),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1014),
.A2(n_581),
.B(n_554),
.C(n_592),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_960),
.A2(n_595),
.B(n_590),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_999),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_SL g1181 ( 
.A1(n_1034),
.A2(n_597),
.B(n_559),
.C(n_592),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_981),
.A2(n_595),
.B(n_590),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_950),
.B(n_339),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_952),
.B(n_507),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_942),
.B(n_1002),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_995),
.A2(n_401),
.B(n_347),
.C(n_356),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_937),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_R g1188 ( 
.A(n_970),
.B(n_357),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_942),
.B(n_1029),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1029),
.B(n_559),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1076),
.B(n_562),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1076),
.B(n_565),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_982),
.A2(n_595),
.B(n_590),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1018),
.B(n_363),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1015),
.A2(n_404),
.B1(n_374),
.B2(n_375),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1013),
.B(n_364),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_956),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_933),
.A2(n_590),
.B(n_591),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_SL g1199 ( 
.A(n_1031),
.B(n_399),
.C(n_377),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_964),
.B(n_295),
.Y(n_1200)
);

INVx4_ASAP7_75t_L g1201 ( 
.A(n_926),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1050),
.A2(n_597),
.B(n_565),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1009),
.B(n_92),
.Y(n_1203)
);

AO32x1_ASAP7_75t_L g1204 ( 
.A1(n_1017),
.A2(n_581),
.A3(n_566),
.B1(n_577),
.B2(n_578),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_R g1205 ( 
.A(n_926),
.B(n_381),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1097),
.B(n_566),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1035),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_959),
.A2(n_586),
.B(n_591),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_R g1209 ( 
.A(n_937),
.B(n_382),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1033),
.B(n_295),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1097),
.B(n_1010),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1051),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1095),
.A2(n_383),
.B1(n_384),
.B2(n_390),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_979),
.A2(n_586),
.B(n_591),
.Y(n_1214)
);

XOR2xp5_ASAP7_75t_L g1215 ( 
.A(n_997),
.B(n_94),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_921),
.B(n_577),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_956),
.B(n_585),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1092),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_SL g1219 ( 
.A1(n_1080),
.A2(n_394),
.B1(n_20),
.B2(n_23),
.Y(n_1219)
);

INVx6_ASAP7_75t_L g1220 ( 
.A(n_1051),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1013),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1009),
.B(n_585),
.Y(n_1222)
);

BUFx12f_ASAP7_75t_L g1223 ( 
.A(n_1036),
.Y(n_1223)
);

AO21x1_ASAP7_75t_L g1224 ( 
.A1(n_953),
.A2(n_588),
.B(n_591),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1084),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_936),
.B(n_943),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1044),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_943),
.B(n_588),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1084),
.Y(n_1229)
);

BUFx12f_ASAP7_75t_L g1230 ( 
.A(n_1080),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_948),
.B(n_587),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_948),
.B(n_19),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_990),
.A2(n_586),
.B(n_23),
.C(n_28),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1005),
.A2(n_596),
.B1(n_587),
.B2(n_30),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1046),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1038),
.A2(n_596),
.B(n_587),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1092),
.B(n_20),
.Y(n_1237)
);

INVx6_ASAP7_75t_SL g1238 ( 
.A(n_985),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1065),
.B(n_573),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1000),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1020),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1092),
.B(n_596),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1092),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_SL g1244 ( 
.A1(n_954),
.A2(n_935),
.B(n_925),
.C(n_1054),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1074),
.B(n_573),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1100),
.B(n_573),
.Y(n_1246)
);

CKINVDCx11_ASAP7_75t_R g1247 ( 
.A(n_1001),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1049),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1060),
.A2(n_596),
.B(n_587),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1052),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1059),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1037),
.B(n_596),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1055),
.Y(n_1253)
);

AO21x1_ASAP7_75t_L g1254 ( 
.A1(n_992),
.A2(n_33),
.B(n_35),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1057),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_977),
.A2(n_596),
.B1(n_587),
.B2(n_37),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_976),
.B(n_1003),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1071),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1011),
.A2(n_596),
.B1(n_587),
.B2(n_38),
.Y(n_1259)
);

CKINVDCx6p67_ASAP7_75t_R g1260 ( 
.A(n_1158),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1189),
.B(n_1211),
.Y(n_1261)
);

AO31x2_ASAP7_75t_L g1262 ( 
.A1(n_1224),
.A2(n_957),
.A3(n_1068),
.B(n_930),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_SL g1263 ( 
.A(n_1166),
.B(n_1049),
.Y(n_1263)
);

CKINVDCx11_ASAP7_75t_R g1264 ( 
.A(n_1168),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1119),
.B(n_1183),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1128),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1215),
.A2(n_1016),
.B(n_1045),
.Y(n_1267)
);

AO22x2_ASAP7_75t_L g1268 ( 
.A1(n_1166),
.A2(n_1024),
.B1(n_1075),
.B2(n_1053),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1211),
.A2(n_1019),
.B1(n_1078),
.B2(n_1053),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1186),
.A2(n_1022),
.A3(n_1089),
.B(n_975),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1113),
.A2(n_1102),
.B(n_1061),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1107),
.A2(n_1102),
.B(n_1061),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1111),
.B(n_1079),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1120),
.A2(n_1062),
.B(n_1081),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1177),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1148),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1124),
.B(n_1086),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1146),
.A2(n_1072),
.B(n_1070),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1103),
.A2(n_1075),
.B(n_986),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1254),
.A2(n_1023),
.A3(n_1008),
.B(n_1026),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1244),
.A2(n_986),
.B(n_1004),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_SL g1282 ( 
.A1(n_1185),
.A2(n_980),
.B(n_955),
.C(n_1101),
.Y(n_1282)
);

CKINVDCx11_ASAP7_75t_R g1283 ( 
.A(n_1223),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1226),
.A2(n_1096),
.B(n_1085),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1157),
.B(n_1043),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1160),
.Y(n_1286)
);

AND2x2_ASAP7_75t_SL g1287 ( 
.A(n_1194),
.B(n_1042),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1170),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1219),
.A2(n_1025),
.B1(n_1049),
.B2(n_1021),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1147),
.A2(n_1099),
.B(n_1098),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1140),
.B(n_1025),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1232),
.A2(n_1163),
.B1(n_1176),
.B2(n_1213),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1175),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1247),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1123),
.B(n_1056),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1153),
.B(n_1078),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_1104),
.B(n_1028),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1207),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1227),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1149),
.B(n_1058),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1108),
.A2(n_1048),
.B(n_1063),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1112),
.A2(n_1094),
.B(n_1064),
.Y(n_1302)
);

AO32x2_ASAP7_75t_L g1303 ( 
.A1(n_1259),
.A2(n_1093),
.A3(n_1007),
.B1(n_1049),
.B2(n_1066),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1139),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1253),
.B(n_1087),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1210),
.A2(n_1093),
.B(n_1040),
.C(n_1039),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1171),
.A2(n_1049),
.B(n_587),
.C(n_39),
.Y(n_1307)
);

NOR4xp25_ASAP7_75t_L g1308 ( 
.A(n_1241),
.B(n_33),
.C(n_36),
.D(n_41),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1229),
.B(n_41),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1259),
.A2(n_573),
.A3(n_44),
.B(n_45),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1225),
.B(n_119),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_SL g1312 ( 
.A1(n_1257),
.A2(n_1109),
.B(n_1156),
.C(n_1118),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1256),
.A2(n_573),
.A3(n_47),
.B(n_48),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1105),
.A2(n_587),
.B(n_47),
.C(n_50),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1163),
.A2(n_43),
.B1(n_53),
.B2(n_54),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1196),
.B(n_43),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1167),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1256),
.A2(n_59),
.A3(n_61),
.B(n_62),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1167),
.B(n_59),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1214),
.A2(n_144),
.B(n_206),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1117),
.A2(n_143),
.B(n_203),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1131),
.A2(n_65),
.B(n_68),
.C(n_69),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1235),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1234),
.A2(n_69),
.A3(n_71),
.B(n_72),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1133),
.B(n_150),
.Y(n_1325)
);

BUFx4f_ASAP7_75t_L g1326 ( 
.A(n_1220),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1161),
.A2(n_151),
.B(n_95),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_SL g1328 ( 
.A1(n_1118),
.A2(n_153),
.B(n_99),
.C(n_105),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1258),
.B(n_74),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1148),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_1221),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1127),
.A2(n_159),
.B(n_110),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1179),
.A2(n_160),
.B(n_112),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1190),
.B(n_74),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1251),
.B(n_115),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1199),
.A2(n_120),
.B(n_135),
.C(n_141),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1180),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1191),
.A2(n_147),
.B1(n_164),
.B2(n_171),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1148),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1129),
.A2(n_173),
.B(n_180),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1191),
.A2(n_183),
.B(n_191),
.Y(n_1341)
);

AOI222xp33_ASAP7_75t_L g1342 ( 
.A1(n_1213),
.A2(n_207),
.B1(n_1195),
.B2(n_1230),
.C1(n_1122),
.C2(n_1234),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1206),
.A2(n_1115),
.B(n_1169),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1192),
.A2(n_1206),
.B(n_1116),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1172),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1203),
.B(n_1173),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_SL g1347 ( 
.A1(n_1233),
.A2(n_1248),
.B(n_1143),
.Y(n_1347)
);

INVx4_ASAP7_75t_L g1348 ( 
.A(n_1133),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1249),
.A2(n_1193),
.B(n_1182),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1121),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1136),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1240),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1243),
.Y(n_1353)
);

OR2x6_ASAP7_75t_L g1354 ( 
.A(n_1220),
.B(n_1172),
.Y(n_1354)
);

AOI221x1_ASAP7_75t_L g1355 ( 
.A1(n_1237),
.A2(n_1192),
.B1(n_1190),
.B2(n_1228),
.C(n_1116),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1126),
.A2(n_1130),
.B(n_1142),
.C(n_1200),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1236),
.A2(n_1208),
.A3(n_1164),
.B(n_1198),
.Y(n_1357)
);

AO31x2_ASAP7_75t_L g1358 ( 
.A1(n_1217),
.A2(n_1141),
.A3(n_1216),
.B(n_1204),
.Y(n_1358)
);

AOI31xp67_ASAP7_75t_L g1359 ( 
.A1(n_1252),
.A2(n_1231),
.A3(n_1242),
.B(n_1216),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1195),
.A2(n_1222),
.B(n_1181),
.C(n_1159),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1255),
.B(n_1173),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1169),
.A2(n_1174),
.B(n_1114),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1176),
.B(n_1203),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1145),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1176),
.B(n_1135),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1154),
.B(n_1172),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1238),
.B(n_1197),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1243),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1220),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1238),
.A2(n_1184),
.B1(n_1205),
.B2(n_1250),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1162),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1165),
.B(n_1184),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1165),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1184),
.B(n_1104),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1110),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1162),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1106),
.B(n_1155),
.Y(n_1377)
);

OAI21xp33_ASAP7_75t_L g1378 ( 
.A1(n_1188),
.A2(n_1209),
.B(n_1162),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1239),
.A2(n_1246),
.B(n_1245),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1151),
.A2(n_1106),
.B(n_1155),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1178),
.A2(n_1245),
.B(n_1239),
.Y(n_1381)
);

NAND3x1_ASAP7_75t_L g1382 ( 
.A(n_1212),
.B(n_1132),
.C(n_1187),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1246),
.A2(n_1218),
.B(n_1197),
.Y(n_1383)
);

AO31x2_ASAP7_75t_L g1384 ( 
.A1(n_1204),
.A2(n_1125),
.A3(n_1137),
.B(n_1138),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1243),
.Y(n_1385)
);

AO22x2_ASAP7_75t_L g1386 ( 
.A1(n_1134),
.A2(n_1201),
.B1(n_1152),
.B2(n_1144),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1150),
.Y(n_1387)
);

AO31x2_ASAP7_75t_L g1388 ( 
.A1(n_1204),
.A2(n_1224),
.A3(n_924),
.B(n_1031),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1134),
.B(n_1201),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1134),
.A2(n_872),
.B(n_1120),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1194),
.A2(n_1002),
.B1(n_1018),
.B2(n_940),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1219),
.A2(n_965),
.B1(n_940),
.B2(n_871),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1185),
.A2(n_965),
.B(n_940),
.C(n_755),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1202),
.A2(n_1146),
.B(n_1077),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1132),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1202),
.A2(n_1146),
.B(n_1077),
.Y(n_1396)
);

AOI221x1_ASAP7_75t_L g1397 ( 
.A1(n_1186),
.A2(n_965),
.B1(n_940),
.B2(n_963),
.C(n_1166),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1120),
.A2(n_872),
.B(n_1103),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1202),
.A2(n_1146),
.B(n_1077),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1189),
.B(n_965),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1170),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_SL g1402 ( 
.A(n_1194),
.B(n_940),
.C(n_965),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1140),
.B(n_846),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1140),
.B(n_927),
.Y(n_1404)
);

AO22x2_ASAP7_75t_L g1405 ( 
.A1(n_1166),
.A2(n_844),
.B1(n_1185),
.B2(n_1163),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1158),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1148),
.Y(n_1407)
);

OR2x6_ASAP7_75t_L g1408 ( 
.A(n_1220),
.B(n_1172),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1113),
.A2(n_965),
.B(n_1189),
.Y(n_1409)
);

AOI221x1_ASAP7_75t_L g1410 ( 
.A1(n_1186),
.A2(n_965),
.B1(n_940),
.B2(n_963),
.C(n_1166),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1113),
.A2(n_965),
.B(n_1189),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1158),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1202),
.A2(n_1146),
.B(n_1077),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1119),
.Y(n_1414)
);

AOI221x1_ASAP7_75t_L g1415 ( 
.A1(n_1186),
.A2(n_965),
.B1(n_940),
.B2(n_963),
.C(n_1166),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1140),
.B(n_846),
.Y(n_1416)
);

BUFx4f_ASAP7_75t_L g1417 ( 
.A(n_1220),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1166),
.A2(n_965),
.B1(n_940),
.B2(n_871),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1148),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1202),
.A2(n_1146),
.B(n_1077),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1185),
.A2(n_965),
.B1(n_940),
.B2(n_844),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1202),
.A2(n_1146),
.B(n_1077),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1119),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1119),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1414),
.Y(n_1425)
);

NAND2x1p5_ASAP7_75t_L g1426 ( 
.A(n_1326),
.B(n_1417),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1392),
.A2(n_1402),
.B1(n_1342),
.B2(n_1391),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1400),
.B(n_1265),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1395),
.Y(n_1429)
);

CKINVDCx12_ASAP7_75t_R g1430 ( 
.A(n_1354),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1293),
.Y(n_1431)
);

INVx6_ASAP7_75t_L g1432 ( 
.A(n_1348),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1392),
.A2(n_1418),
.B1(n_1342),
.B2(n_1421),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1401),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1393),
.A2(n_1418),
.B(n_1410),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1405),
.A2(n_1411),
.B1(n_1409),
.B2(n_1292),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1283),
.Y(n_1437)
);

CKINVDCx11_ASAP7_75t_R g1438 ( 
.A(n_1264),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1405),
.A2(n_1409),
.B1(n_1411),
.B2(n_1292),
.Y(n_1439)
);

OAI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1315),
.A2(n_1397),
.B1(n_1415),
.B2(n_1261),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1276),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1288),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1304),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1317),
.A2(n_1315),
.B1(n_1316),
.B2(n_1319),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1326),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1423),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1298),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1266),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1334),
.A2(n_1287),
.B1(n_1295),
.B2(n_1263),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1330),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1263),
.A2(n_1285),
.B1(n_1378),
.B2(n_1416),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1378),
.A2(n_1403),
.B1(n_1273),
.B2(n_1365),
.Y(n_1452)
);

INVx8_ASAP7_75t_L g1453 ( 
.A(n_1354),
.Y(n_1453)
);

BUFx4f_ASAP7_75t_SL g1454 ( 
.A(n_1260),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1337),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1286),
.Y(n_1456)
);

OAI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1267),
.A2(n_1354),
.B1(n_1408),
.B2(n_1289),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1404),
.B(n_1300),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1417),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1296),
.A2(n_1376),
.B1(n_1371),
.B2(n_1346),
.Y(n_1460)
);

BUFx2_ASAP7_75t_SL g1461 ( 
.A(n_1406),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1424),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1352),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1299),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1309),
.B(n_1361),
.Y(n_1465)
);

BUFx8_ASAP7_75t_SL g1466 ( 
.A(n_1294),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1305),
.B(n_1277),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1344),
.A2(n_1338),
.B1(n_1408),
.B2(n_1268),
.Y(n_1468)
);

BUFx8_ASAP7_75t_SL g1469 ( 
.A(n_1275),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1331),
.B(n_1291),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1408),
.A2(n_1268),
.B1(n_1364),
.B2(n_1329),
.Y(n_1471)
);

NAND2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1374),
.B(n_1372),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1363),
.A2(n_1366),
.B1(n_1289),
.B2(n_1331),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1412),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1330),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1407),
.Y(n_1476)
);

OAI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1267),
.A2(n_1355),
.B1(n_1345),
.B2(n_1350),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1347),
.A2(n_1370),
.B1(n_1335),
.B2(n_1311),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_SL g1479 ( 
.A(n_1369),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1308),
.A2(n_1389),
.B1(n_1362),
.B2(n_1325),
.Y(n_1480)
);

BUFx12f_ASAP7_75t_L g1481 ( 
.A(n_1330),
.Y(n_1481)
);

OAI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1323),
.A2(n_1351),
.B1(n_1375),
.B2(n_1269),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1384),
.Y(n_1483)
);

BUFx8_ASAP7_75t_L g1484 ( 
.A(n_1339),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1384),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1339),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1322),
.A2(n_1360),
.B(n_1336),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1374),
.A2(n_1356),
.B1(n_1386),
.B2(n_1372),
.Y(n_1488)
);

BUFx10_ASAP7_75t_L g1489 ( 
.A(n_1367),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1419),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1308),
.A2(n_1362),
.B1(n_1390),
.B2(n_1341),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1343),
.A2(n_1311),
.B1(n_1386),
.B2(n_1271),
.Y(n_1492)
);

INVx6_ASAP7_75t_L g1493 ( 
.A(n_1348),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1387),
.B(n_1407),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1343),
.A2(n_1381),
.B1(n_1271),
.B2(n_1321),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1381),
.A2(n_1332),
.B1(n_1340),
.B2(n_1284),
.Y(n_1496)
);

BUFx8_ASAP7_75t_L g1497 ( 
.A(n_1419),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1385),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1353),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1324),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1419),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1324),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1324),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1314),
.B(n_1377),
.Y(n_1504)
);

BUFx2_ASAP7_75t_SL g1505 ( 
.A(n_1382),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_SL g1506 ( 
.A1(n_1318),
.A2(n_1327),
.B1(n_1272),
.B2(n_1310),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1318),
.Y(n_1507)
);

BUFx12f_ASAP7_75t_L g1508 ( 
.A(n_1353),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1297),
.A2(n_1281),
.B1(n_1373),
.B2(n_1380),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1318),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1272),
.A2(n_1297),
.B1(n_1279),
.B2(n_1302),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1368),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1307),
.A2(n_1312),
.B1(n_1373),
.B2(n_1282),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1368),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1368),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1379),
.A2(n_1333),
.B1(n_1320),
.B2(n_1301),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1328),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1310),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1310),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1313),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1313),
.Y(n_1521)
);

INVx4_ASAP7_75t_L g1522 ( 
.A(n_1383),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1280),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1359),
.Y(n_1524)
);

INVx6_ASAP7_75t_L g1525 ( 
.A(n_1306),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1280),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1303),
.A2(n_1388),
.B1(n_1270),
.B2(n_1262),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1358),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1274),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1358),
.Y(n_1530)
);

BUFx8_ASAP7_75t_SL g1531 ( 
.A(n_1388),
.Y(n_1531)
);

BUFx12f_ASAP7_75t_L g1532 ( 
.A(n_1270),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_SL g1533 ( 
.A(n_1303),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1398),
.A2(n_1349),
.B1(n_1290),
.B2(n_1422),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1270),
.Y(n_1535)
);

CKINVDCx11_ASAP7_75t_R g1536 ( 
.A(n_1262),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1394),
.A2(n_1420),
.B1(n_1413),
.B2(n_1399),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1388),
.Y(n_1538)
);

BUFx8_ASAP7_75t_L g1539 ( 
.A(n_1303),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1396),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1278),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1262),
.A2(n_940),
.B1(n_965),
.B2(n_1392),
.Y(n_1542)
);

CKINVDCx11_ASAP7_75t_R g1543 ( 
.A(n_1357),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1357),
.A2(n_965),
.B1(n_1392),
.B2(n_1402),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1293),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1392),
.A2(n_940),
.B1(n_965),
.B2(n_1418),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1293),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1395),
.Y(n_1548)
);

INVx3_ASAP7_75t_SL g1549 ( 
.A(n_1260),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1293),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1392),
.A2(n_940),
.B1(n_1402),
.B2(n_965),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1414),
.Y(n_1552)
);

INVx6_ASAP7_75t_L g1553 ( 
.A(n_1348),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1293),
.Y(n_1554)
);

CKINVDCx11_ASAP7_75t_R g1555 ( 
.A(n_1395),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1392),
.A2(n_965),
.B1(n_1402),
.B2(n_940),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1293),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1293),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1392),
.A2(n_965),
.B1(n_1402),
.B2(n_940),
.Y(n_1559)
);

INVx6_ASAP7_75t_L g1560 ( 
.A(n_1348),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1392),
.A2(n_965),
.B1(n_1402),
.B2(n_940),
.Y(n_1561)
);

OAI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1418),
.A2(n_1315),
.B1(n_965),
.B2(n_1292),
.Y(n_1562)
);

OAI21xp33_ASAP7_75t_L g1563 ( 
.A1(n_1402),
.A2(n_965),
.B(n_940),
.Y(n_1563)
);

OAI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1418),
.A2(n_1315),
.B1(n_965),
.B2(n_1292),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1392),
.A2(n_940),
.B1(n_965),
.B2(n_1418),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1293),
.Y(n_1566)
);

INVx6_ASAP7_75t_L g1567 ( 
.A(n_1348),
.Y(n_1567)
);

INVx3_ASAP7_75t_SL g1568 ( 
.A(n_1260),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1400),
.B(n_940),
.Y(n_1569)
);

CKINVDCx6p67_ASAP7_75t_R g1570 ( 
.A(n_1264),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1293),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1392),
.A2(n_940),
.B1(n_792),
.B2(n_755),
.Y(n_1572)
);

INVxp67_ASAP7_75t_SL g1573 ( 
.A(n_1344),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1392),
.A2(n_940),
.B1(n_792),
.B2(n_755),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1392),
.A2(n_965),
.B1(n_1402),
.B2(n_940),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1392),
.A2(n_940),
.B1(n_792),
.B2(n_755),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1293),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1326),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1392),
.A2(n_965),
.B1(n_940),
.B2(n_1219),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1392),
.A2(n_940),
.B1(n_1402),
.B2(n_965),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1392),
.A2(n_965),
.B1(n_1402),
.B2(n_940),
.Y(n_1581)
);

INVx4_ASAP7_75t_L g1582 ( 
.A(n_1276),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1500),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1502),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1532),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1453),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1436),
.B(n_1439),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1537),
.A2(n_1516),
.B(n_1534),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1503),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1436),
.B(n_1439),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1537),
.A2(n_1516),
.B(n_1511),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1528),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1507),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1574),
.A2(n_1433),
.B1(n_1572),
.B2(n_1576),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1522),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1442),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1470),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1453),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1435),
.B(n_1510),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1447),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1464),
.Y(n_1601)
);

OA21x2_ASAP7_75t_L g1602 ( 
.A1(n_1518),
.A2(n_1520),
.B(n_1519),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1428),
.B(n_1569),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1521),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1538),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1544),
.B(n_1492),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1531),
.Y(n_1607)
);

OAI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1546),
.A2(n_1565),
.B1(n_1562),
.B2(n_1564),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1544),
.B(n_1492),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1483),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1511),
.A2(n_1524),
.B(n_1509),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1453),
.Y(n_1612)
);

NAND2x1_ASAP7_75t_L g1613 ( 
.A(n_1525),
.B(n_1522),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1472),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1485),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1433),
.A2(n_1427),
.B1(n_1579),
.B2(n_1562),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1432),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1530),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1431),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1526),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1472),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1480),
.B(n_1471),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1527),
.Y(n_1623)
);

AOI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1542),
.A2(n_1504),
.B(n_1535),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1495),
.A2(n_1496),
.B(n_1523),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1552),
.Y(n_1626)
);

OR2x2_ASAP7_75t_SL g1627 ( 
.A(n_1525),
.B(n_1564),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1495),
.A2(n_1496),
.B(n_1573),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1434),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1529),
.B(n_1540),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1468),
.A2(n_1513),
.B(n_1488),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1545),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1533),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1541),
.B(n_1471),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1525),
.Y(n_1635)
);

AO31x2_ASAP7_75t_L g1636 ( 
.A1(n_1517),
.A2(n_1491),
.A3(n_1533),
.B(n_1506),
.Y(n_1636)
);

AO21x2_ASAP7_75t_L g1637 ( 
.A1(n_1491),
.A2(n_1440),
.B(n_1482),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1550),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1539),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1554),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1539),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1480),
.B(n_1506),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1541),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1482),
.Y(n_1644)
);

AOI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1557),
.A2(n_1571),
.B(n_1558),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1432),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1468),
.A2(n_1487),
.B(n_1449),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1543),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1547),
.Y(n_1649)
);

BUFx4f_ASAP7_75t_SL g1650 ( 
.A(n_1548),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1536),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1517),
.Y(n_1652)
);

AO21x2_ASAP7_75t_L g1653 ( 
.A1(n_1440),
.A2(n_1477),
.B(n_1457),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1566),
.B(n_1577),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1477),
.Y(n_1655)
);

INVx4_ASAP7_75t_L g1656 ( 
.A(n_1432),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1449),
.B(n_1443),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1484),
.Y(n_1658)
);

INVx6_ASAP7_75t_L g1659 ( 
.A(n_1484),
.Y(n_1659)
);

BUFx2_ASAP7_75t_R g1660 ( 
.A(n_1469),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1430),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1457),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1455),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1473),
.A2(n_1579),
.B1(n_1505),
.B2(n_1551),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1463),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1425),
.Y(n_1666)
);

AO21x2_ASAP7_75t_L g1667 ( 
.A1(n_1563),
.A2(n_1498),
.B(n_1467),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1476),
.Y(n_1668)
);

OAI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1556),
.A2(n_1575),
.B(n_1581),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1580),
.A2(n_1581),
.B1(n_1561),
.B2(n_1559),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1458),
.B(n_1556),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1446),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1512),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1451),
.A2(n_1460),
.B(n_1478),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1448),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1515),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1499),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1452),
.B(n_1451),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1514),
.Y(n_1679)
);

AO21x2_ASAP7_75t_L g1680 ( 
.A1(n_1559),
.A2(n_1575),
.B(n_1561),
.Y(n_1680)
);

OR2x6_ASAP7_75t_L g1681 ( 
.A(n_1426),
.B(n_1459),
.Y(n_1681)
);

CKINVDCx11_ASAP7_75t_R g1682 ( 
.A(n_1437),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1465),
.B(n_1452),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1475),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_SL g1685 ( 
.A1(n_1462),
.A2(n_1461),
.B1(n_1454),
.B2(n_1494),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1444),
.A2(n_1479),
.B1(n_1570),
.B2(n_1474),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1493),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1444),
.B(n_1441),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1490),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1493),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1493),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1553),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1582),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1553),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1553),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1560),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1560),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1560),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1479),
.A2(n_1489),
.B1(n_1445),
.B2(n_1578),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1426),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1567),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1567),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1567),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1501),
.B(n_1489),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1456),
.A2(n_1438),
.B1(n_1568),
.B2(n_1549),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1450),
.B(n_1486),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1549),
.A2(n_1568),
.B1(n_1454),
.B2(n_1555),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1450),
.B(n_1486),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1429),
.B(n_1497),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1497),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1481),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1508),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1466),
.Y(n_1713)
);

OR2x6_ASAP7_75t_L g1714 ( 
.A(n_1681),
.B(n_1635),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1597),
.B(n_1633),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1603),
.B(n_1683),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1626),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1683),
.B(n_1671),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_R g1719 ( 
.A(n_1682),
.B(n_1713),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1594),
.A2(n_1616),
.B1(n_1608),
.B2(n_1670),
.Y(n_1720)
);

AO32x2_ASAP7_75t_L g1721 ( 
.A1(n_1637),
.A2(n_1598),
.A3(n_1586),
.B1(n_1636),
.B2(n_1633),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1630),
.B(n_1648),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1630),
.B(n_1648),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1599),
.B(n_1596),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1614),
.B(n_1621),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1610),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1600),
.B(n_1601),
.Y(n_1727)
);

AO32x2_ASAP7_75t_L g1728 ( 
.A1(n_1637),
.A2(n_1598),
.A3(n_1586),
.B1(n_1636),
.B2(n_1617),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1650),
.Y(n_1729)
);

OAI211xp5_ASAP7_75t_L g1730 ( 
.A1(n_1594),
.A2(n_1664),
.B(n_1669),
.C(n_1670),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1666),
.B(n_1704),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1654),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1668),
.B(n_1639),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1614),
.B(n_1621),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1672),
.B(n_1675),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1591),
.A2(n_1588),
.B(n_1625),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1610),
.Y(n_1737)
);

OAI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1647),
.A2(n_1674),
.B(n_1686),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1661),
.B(n_1709),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1619),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1647),
.A2(n_1674),
.B(n_1631),
.Y(n_1741)
);

NOR4xp25_ASAP7_75t_SL g1742 ( 
.A(n_1607),
.B(n_1635),
.C(n_1662),
.D(n_1585),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1627),
.A2(n_1678),
.B1(n_1607),
.B2(n_1699),
.Y(n_1743)
);

AO32x2_ASAP7_75t_L g1744 ( 
.A1(n_1637),
.A2(n_1636),
.A3(n_1687),
.B1(n_1617),
.B2(n_1701),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1631),
.A2(n_1678),
.B(n_1628),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1713),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1709),
.B(n_1660),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1668),
.B(n_1639),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1614),
.B(n_1621),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1585),
.B(n_1681),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1629),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1641),
.B(n_1651),
.Y(n_1752)
);

AO22x2_ASAP7_75t_L g1753 ( 
.A1(n_1642),
.A2(n_1655),
.B1(n_1622),
.B2(n_1620),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1641),
.B(n_1651),
.Y(n_1754)
);

CKINVDCx6p67_ASAP7_75t_R g1755 ( 
.A(n_1658),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1657),
.B(n_1688),
.Y(n_1756)
);

NAND3xp33_ASAP7_75t_L g1757 ( 
.A(n_1655),
.B(n_1587),
.C(n_1590),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1657),
.B(n_1688),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1627),
.A2(n_1685),
.B1(n_1659),
.B2(n_1642),
.Y(n_1759)
);

OA21x2_ASAP7_75t_L g1760 ( 
.A1(n_1591),
.A2(n_1588),
.B(n_1625),
.Y(n_1760)
);

OAI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1628),
.A2(n_1644),
.B(n_1611),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1606),
.B(n_1609),
.Y(n_1762)
);

OR2x6_ASAP7_75t_L g1763 ( 
.A(n_1681),
.B(n_1613),
.Y(n_1763)
);

OA21x2_ASAP7_75t_L g1764 ( 
.A1(n_1611),
.A2(n_1583),
.B(n_1584),
.Y(n_1764)
);

INVx2_ASAP7_75t_SL g1765 ( 
.A(n_1659),
.Y(n_1765)
);

NAND2x1p5_ASAP7_75t_L g1766 ( 
.A(n_1656),
.B(n_1703),
.Y(n_1766)
);

A2O1A1Ixp33_ASAP7_75t_L g1767 ( 
.A1(n_1609),
.A2(n_1644),
.B(n_1623),
.C(n_1634),
.Y(n_1767)
);

A2O1A1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1623),
.A2(n_1634),
.B(n_1613),
.C(n_1658),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1667),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1654),
.B(n_1632),
.Y(n_1770)
);

O2A1O1Ixp33_ASAP7_75t_SL g1771 ( 
.A1(n_1710),
.A2(n_1646),
.B(n_1687),
.C(n_1701),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1659),
.A2(n_1705),
.B1(n_1707),
.B2(n_1681),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1695),
.B(n_1696),
.Y(n_1773)
);

OA21x2_ASAP7_75t_L g1774 ( 
.A1(n_1584),
.A2(n_1589),
.B(n_1593),
.Y(n_1774)
);

BUFx4f_ASAP7_75t_SL g1775 ( 
.A(n_1658),
.Y(n_1775)
);

OA21x2_ASAP7_75t_L g1776 ( 
.A1(n_1589),
.A2(n_1593),
.B(n_1604),
.Y(n_1776)
);

INVxp67_ASAP7_75t_SL g1777 ( 
.A(n_1643),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1711),
.B(n_1712),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1680),
.A2(n_1653),
.B1(n_1659),
.B2(n_1634),
.Y(n_1779)
);

NOR2x1_ASAP7_75t_SL g1780 ( 
.A(n_1653),
.B(n_1667),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1638),
.B(n_1640),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1710),
.Y(n_1782)
);

NAND2x1p5_ASAP7_75t_L g1783 ( 
.A(n_1656),
.B(n_1703),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1680),
.A2(n_1634),
.B1(n_1700),
.B2(n_1654),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1695),
.B(n_1696),
.Y(n_1785)
);

AOI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1673),
.A2(n_1676),
.B1(n_1665),
.B2(n_1663),
.C(n_1604),
.Y(n_1786)
);

OAI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1624),
.A2(n_1693),
.B(n_1645),
.Y(n_1787)
);

BUFx8_ASAP7_75t_L g1788 ( 
.A(n_1711),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1689),
.B(n_1684),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1774),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1759),
.B(n_1612),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1718),
.B(n_1676),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1774),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1726),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1716),
.B(n_1712),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1732),
.B(n_1595),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1756),
.B(n_1636),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1776),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1776),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1758),
.B(n_1636),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1735),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1784),
.B(n_1615),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1784),
.B(n_1615),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1762),
.B(n_1643),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1724),
.B(n_1602),
.Y(n_1805)
);

AOI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1730),
.A2(n_1679),
.B1(n_1663),
.B2(n_1649),
.C(n_1677),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1779),
.B(n_1602),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1737),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1764),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1779),
.B(n_1753),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1720),
.A2(n_1700),
.B1(n_1612),
.B2(n_1691),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1770),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1753),
.B(n_1602),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1715),
.B(n_1602),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1745),
.B(n_1618),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1773),
.Y(n_1816)
);

INVx4_ASAP7_75t_L g1817 ( 
.A(n_1763),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1720),
.A2(n_1700),
.B1(n_1612),
.B2(n_1696),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1739),
.B(n_1700),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1767),
.A2(n_1612),
.B1(n_1690),
.B2(n_1691),
.Y(n_1820)
);

INVxp67_ASAP7_75t_L g1821 ( 
.A(n_1717),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1744),
.Y(n_1822)
);

NOR2x1_ASAP7_75t_L g1823 ( 
.A(n_1787),
.B(n_1595),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1738),
.A2(n_1612),
.B1(n_1702),
.B2(n_1652),
.Y(n_1824)
);

INVxp67_ASAP7_75t_L g1825 ( 
.A(n_1789),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1733),
.B(n_1748),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1757),
.A2(n_1697),
.B1(n_1692),
.B2(n_1694),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1761),
.B(n_1592),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1769),
.B(n_1592),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1721),
.B(n_1605),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1721),
.B(n_1605),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1785),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1727),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_1794),
.Y(n_1834)
);

OAI31xp33_ASAP7_75t_L g1835 ( 
.A1(n_1791),
.A2(n_1743),
.A3(n_1757),
.B(n_1772),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1805),
.B(n_1777),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1808),
.Y(n_1837)
);

INVx4_ASAP7_75t_L g1838 ( 
.A(n_1817),
.Y(n_1838)
);

NAND3xp33_ASAP7_75t_L g1839 ( 
.A(n_1806),
.B(n_1741),
.C(n_1742),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1801),
.B(n_1719),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1810),
.B(n_1752),
.Y(n_1841)
);

OAI31xp33_ASAP7_75t_L g1842 ( 
.A1(n_1820),
.A2(n_1768),
.A3(n_1722),
.B(n_1723),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1810),
.B(n_1754),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1814),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1797),
.B(n_1721),
.Y(n_1845)
);

BUFx3_ASAP7_75t_L g1846 ( 
.A(n_1796),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1814),
.B(n_1736),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1817),
.B(n_1750),
.Y(n_1848)
);

AOI221xp5_ASAP7_75t_L g1849 ( 
.A1(n_1822),
.A2(n_1778),
.B1(n_1731),
.B2(n_1786),
.C(n_1747),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1790),
.Y(n_1850)
);

OAI31xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1811),
.A2(n_1749),
.A3(n_1734),
.B(n_1725),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1808),
.Y(n_1852)
);

INVx4_ASAP7_75t_L g1853 ( 
.A(n_1817),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1797),
.B(n_1744),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1812),
.B(n_1736),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_R g1856 ( 
.A(n_1819),
.B(n_1746),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1800),
.B(n_1744),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1795),
.A2(n_1714),
.B1(n_1749),
.B2(n_1734),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1802),
.Y(n_1859)
);

BUFx3_ASAP7_75t_L g1860 ( 
.A(n_1796),
.Y(n_1860)
);

AOI33xp33_ASAP7_75t_L g1861 ( 
.A1(n_1807),
.A2(n_1781),
.A3(n_1771),
.B1(n_1765),
.B2(n_1740),
.B3(n_1751),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1800),
.B(n_1728),
.Y(n_1862)
);

NOR3xp33_ASAP7_75t_SL g1863 ( 
.A(n_1827),
.B(n_1782),
.C(n_1697),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1790),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1813),
.B(n_1760),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1793),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1793),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1809),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1815),
.B(n_1780),
.Y(n_1869)
);

INVxp67_ASAP7_75t_SL g1870 ( 
.A(n_1798),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1824),
.A2(n_1714),
.B1(n_1725),
.B2(n_1788),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1815),
.B(n_1792),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1813),
.B(n_1760),
.Y(n_1873)
);

OAI221xp5_ASAP7_75t_SL g1874 ( 
.A1(n_1818),
.A2(n_1755),
.B1(n_1763),
.B2(n_1729),
.C(n_1719),
.Y(n_1874)
);

HB1xp67_ASAP7_75t_L g1875 ( 
.A(n_1802),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1803),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1816),
.B(n_1832),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1822),
.A2(n_1775),
.B1(n_1652),
.B2(n_1624),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1833),
.B(n_1780),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1821),
.A2(n_1652),
.B1(n_1783),
.B2(n_1766),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1816),
.B(n_1728),
.Y(n_1881)
);

BUFx3_ASAP7_75t_L g1882 ( 
.A(n_1796),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1850),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1881),
.B(n_1830),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1850),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1850),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1849),
.B(n_1817),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1847),
.B(n_1799),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1836),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1881),
.B(n_1830),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1862),
.B(n_1831),
.Y(n_1891)
);

INVx2_ASAP7_75t_SL g1892 ( 
.A(n_1864),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1834),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1862),
.B(n_1831),
.Y(n_1894)
);

INVx4_ASAP7_75t_L g1895 ( 
.A(n_1838),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1864),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1868),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1837),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1837),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1852),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1854),
.B(n_1803),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1866),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1849),
.B(n_1823),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1857),
.B(n_1823),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1857),
.B(n_1826),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1845),
.B(n_1826),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1845),
.B(n_1804),
.Y(n_1907)
);

BUFx2_ASAP7_75t_L g1908 ( 
.A(n_1870),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1866),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1852),
.Y(n_1910)
);

BUFx2_ASAP7_75t_L g1911 ( 
.A(n_1870),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1855),
.B(n_1829),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1859),
.B(n_1875),
.Y(n_1913)
);

NOR2xp67_ASAP7_75t_L g1914 ( 
.A(n_1839),
.B(n_1809),
.Y(n_1914)
);

BUFx3_ASAP7_75t_L g1915 ( 
.A(n_1838),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1872),
.B(n_1804),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1866),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1876),
.B(n_1825),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1867),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1844),
.B(n_1809),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1867),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1835),
.A2(n_1839),
.B1(n_1863),
.B2(n_1874),
.C(n_1878),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1872),
.B(n_1833),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1841),
.B(n_1809),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1841),
.B(n_1843),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1855),
.B(n_1828),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1898),
.Y(n_1927)
);

INVxp67_ASAP7_75t_SL g1928 ( 
.A(n_1914),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1898),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1908),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1914),
.B(n_1838),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1899),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1908),
.Y(n_1933)
);

INVx2_ASAP7_75t_SL g1934 ( 
.A(n_1915),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1901),
.B(n_1846),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1901),
.B(n_1846),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_R g1937 ( 
.A(n_1915),
.B(n_1788),
.Y(n_1937)
);

NAND2xp33_ASAP7_75t_SL g1938 ( 
.A(n_1903),
.B(n_1863),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1913),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1903),
.B(n_1861),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1901),
.B(n_1860),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1915),
.B(n_1838),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1908),
.Y(n_1943)
);

OR2x6_ASAP7_75t_L g1944 ( 
.A(n_1895),
.B(n_1853),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1889),
.B(n_1879),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1911),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1899),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1900),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1925),
.B(n_1860),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1900),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1925),
.B(n_1860),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1910),
.Y(n_1952)
);

INVxp67_ASAP7_75t_L g1953 ( 
.A(n_1887),
.Y(n_1953)
);

INVx1_ASAP7_75t_SL g1954 ( 
.A(n_1915),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1913),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1889),
.B(n_1879),
.Y(n_1956)
);

NAND3xp33_ASAP7_75t_SL g1957 ( 
.A(n_1922),
.B(n_1835),
.C(n_1842),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1925),
.B(n_1882),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1904),
.B(n_1882),
.Y(n_1959)
);

NOR2x1_ASAP7_75t_SL g1960 ( 
.A(n_1913),
.B(n_1853),
.Y(n_1960)
);

NOR2x1_ASAP7_75t_L g1961 ( 
.A(n_1895),
.B(n_1840),
.Y(n_1961)
);

NAND2x1_ASAP7_75t_L g1962 ( 
.A(n_1911),
.B(n_1904),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1926),
.B(n_1865),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1904),
.B(n_1882),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1911),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1910),
.Y(n_1966)
);

AOI221xp5_ASAP7_75t_L g1967 ( 
.A1(n_1922),
.A2(n_1869),
.B1(n_1878),
.B2(n_1874),
.C(n_1842),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1885),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1885),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1885),
.Y(n_1970)
);

AOI32xp33_ASAP7_75t_L g1971 ( 
.A1(n_1887),
.A2(n_1843),
.A3(n_1869),
.B1(n_1848),
.B2(n_1853),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1892),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1906),
.B(n_1877),
.Y(n_1973)
);

NAND3xp33_ASAP7_75t_L g1974 ( 
.A(n_1895),
.B(n_1871),
.C(n_1851),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1906),
.B(n_1877),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1886),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1940),
.B(n_1891),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1928),
.B(n_1891),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1957),
.A2(n_1895),
.B1(n_1848),
.B2(n_1853),
.Y(n_1979)
);

NOR3xp33_ASAP7_75t_L g1980 ( 
.A(n_1938),
.B(n_1895),
.C(n_1880),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1927),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1935),
.B(n_1891),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1927),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1953),
.B(n_1894),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1935),
.B(n_1894),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1939),
.B(n_1894),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1955),
.B(n_1945),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1961),
.B(n_1916),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1954),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1967),
.B(n_1856),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1936),
.B(n_1884),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1929),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1960),
.B(n_1884),
.Y(n_1993)
);

AOI221xp5_ASAP7_75t_L g1994 ( 
.A1(n_1974),
.A2(n_1926),
.B1(n_1890),
.B2(n_1884),
.C(n_1865),
.Y(n_1994)
);

NAND4xp75_ASAP7_75t_L g1995 ( 
.A(n_1934),
.B(n_1690),
.C(n_1698),
.D(n_1692),
.Y(n_1995)
);

AND2x4_ASAP7_75t_L g1996 ( 
.A(n_1960),
.B(n_1892),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1929),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1972),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1942),
.B(n_1916),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1931),
.B(n_1890),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1930),
.Y(n_2001)
);

INVxp67_ASAP7_75t_SL g2002 ( 
.A(n_1962),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1972),
.Y(n_2003)
);

INVx2_ASAP7_75t_SL g2004 ( 
.A(n_1962),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1932),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1936),
.B(n_1890),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1941),
.B(n_1905),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1941),
.B(n_1905),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1930),
.B(n_1906),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1933),
.B(n_1905),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1933),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1943),
.B(n_1907),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1949),
.B(n_1924),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1945),
.B(n_1926),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1943),
.B(n_1907),
.Y(n_2015)
);

INVx1_ASAP7_75t_SL g2016 ( 
.A(n_1931),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1946),
.B(n_1907),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_2001),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2001),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1981),
.Y(n_2020)
);

NAND2x1_ASAP7_75t_L g2021 ( 
.A(n_1996),
.B(n_1931),
.Y(n_2021)
);

AOI221x1_ASAP7_75t_SL g2022 ( 
.A1(n_1977),
.A2(n_1931),
.B1(n_1946),
.B2(n_1965),
.C(n_1932),
.Y(n_2022)
);

AOI221xp5_ASAP7_75t_L g2023 ( 
.A1(n_1994),
.A2(n_1971),
.B1(n_1965),
.B2(n_1934),
.C(n_1942),
.Y(n_2023)
);

AOI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1990),
.A2(n_1942),
.B1(n_1944),
.B2(n_1959),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1981),
.Y(n_2025)
);

AOI322xp5_ASAP7_75t_L g2026 ( 
.A1(n_1994),
.A2(n_1975),
.A3(n_1973),
.B1(n_1951),
.B2(n_1958),
.C1(n_1949),
.C2(n_1959),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_2004),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1983),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1983),
.Y(n_2029)
);

OAI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1980),
.A2(n_1942),
.B(n_1944),
.Y(n_2030)
);

INVx1_ASAP7_75t_SL g2031 ( 
.A(n_1989),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1992),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1978),
.B(n_1964),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_2004),
.B(n_1944),
.Y(n_2034)
);

AOI21xp33_ASAP7_75t_L g2035 ( 
.A1(n_1989),
.A2(n_1944),
.B(n_1956),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1992),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_1984),
.B(n_1956),
.Y(n_2037)
);

HB1xp67_ASAP7_75t_L g2038 ( 
.A(n_1978),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1977),
.B(n_1973),
.Y(n_2039)
);

INVx1_ASAP7_75t_SL g2040 ( 
.A(n_1978),
.Y(n_2040)
);

INVxp67_ASAP7_75t_L g2041 ( 
.A(n_2002),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1988),
.B(n_1975),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1997),
.Y(n_2043)
);

AOI21xp33_ASAP7_75t_L g2044 ( 
.A1(n_1979),
.A2(n_1944),
.B(n_1947),
.Y(n_2044)
);

INVx1_ASAP7_75t_SL g2045 ( 
.A(n_2016),
.Y(n_2045)
);

AO22x1_ASAP7_75t_L g2046 ( 
.A1(n_2002),
.A2(n_1964),
.B1(n_1951),
.B2(n_1958),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_1980),
.A2(n_1880),
.B1(n_1848),
.B2(n_1924),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2038),
.Y(n_2048)
);

NAND2x1p5_ASAP7_75t_L g2049 ( 
.A(n_2031),
.B(n_2016),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_2038),
.B(n_1993),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2018),
.Y(n_2051)
);

A2O1A1Ixp33_ASAP7_75t_L g2052 ( 
.A1(n_2022),
.A2(n_1993),
.B(n_2004),
.C(n_1984),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2019),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2040),
.Y(n_2054)
);

NOR3xp33_ASAP7_75t_L g2055 ( 
.A(n_2030),
.B(n_2011),
.C(n_1987),
.Y(n_2055)
);

OAI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_2023),
.A2(n_1986),
.B1(n_1993),
.B2(n_1987),
.Y(n_2056)
);

AOI22xp5_ASAP7_75t_SL g2057 ( 
.A1(n_2041),
.A2(n_1996),
.B1(n_2000),
.B2(n_2011),
.Y(n_2057)
);

OAI221xp5_ASAP7_75t_L g2058 ( 
.A1(n_2024),
.A2(n_1999),
.B1(n_1986),
.B2(n_2010),
.C(n_2009),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2047),
.A2(n_1995),
.B1(n_2000),
.B2(n_1985),
.Y(n_2059)
);

AOI221xp5_ASAP7_75t_L g2060 ( 
.A1(n_2035),
.A2(n_2000),
.B1(n_2009),
.B2(n_2010),
.C(n_1997),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2020),
.Y(n_2061)
);

INVx1_ASAP7_75t_SL g2062 ( 
.A(n_2045),
.Y(n_2062)
);

OAI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_2021),
.A2(n_2017),
.B1(n_2015),
.B2(n_2012),
.Y(n_2063)
);

NAND2xp33_ASAP7_75t_L g2064 ( 
.A(n_2033),
.B(n_1937),
.Y(n_2064)
);

AOI21xp33_ASAP7_75t_L g2065 ( 
.A1(n_2044),
.A2(n_2011),
.B(n_2014),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2033),
.B(n_1982),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2025),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2028),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2029),
.Y(n_2069)
);

AOI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_2042),
.A2(n_1982),
.B1(n_1985),
.B2(n_1991),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2039),
.B(n_1991),
.Y(n_2071)
);

AOI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_2056),
.A2(n_2046),
.B1(n_2034),
.B2(n_2041),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2048),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2062),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_2062),
.B(n_2026),
.Y(n_2075)
);

AOI211x1_ASAP7_75t_L g2076 ( 
.A1(n_2063),
.A2(n_2012),
.B(n_2015),
.C(n_2017),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2050),
.Y(n_2077)
);

AOI32xp33_ASAP7_75t_L g2078 ( 
.A1(n_2055),
.A2(n_2034),
.A3(n_1996),
.B1(n_2006),
.B2(n_2043),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2050),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2049),
.Y(n_2080)
);

O2A1O1Ixp33_ASAP7_75t_L g2081 ( 
.A1(n_2049),
.A2(n_2052),
.B(n_2065),
.C(n_2059),
.Y(n_2081)
);

NAND2xp33_ASAP7_75t_L g2082 ( 
.A(n_2066),
.B(n_2037),
.Y(n_2082)
);

OA22x2_ASAP7_75t_SL g2083 ( 
.A1(n_2054),
.A2(n_2027),
.B1(n_2032),
.B2(n_2036),
.Y(n_2083)
);

AOI222xp33_ASAP7_75t_L g2084 ( 
.A1(n_2060),
.A2(n_1996),
.B1(n_2034),
.B2(n_2027),
.C1(n_2005),
.C2(n_2006),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_2071),
.B(n_2014),
.Y(n_2085)
);

OAI22xp33_ASAP7_75t_SL g2086 ( 
.A1(n_2058),
.A2(n_2005),
.B1(n_2003),
.B2(n_1998),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_2051),
.Y(n_2087)
);

INVxp67_ASAP7_75t_L g2088 ( 
.A(n_2080),
.Y(n_2088)
);

NAND4xp25_ASAP7_75t_L g2089 ( 
.A(n_2081),
.B(n_2053),
.C(n_2070),
.D(n_2057),
.Y(n_2089)
);

NAND5xp2_ASAP7_75t_L g2090 ( 
.A(n_2084),
.B(n_2069),
.C(n_2068),
.D(n_2067),
.E(n_2061),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2074),
.Y(n_2091)
);

AOI321xp33_ASAP7_75t_L g2092 ( 
.A1(n_2075),
.A2(n_2064),
.A3(n_2003),
.B1(n_1998),
.B2(n_2007),
.C(n_2008),
.Y(n_2092)
);

NAND2x1p5_ASAP7_75t_L g2093 ( 
.A(n_2077),
.B(n_2007),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_2085),
.B(n_2008),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2079),
.Y(n_2095)
);

AND4x1_ASAP7_75t_L g2096 ( 
.A(n_2072),
.B(n_1851),
.C(n_2013),
.D(n_1858),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2078),
.B(n_2013),
.Y(n_2097)
);

OAI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2076),
.A2(n_1995),
.B1(n_1998),
.B2(n_2003),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2073),
.B(n_1947),
.Y(n_2099)
);

AOI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_2086),
.A2(n_1966),
.B(n_1952),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2087),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2093),
.B(n_2082),
.Y(n_2102)
);

AOI21xp5_ASAP7_75t_L g2103 ( 
.A1(n_2090),
.A2(n_2083),
.B(n_1952),
.Y(n_2103)
);

AOI221xp5_ASAP7_75t_L g2104 ( 
.A1(n_2089),
.A2(n_2098),
.B1(n_2091),
.B2(n_2088),
.C(n_2097),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2094),
.Y(n_2105)
);

INVx1_ASAP7_75t_SL g2106 ( 
.A(n_2095),
.Y(n_2106)
);

OAI211xp5_ASAP7_75t_SL g2107 ( 
.A1(n_2092),
.A2(n_2083),
.B(n_1963),
.C(n_1950),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2101),
.B(n_1924),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2099),
.Y(n_2109)
);

AOI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_2103),
.A2(n_2100),
.B(n_2092),
.Y(n_2110)
);

AOI211xp5_ASAP7_75t_L g2111 ( 
.A1(n_2107),
.A2(n_2096),
.B(n_1963),
.C(n_1966),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2105),
.Y(n_2112)
);

AOI221xp5_ASAP7_75t_L g2113 ( 
.A1(n_2104),
.A2(n_2106),
.B1(n_2102),
.B2(n_2108),
.C(n_2109),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2103),
.B(n_1948),
.Y(n_2114)
);

O2A1O1Ixp33_ASAP7_75t_L g2115 ( 
.A1(n_2107),
.A2(n_1948),
.B(n_1950),
.C(n_1893),
.Y(n_2115)
);

AOI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_2104),
.A2(n_1976),
.B1(n_1970),
.B2(n_1969),
.Y(n_2116)
);

NAND4xp75_ASAP7_75t_L g2117 ( 
.A(n_2104),
.B(n_1976),
.C(n_1970),
.D(n_1969),
.Y(n_2117)
);

OAI221xp5_ASAP7_75t_SL g2118 ( 
.A1(n_2103),
.A2(n_1873),
.B1(n_1968),
.B2(n_1888),
.C(n_1912),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2112),
.Y(n_2119)
);

XNOR2x1_ASAP7_75t_L g2120 ( 
.A(n_2117),
.B(n_1848),
.Y(n_2120)
);

NAND2x1_ASAP7_75t_L g2121 ( 
.A(n_2116),
.B(n_1968),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_2113),
.A2(n_1897),
.B1(n_1920),
.B2(n_1918),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2114),
.Y(n_2123)
);

AND5x1_ASAP7_75t_L g2124 ( 
.A(n_2111),
.B(n_2110),
.C(n_2115),
.D(n_2118),
.E(n_1897),
.Y(n_2124)
);

OAI22xp5_ASAP7_75t_L g2125 ( 
.A1(n_2122),
.A2(n_1897),
.B1(n_1888),
.B2(n_1893),
.Y(n_2125)
);

NOR3xp33_ASAP7_75t_L g2126 ( 
.A(n_2123),
.B(n_1897),
.C(n_1873),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2119),
.Y(n_2127)
);

NOR3xp33_ASAP7_75t_L g2128 ( 
.A(n_2121),
.B(n_1897),
.C(n_1923),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2127),
.B(n_2120),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2125),
.Y(n_2130)
);

AOI22xp33_ASAP7_75t_L g2131 ( 
.A1(n_2130),
.A2(n_2126),
.B1(n_2128),
.B2(n_2124),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2131),
.A2(n_2129),
.B1(n_1888),
.B2(n_1892),
.Y(n_2132)
);

AO22x2_ASAP7_75t_L g2133 ( 
.A1(n_2131),
.A2(n_1883),
.B1(n_1909),
.B2(n_1896),
.Y(n_2133)
);

INVx4_ASAP7_75t_L g2134 ( 
.A(n_2133),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_2132),
.B(n_1918),
.Y(n_2135)
);

AOI22xp33_ASAP7_75t_L g2136 ( 
.A1(n_2135),
.A2(n_1868),
.B1(n_1920),
.B2(n_1896),
.Y(n_2136)
);

XNOR2x1_ASAP7_75t_L g2137 ( 
.A(n_2136),
.B(n_2134),
.Y(n_2137)
);

OAI21xp5_ASAP7_75t_L g2138 ( 
.A1(n_2137),
.A2(n_1923),
.B(n_1920),
.Y(n_2138)
);

INVxp67_ASAP7_75t_L g2139 ( 
.A(n_2138),
.Y(n_2139)
);

AOI221xp5_ASAP7_75t_L g2140 ( 
.A1(n_2139),
.A2(n_1921),
.B1(n_1919),
.B2(n_1902),
.C(n_1917),
.Y(n_2140)
);

AOI211xp5_ASAP7_75t_L g2141 ( 
.A1(n_2140),
.A2(n_1706),
.B(n_1708),
.C(n_1698),
.Y(n_2141)
);


endmodule