module fake_netlist_6_3701_n_1147 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1147);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1147;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_222;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_1017;
wire n_1004;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_901;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_1121;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_934;
wire n_482;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_811;
wire n_1060;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx2_ASAP7_75t_L g222 ( 
.A(n_43),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_207),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_91),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_130),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_69),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_85),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_165),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_49),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_48),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_143),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_119),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_103),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_96),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_19),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_169),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_201),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_25),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_101),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_11),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_6),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_97),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_93),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_31),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_64),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_22),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_127),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_105),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_198),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_99),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_139),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_155),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_21),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_132),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_150),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_98),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_100),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_16),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_47),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_205),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_24),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_46),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_95),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_200),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_86),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_173),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_121),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_104),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_2),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_212),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_40),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_168),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_219),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_166),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_220),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_123),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_114),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_175),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_70),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_188),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_60),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_12),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_141),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_82),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_65),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_52),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_176),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_0),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_81),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_133),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_162),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_57),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_236),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_223),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_237),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_259),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_232),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_241),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_227),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_222),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_239),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_232),
.Y(n_306)
);

BUFx2_ASAP7_75t_SL g307 ( 
.A(n_272),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_257),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_272),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_273),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_242),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_228),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_230),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_240),
.Y(n_315)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_245),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_264),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_265),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_266),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_247),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_269),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_288),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_262),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_222),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_270),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_224),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_224),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_243),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_243),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_288),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_257),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_234),
.B(n_0),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_260),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_260),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_234),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_279),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_279),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_283),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_305),
.B(n_257),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_302),
.B(n_291),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_306),
.A2(n_289),
.B1(n_256),
.B2(n_229),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_295),
.B(n_225),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_328),
.A2(n_253),
.B1(n_293),
.B2(n_251),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_329),
.Y(n_350)
);

CKINVDCx6p67_ASAP7_75t_R g351 ( 
.A(n_334),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_329),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_229),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_256),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_292),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_298),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_298),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_330),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_226),
.Y(n_361)
);

CKINVDCx8_ASAP7_75t_R g362 ( 
.A(n_307),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_231),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_294),
.Y(n_365)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_296),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_300),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_335),
.A2(n_290),
.B1(n_286),
.B2(n_284),
.Y(n_368)
);

OAI21x1_ASAP7_75t_L g369 ( 
.A1(n_336),
.A2(n_235),
.B(n_233),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_337),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_303),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_308),
.A2(n_282),
.B1(n_280),
.B2(n_278),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_313),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_314),
.B(n_238),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_315),
.B(n_277),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_244),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_297),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_317),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_318),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_322),
.B(n_276),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_324),
.A2(n_248),
.B(n_246),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_325),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_306),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_320),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_326),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_342),
.B(n_249),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_342),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_316),
.B(n_250),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_299),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_309),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_362),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_353),
.B(n_309),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_362),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_393),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_R g404 ( 
.A(n_392),
.B(n_310),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_386),
.Y(n_405)
);

BUFx8_ASAP7_75t_SL g406 ( 
.A(n_387),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_348),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_397),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_R g409 ( 
.A(n_392),
.B(n_310),
.Y(n_409)
);

NAND2xp33_ASAP7_75t_R g410 ( 
.A(n_383),
.B(n_384),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_351),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_351),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_347),
.B(n_312),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_397),
.Y(n_414)
);

CKINVDCx11_ASAP7_75t_R g415 ( 
.A(n_397),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_391),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_393),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_391),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_365),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_365),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_348),
.Y(n_421)
);

AO22x2_ASAP7_75t_L g422 ( 
.A1(n_389),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_391),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_348),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_391),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_343),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_391),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_397),
.Y(n_429)
);

INVxp33_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_383),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_384),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_395),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_348),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_366),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_361),
.B(n_312),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_379),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_345),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_377),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_366),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_372),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_357),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_354),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_356),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_392),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_366),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_366),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_396),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_366),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_379),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_350),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_378),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_366),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_367),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_367),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_394),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_350),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_345),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_394),
.B(n_252),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_390),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_378),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_389),
.B(n_323),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_361),
.B(n_323),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_368),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_349),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_350),
.Y(n_468)
);

OA21x2_ASAP7_75t_L g469 ( 
.A1(n_369),
.A2(n_258),
.B(n_255),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_378),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_368),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_390),
.B(n_356),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_462),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_416),
.B(n_356),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_400),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_356),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_452),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_405),
.Y(n_479)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_452),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_462),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_344),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_410),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_433),
.B(n_333),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_419),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_418),
.B(n_374),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_406),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_437),
.B(n_364),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_420),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_425),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_451),
.B(n_364),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_439),
.Y(n_492)
);

AND2x6_ASAP7_75t_L g493 ( 
.A(n_436),
.B(n_344),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_443),
.B(n_333),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_406),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_423),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_426),
.B(n_374),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_404),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_428),
.B(n_374),
.Y(n_499)
);

BUFx4f_ASAP7_75t_L g500 ( 
.A(n_465),
.Y(n_500)
);

AO22x2_ASAP7_75t_L g501 ( 
.A1(n_444),
.A2(n_396),
.B1(n_374),
.B2(n_376),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_452),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_449),
.B(n_376),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_466),
.A2(n_385),
.B1(n_369),
.B2(n_371),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_461),
.B(n_446),
.Y(n_505)
);

AND2x2_ASAP7_75t_SL g506 ( 
.A(n_408),
.B(n_385),
.Y(n_506)
);

BUFx4f_ASAP7_75t_L g507 ( 
.A(n_399),
.Y(n_507)
);

AND2x6_ASAP7_75t_L g508 ( 
.A(n_403),
.B(n_388),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_427),
.B(n_375),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_460),
.B(n_385),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_402),
.B(n_417),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_435),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_466),
.A2(n_385),
.B1(n_371),
.B2(n_382),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_453),
.B(n_378),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_463),
.B(n_371),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_435),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_467),
.B(n_373),
.Y(n_517)
);

AND2x4_ASAP7_75t_SL g518 ( 
.A(n_414),
.B(n_373),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_471),
.A2(n_261),
.B1(n_275),
.B2(n_274),
.Y(n_519)
);

BUFx10_ASAP7_75t_L g520 ( 
.A(n_464),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_455),
.B(n_380),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_470),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_471),
.A2(n_360),
.B1(n_370),
.B2(n_355),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_456),
.B(n_263),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_457),
.B(n_388),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_422),
.B(n_380),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_403),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_407),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_407),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_421),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_421),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_411),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_412),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_424),
.B(n_363),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_434),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_458),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_414),
.B(n_381),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g540 ( 
.A(n_441),
.B(n_268),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_458),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_413),
.B(n_381),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_429),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_431),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_468),
.B(n_363),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_468),
.B(n_363),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_440),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_430),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_429),
.B(n_358),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_422),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_398),
.B(n_358),
.Y(n_551)
);

CKINVDCx8_ASAP7_75t_R g552 ( 
.A(n_401),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_432),
.B(n_359),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_442),
.B(n_271),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_447),
.B(n_359),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_422),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_469),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_448),
.B(n_355),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_509),
.B(n_409),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_542),
.B(n_440),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_521),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_527),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_527),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_552),
.Y(n_564)
);

A2O1A1Ixp33_ASAP7_75t_L g565 ( 
.A1(n_482),
.A2(n_454),
.B(n_450),
.C(n_459),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_518),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_543),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_483),
.B(n_438),
.Y(n_568)
);

AO22x2_ASAP7_75t_L g569 ( 
.A1(n_550),
.A2(n_438),
.B1(n_459),
.B2(n_415),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_541),
.Y(n_570)
);

AO22x2_ASAP7_75t_L g571 ( 
.A1(n_556),
.A2(n_415),
.B1(n_3),
.B2(n_4),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_525),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_474),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_476),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_539),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_479),
.Y(n_576)
);

A2O1A1Ixp33_ASAP7_75t_L g577 ( 
.A1(n_517),
.A2(n_346),
.B(n_370),
.C(n_360),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_490),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_488),
.B(n_346),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_557),
.B(n_477),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_488),
.B(n_35),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_493),
.A2(n_469),
.B1(n_370),
.B2(n_360),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_492),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_541),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_548),
.B(n_36),
.Y(n_585)
);

AO22x2_ASAP7_75t_L g586 ( 
.A1(n_549),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_553),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_531),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_511),
.B(n_469),
.Y(n_589)
);

NAND2x1p5_ASAP7_75t_L g590 ( 
.A(n_496),
.B(n_539),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_505),
.B(n_5),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_497),
.B(n_355),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_549),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_496),
.B(n_37),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_533),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_538),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_485),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_499),
.B(n_355),
.Y(n_598)
);

AO22x2_ASAP7_75t_L g599 ( 
.A1(n_526),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_489),
.B(n_38),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_551),
.Y(n_601)
);

OR2x2_ASAP7_75t_SL g602 ( 
.A(n_503),
.B(n_7),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_538),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_522),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_515),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_511),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_536),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_493),
.B(n_355),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_551),
.B(n_360),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_528),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_500),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_535),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_493),
.B(n_360),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_532),
.Y(n_614)
);

O2A1O1Ixp33_ASAP7_75t_L g615 ( 
.A1(n_475),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_513),
.A2(n_352),
.B1(n_350),
.B2(n_370),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_493),
.B(n_370),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_500),
.B(n_350),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_529),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_530),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_L g621 ( 
.A1(n_507),
.A2(n_352),
.B1(n_10),
.B2(n_11),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_502),
.Y(n_622)
);

NAND2x1p5_ASAP7_75t_L g623 ( 
.A(n_507),
.B(n_352),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_545),
.Y(n_624)
);

NAND2x1p5_ASAP7_75t_L g625 ( 
.A(n_512),
.B(n_352),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_561),
.B(n_498),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_568),
.A2(n_486),
.B1(n_540),
.B2(n_484),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_560),
.B(n_501),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_592),
.A2(n_481),
.B(n_473),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_608),
.A2(n_481),
.B(n_473),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_587),
.B(n_494),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_572),
.B(n_501),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_601),
.B(n_544),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_593),
.B(n_520),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_613),
.A2(n_510),
.B(n_478),
.Y(n_635)
);

A2O1A1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_591),
.A2(n_506),
.B(n_555),
.C(n_491),
.Y(n_636)
);

A2O1A1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_565),
.A2(n_491),
.B(n_554),
.C(n_504),
.Y(n_637)
);

BUFx4f_ASAP7_75t_L g638 ( 
.A(n_590),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_567),
.Y(n_639)
);

NOR3xp33_ASAP7_75t_L g640 ( 
.A(n_559),
.B(n_524),
.C(n_519),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_617),
.A2(n_558),
.B(n_480),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_606),
.B(n_520),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_618),
.A2(n_480),
.B(n_514),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_611),
.B(n_532),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_574),
.B(n_523),
.Y(n_645)
);

AO32x2_ASAP7_75t_L g646 ( 
.A1(n_616),
.A2(n_547),
.A3(n_516),
.B1(n_512),
.B2(n_526),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_575),
.B(n_534),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_562),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_605),
.A2(n_578),
.B1(n_583),
.B2(n_576),
.Y(n_649)
);

AOI21x1_ASAP7_75t_L g650 ( 
.A1(n_598),
.A2(n_546),
.B(n_537),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_579),
.Y(n_651)
);

AOI21x1_ASAP7_75t_L g652 ( 
.A1(n_589),
.A2(n_537),
.B(n_480),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_612),
.A2(n_547),
.B1(n_516),
.B2(n_537),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_624),
.A2(n_609),
.B(n_585),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_570),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_585),
.B(n_534),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_624),
.A2(n_352),
.B(n_508),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_577),
.A2(n_508),
.B(n_487),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_562),
.A2(n_508),
.B(n_41),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_573),
.B(n_495),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_SL g661 ( 
.A1(n_621),
.A2(n_508),
.B(n_120),
.C(n_122),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_563),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_563),
.A2(n_42),
.B(n_39),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_581),
.B(n_44),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_580),
.A2(n_50),
.B(n_45),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_604),
.B(n_9),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_597),
.B(n_12),
.Y(n_667)
);

O2A1O1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_615),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_584),
.A2(n_53),
.B(n_51),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_579),
.B(n_13),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_573),
.B(n_14),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_573),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_584),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_588),
.Y(n_674)
);

BUFx8_ASAP7_75t_L g675 ( 
.A(n_614),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_581),
.B(n_15),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_594),
.Y(n_677)
);

OAI21xp33_ASAP7_75t_L g678 ( 
.A1(n_586),
.A2(n_16),
.B(n_17),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_600),
.B(n_17),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_564),
.B(n_18),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_600),
.A2(n_55),
.B(n_54),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_582),
.A2(n_58),
.B(n_56),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_594),
.B(n_59),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_566),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_580),
.A2(n_136),
.B1(n_218),
.B2(n_217),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_602),
.B(n_18),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_588),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_596),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_SL g689 ( 
.A(n_627),
.B(n_623),
.C(n_625),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_635),
.A2(n_595),
.B(n_620),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_662),
.Y(n_691)
);

O2A1O1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_636),
.A2(n_607),
.B(n_595),
.C(n_620),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_SL g693 ( 
.A(n_678),
.B(n_686),
.C(n_680),
.Y(n_693)
);

INVx8_ASAP7_75t_L g694 ( 
.A(n_677),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_639),
.Y(n_695)
);

NAND2x1p5_ASAP7_75t_L g696 ( 
.A(n_638),
.B(n_677),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_677),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_651),
.B(n_569),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_654),
.A2(n_603),
.B(n_622),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_640),
.B(n_610),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_638),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_674),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_687),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_647),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_631),
.B(n_626),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_649),
.B(n_619),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_648),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_673),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_655),
.Y(n_709)
);

CKINVDCx16_ASAP7_75t_R g710 ( 
.A(n_660),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_637),
.A2(n_622),
.B(n_586),
.C(n_599),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_678),
.A2(n_599),
.B(n_571),
.C(n_569),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_634),
.B(n_571),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_679),
.A2(n_580),
.B1(n_20),
.B2(n_21),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_632),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_644),
.B(n_580),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_SL g717 ( 
.A1(n_665),
.A2(n_137),
.B(n_216),
.C(n_215),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_681),
.A2(n_19),
.B(n_20),
.C(n_22),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_675),
.Y(n_719)
);

OAI22x1_ASAP7_75t_L g720 ( 
.A1(n_656),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_671),
.B(n_23),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_629),
.A2(n_140),
.B(n_214),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_688),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_642),
.B(n_676),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_688),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_645),
.B(n_26),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_628),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_630),
.A2(n_643),
.B(n_657),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_683),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_668),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_672),
.B(n_61),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_688),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_666),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_667),
.Y(n_734)
);

OR2x6_ASAP7_75t_L g735 ( 
.A(n_664),
.B(n_62),
.Y(n_735)
);

OAI21xp33_ASAP7_75t_L g736 ( 
.A1(n_670),
.A2(n_30),
.B(n_32),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_653),
.B(n_32),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_641),
.A2(n_147),
.B(n_213),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_652),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_682),
.A2(n_146),
.B(n_211),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_650),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_658),
.A2(n_33),
.B(n_34),
.C(n_63),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_684),
.B(n_33),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_659),
.A2(n_661),
.B(n_669),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_675),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_SL g746 ( 
.A1(n_685),
.A2(n_34),
.B1(n_66),
.B2(n_67),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_663),
.A2(n_68),
.B(n_71),
.Y(n_747)
);

OAI21xp33_ASAP7_75t_SL g748 ( 
.A1(n_633),
.A2(n_72),
.B(n_73),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_691),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_695),
.Y(n_750)
);

BUFx4_ASAP7_75t_SL g751 ( 
.A(n_719),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_702),
.Y(n_752)
);

BUFx12f_ASAP7_75t_L g753 ( 
.A(n_745),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_704),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_723),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_725),
.Y(n_756)
);

BUFx12f_ASAP7_75t_L g757 ( 
.A(n_701),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_707),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_705),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_704),
.Y(n_760)
);

BUFx12f_ASAP7_75t_L g761 ( 
.A(n_701),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_723),
.Y(n_762)
);

INVx6_ASAP7_75t_L g763 ( 
.A(n_704),
.Y(n_763)
);

BUFx4_ASAP7_75t_R g764 ( 
.A(n_703),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_723),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_736),
.A2(n_646),
.B1(n_75),
.B2(n_76),
.Y(n_766)
);

CKINVDCx6p67_ASAP7_75t_R g767 ( 
.A(n_694),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_694),
.Y(n_768)
);

BUFx2_ASAP7_75t_SL g769 ( 
.A(n_732),
.Y(n_769)
);

BUFx12f_ASAP7_75t_L g770 ( 
.A(n_697),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_732),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_708),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_732),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_709),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_696),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_693),
.B(n_646),
.Y(n_776)
);

INVx6_ASAP7_75t_SL g777 ( 
.A(n_731),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_741),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_697),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_697),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_731),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_739),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_715),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_710),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_706),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_733),
.Y(n_786)
);

OR2x6_ASAP7_75t_L g787 ( 
.A(n_711),
.B(n_646),
.Y(n_787)
);

CKINVDCx11_ASAP7_75t_R g788 ( 
.A(n_735),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_735),
.Y(n_789)
);

INVx6_ASAP7_75t_L g790 ( 
.A(n_698),
.Y(n_790)
);

NAND2x1p5_ASAP7_75t_L g791 ( 
.A(n_716),
.B(n_74),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_734),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_746),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_700),
.Y(n_794)
);

BUFx4_ASAP7_75t_SL g795 ( 
.A(n_720),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_737),
.Y(n_796)
);

BUFx12f_ASAP7_75t_L g797 ( 
.A(n_721),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_726),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_692),
.Y(n_799)
);

CKINVDCx11_ASAP7_75t_R g800 ( 
.A(n_727),
.Y(n_800)
);

BUFx12f_ASAP7_75t_L g801 ( 
.A(n_743),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_713),
.Y(n_802)
);

INVx8_ASAP7_75t_L g803 ( 
.A(n_748),
.Y(n_803)
);

INVx8_ASAP7_75t_L g804 ( 
.A(n_718),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_724),
.Y(n_805)
);

NAND2x1p5_ASAP7_75t_L g806 ( 
.A(n_699),
.B(n_738),
.Y(n_806)
);

OAI22xp33_ASAP7_75t_SL g807 ( 
.A1(n_729),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_689),
.Y(n_808)
);

INVx5_ASAP7_75t_L g809 ( 
.A(n_717),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_690),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_712),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_714),
.B(n_87),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_742),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_728),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_722),
.Y(n_815)
);

BUFx6f_ASAP7_75t_SL g816 ( 
.A(n_730),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_747),
.Y(n_817)
);

NAND2x1p5_ASAP7_75t_L g818 ( 
.A(n_740),
.B(n_88),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_744),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_800),
.B(n_89),
.C(n_90),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_778),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_805),
.A2(n_92),
.B1(n_94),
.B2(n_102),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_SL g823 ( 
.A(n_793),
.B(n_106),
.C(n_107),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_779),
.Y(n_824)
);

NAND3x1_ASAP7_75t_L g825 ( 
.A(n_789),
.B(n_108),
.C(n_109),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_806),
.A2(n_110),
.B(n_111),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_806),
.A2(n_112),
.B(n_113),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_SL g828 ( 
.A1(n_793),
.A2(n_797),
.B1(n_801),
.B2(n_784),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_778),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_749),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_752),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_794),
.B(n_115),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_813),
.A2(n_116),
.B(n_117),
.C(n_118),
.Y(n_833)
);

OA21x2_ASAP7_75t_L g834 ( 
.A1(n_819),
.A2(n_124),
.B(n_125),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_798),
.B(n_796),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_814),
.A2(n_126),
.B(n_128),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_749),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_782),
.Y(n_838)
);

OAI21x1_ASAP7_75t_L g839 ( 
.A1(n_814),
.A2(n_129),
.B(n_131),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_750),
.Y(n_840)
);

OAI21x1_ASAP7_75t_L g841 ( 
.A1(n_815),
.A2(n_808),
.B(n_818),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_764),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_816),
.A2(n_134),
.B1(n_135),
.B2(n_138),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_808),
.A2(n_142),
.B(n_144),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_818),
.A2(n_145),
.B(n_149),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_750),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_760),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_800),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_794),
.B(n_154),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_781),
.B(n_156),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_792),
.Y(n_851)
);

CKINVDCx11_ASAP7_75t_R g852 ( 
.A(n_753),
.Y(n_852)
);

INVxp67_ASAP7_75t_SL g853 ( 
.A(n_792),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_816),
.A2(n_789),
.B1(n_811),
.B2(n_813),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_751),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_756),
.Y(n_856)
);

INVx4_ASAP7_75t_SL g857 ( 
.A(n_757),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_798),
.A2(n_157),
.B(n_158),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_783),
.B(n_159),
.Y(n_859)
);

OAI22xp33_ASAP7_75t_L g860 ( 
.A1(n_804),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_783),
.B(n_164),
.Y(n_861)
);

AO21x2_ASAP7_75t_L g862 ( 
.A1(n_799),
.A2(n_167),
.B(n_170),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_758),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_SL g864 ( 
.A1(n_812),
.A2(n_759),
.B(n_754),
.C(n_799),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_751),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_759),
.A2(n_171),
.B1(n_172),
.B2(n_174),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_786),
.B(n_177),
.Y(n_867)
);

OAI21xp33_ASAP7_75t_L g868 ( 
.A1(n_766),
.A2(n_178),
.B(n_179),
.Y(n_868)
);

INVx3_ASAP7_75t_SL g869 ( 
.A(n_767),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_770),
.Y(n_870)
);

AO21x1_ASAP7_75t_L g871 ( 
.A1(n_807),
.A2(n_180),
.B(n_181),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_SL g872 ( 
.A1(n_804),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_804),
.A2(n_185),
.B(n_186),
.C(n_187),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_774),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_781),
.B(n_189),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_785),
.A2(n_190),
.B(n_191),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_764),
.Y(n_877)
);

OR2x6_ASAP7_75t_L g878 ( 
.A(n_763),
.B(n_192),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_786),
.B(n_193),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_853),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_835),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_821),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_841),
.A2(n_791),
.B(n_766),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_840),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_SL g885 ( 
.A1(n_828),
.A2(n_803),
.B1(n_802),
.B2(n_776),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_821),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_829),
.Y(n_887)
);

AOI21x1_ASAP7_75t_L g888 ( 
.A1(n_854),
.A2(n_787),
.B(n_772),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_831),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_838),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_826),
.A2(n_791),
.B(n_817),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_840),
.Y(n_892)
);

OAI21x1_ASAP7_75t_L g893 ( 
.A1(n_827),
.A2(n_810),
.B(n_809),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_863),
.B(n_787),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_874),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_868),
.A2(n_788),
.B1(n_802),
.B2(n_790),
.Y(n_896)
);

AO21x2_ASAP7_75t_L g897 ( 
.A1(n_823),
.A2(n_809),
.B(n_787),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_852),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_SL g899 ( 
.A1(n_842),
.A2(n_803),
.B1(n_802),
.B2(n_790),
.Y(n_899)
);

AOI21x1_ASAP7_75t_L g900 ( 
.A1(n_871),
.A2(n_809),
.B(n_803),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_851),
.B(n_790),
.Y(n_901)
);

INVxp33_ASAP7_75t_L g902 ( 
.A(n_840),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_830),
.Y(n_903)
);

OA21x2_ASAP7_75t_L g904 ( 
.A1(n_876),
.A2(n_836),
.B(n_839),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_870),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_837),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_834),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_842),
.B(n_788),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_847),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_834),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_879),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_862),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_867),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_846),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_856),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_824),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_855),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_824),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_870),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_845),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_844),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_870),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_869),
.Y(n_923)
);

BUFx2_ASAP7_75t_SL g924 ( 
.A(n_877),
.Y(n_924)
);

BUFx4f_ASAP7_75t_SL g925 ( 
.A(n_865),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_864),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_R g927 ( 
.A(n_898),
.B(n_877),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_880),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_894),
.B(n_857),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_881),
.B(n_802),
.Y(n_930)
);

NAND2xp33_ASAP7_75t_R g931 ( 
.A(n_926),
.B(n_878),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_887),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_914),
.B(n_849),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_889),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_909),
.B(n_760),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_914),
.B(n_832),
.Y(n_936)
);

CKINVDCx16_ASAP7_75t_R g937 ( 
.A(n_898),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_899),
.B(n_820),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_913),
.B(n_859),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_886),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_902),
.B(n_857),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_884),
.B(n_878),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_924),
.A2(n_848),
.B1(n_872),
.B2(n_858),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_886),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_R g945 ( 
.A(n_917),
.B(n_761),
.Y(n_945)
);

CKINVDCx16_ASAP7_75t_R g946 ( 
.A(n_923),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_892),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_924),
.B(n_825),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_SL g949 ( 
.A(n_905),
.B(n_861),
.Y(n_949)
);

NOR3xp33_ASAP7_75t_SL g950 ( 
.A(n_917),
.B(n_822),
.C(n_860),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_895),
.B(n_875),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_894),
.B(n_763),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_925),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_890),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_894),
.B(n_763),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_905),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_R g957 ( 
.A(n_900),
.B(n_770),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_SL g958 ( 
.A1(n_885),
.A2(n_843),
.B(n_873),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_887),
.B(n_875),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_SL g960 ( 
.A1(n_897),
.A2(n_809),
.B1(n_795),
.B2(n_850),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_890),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_932),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_929),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_928),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_929),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_932),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_929),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_933),
.B(n_915),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_948),
.Y(n_969)
);

NAND2x1_ASAP7_75t_L g970 ( 
.A(n_948),
.B(n_912),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_940),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_944),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_934),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_954),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_947),
.B(n_888),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_933),
.B(n_911),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_930),
.B(n_888),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_936),
.B(n_911),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_936),
.B(n_913),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_961),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_956),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_941),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_935),
.B(n_903),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_956),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_959),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_971),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_972),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_962),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_982),
.Y(n_989)
);

AO21x2_ASAP7_75t_L g990 ( 
.A1(n_975),
.A2(n_957),
.B(n_912),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_973),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_967),
.B(n_952),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_962),
.Y(n_993)
);

OA21x2_ASAP7_75t_L g994 ( 
.A1(n_975),
.A2(n_910),
.B(n_907),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_972),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_971),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_966),
.Y(n_997)
);

NOR2x1_ASAP7_75t_SL g998 ( 
.A(n_969),
.B(n_948),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_979),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_974),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_974),
.Y(n_1001)
);

AOI21xp33_ASAP7_75t_L g1002 ( 
.A1(n_970),
.A2(n_931),
.B(n_938),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_967),
.B(n_955),
.Y(n_1003)
);

NAND4xp25_ASAP7_75t_L g1004 ( 
.A(n_968),
.B(n_960),
.C(n_938),
.D(n_958),
.Y(n_1004)
);

OAI211xp5_ASAP7_75t_SL g1005 ( 
.A1(n_1002),
.A2(n_999),
.B(n_950),
.C(n_964),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_1004),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_991),
.B(n_977),
.Y(n_1007)
);

NAND4xp25_ASAP7_75t_L g1008 ( 
.A(n_986),
.B(n_931),
.C(n_908),
.D(n_896),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_996),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_992),
.B(n_967),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_987),
.Y(n_1011)
);

OAI221xp5_ASAP7_75t_L g1012 ( 
.A1(n_989),
.A2(n_943),
.B1(n_969),
.B2(n_970),
.C(n_949),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_992),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_987),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_992),
.B(n_963),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_989),
.B(n_937),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_1010),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_1015),
.B(n_998),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_1013),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_1012),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_1006),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1016),
.B(n_998),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1011),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1009),
.B(n_995),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_1007),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1020),
.B(n_977),
.Y(n_1026)
);

NAND4xp75_ASAP7_75t_L g1027 ( 
.A(n_1022),
.B(n_1005),
.C(n_1014),
.D(n_994),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1018),
.B(n_1003),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1023),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_1021),
.A2(n_1005),
.B(n_1012),
.Y(n_1030)
);

AOI32xp33_ASAP7_75t_SL g1031 ( 
.A1(n_1024),
.A2(n_995),
.A3(n_1001),
.B1(n_1000),
.B2(n_1008),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_1021),
.A2(n_969),
.B1(n_965),
.B2(n_963),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1029),
.B(n_1025),
.Y(n_1033)
);

INVxp33_ASAP7_75t_L g1034 ( 
.A(n_1026),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1028),
.B(n_1017),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1032),
.Y(n_1036)
);

NAND4xp25_ASAP7_75t_L g1037 ( 
.A(n_1030),
.B(n_1019),
.C(n_1024),
.D(n_965),
.Y(n_1037)
);

CKINVDCx16_ASAP7_75t_R g1038 ( 
.A(n_1031),
.Y(n_1038)
);

CKINVDCx16_ASAP7_75t_R g1039 ( 
.A(n_1027),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1029),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_1030),
.B(n_946),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1029),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_L g1043 ( 
.A(n_1030),
.B(n_969),
.C(n_833),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_1035),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_1039),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_1033),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1033),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1040),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1042),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1036),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1038),
.B(n_990),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1034),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1052),
.Y(n_1053)
);

OAI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1051),
.A2(n_1043),
.B1(n_1037),
.B2(n_1041),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1045),
.B(n_1003),
.Y(n_1055)
);

OAI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_1045),
.A2(n_969),
.B1(n_982),
.B2(n_949),
.C(n_953),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_1046),
.A2(n_1003),
.B(n_981),
.C(n_883),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_1044),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1050),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1047),
.A2(n_990),
.B1(n_922),
.B2(n_919),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_1055),
.B(n_1048),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1058),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1053),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1059),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1054),
.B(n_1049),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_1061),
.B(n_1060),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1062),
.Y(n_1067)
);

HAxp5_ASAP7_75t_SL g1068 ( 
.A(n_1063),
.B(n_1056),
.CON(n_1068),
.SN(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1064),
.B(n_1057),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1065),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1062),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1067),
.Y(n_1072)
);

NAND3xp33_ASAP7_75t_L g1073 ( 
.A(n_1068),
.B(n_905),
.C(n_919),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1071),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_1066),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1070),
.B(n_990),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1075),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_L g1078 ( 
.A(n_1073),
.B(n_1069),
.Y(n_1078)
);

OAI211xp5_ASAP7_75t_L g1079 ( 
.A1(n_1074),
.A2(n_945),
.B(n_927),
.C(n_768),
.Y(n_1079)
);

OAI21xp33_ASAP7_75t_SL g1080 ( 
.A1(n_1076),
.A2(n_993),
.B(n_988),
.Y(n_1080)
);

AOI21xp33_ASAP7_75t_SL g1081 ( 
.A1(n_1072),
.A2(n_945),
.B(n_994),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_1077),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_1078),
.B(n_905),
.C(n_919),
.Y(n_1083)
);

NAND4xp25_ASAP7_75t_L g1084 ( 
.A(n_1079),
.B(n_768),
.C(n_850),
.D(n_775),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_1081),
.Y(n_1085)
);

AOI31xp33_ASAP7_75t_L g1086 ( 
.A1(n_1080),
.A2(n_866),
.A3(n_927),
.B(n_939),
.Y(n_1086)
);

AOI32xp33_ASAP7_75t_L g1087 ( 
.A1(n_1078),
.A2(n_981),
.A3(n_775),
.B1(n_942),
.B2(n_984),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1077),
.A2(n_994),
.B(n_993),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1077),
.A2(n_922),
.B1(n_919),
.B2(n_905),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1082),
.B(n_988),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_L g1091 ( 
.A(n_1085),
.B(n_939),
.C(n_976),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1083),
.A2(n_997),
.B(n_919),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1084),
.A2(n_978),
.B(n_997),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_1089),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_1088),
.Y(n_1095)
);

AOI222xp33_ASAP7_75t_L g1096 ( 
.A1(n_1086),
.A2(n_922),
.B1(n_795),
.B2(n_985),
.C1(n_984),
.C2(n_921),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1087),
.B(n_966),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_L g1098 ( 
.A(n_1085),
.B(n_951),
.C(n_921),
.Y(n_1098)
);

NOR3xp33_ASAP7_75t_L g1099 ( 
.A(n_1094),
.B(n_900),
.C(n_777),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_1090),
.B(n_1091),
.Y(n_1100)
);

NOR3x1_ASAP7_75t_L g1101 ( 
.A(n_1097),
.B(n_983),
.C(n_985),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_1093),
.B(n_922),
.Y(n_1102)
);

AOI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_1095),
.A2(n_922),
.B(n_195),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1096),
.B(n_980),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_SL g1105 ( 
.A(n_1098),
.B(n_957),
.C(n_777),
.Y(n_1105)
);

INVxp67_ASAP7_75t_L g1106 ( 
.A(n_1092),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1094),
.B(n_780),
.Y(n_1107)
);

AND2x2_ASAP7_75t_SL g1108 ( 
.A(n_1090),
.B(n_780),
.Y(n_1108)
);

OAI211xp5_ASAP7_75t_L g1109 ( 
.A1(n_1094),
.A2(n_779),
.B(n_780),
.C(n_755),
.Y(n_1109)
);

NOR2x1_ASAP7_75t_L g1110 ( 
.A(n_1095),
.B(n_769),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_1110),
.B(n_779),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1107),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_1100),
.Y(n_1113)
);

XOR2xp5_ASAP7_75t_L g1114 ( 
.A(n_1102),
.B(n_194),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_1106),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_1103),
.Y(n_1116)
);

CKINVDCx16_ASAP7_75t_R g1117 ( 
.A(n_1105),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1104),
.A2(n_897),
.B(n_920),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1113),
.A2(n_1108),
.B(n_1099),
.Y(n_1119)
);

NAND4xp75_ASAP7_75t_L g1120 ( 
.A(n_1112),
.B(n_1101),
.C(n_1109),
.D(n_199),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1114),
.Y(n_1121)
);

OAI22x1_ASAP7_75t_L g1122 ( 
.A1(n_1115),
.A2(n_980),
.B1(n_918),
.B2(n_916),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_SL g1123 ( 
.A1(n_1117),
.A2(n_779),
.B1(n_780),
.B2(n_755),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_SL g1124 ( 
.A1(n_1116),
.A2(n_773),
.B1(n_762),
.B2(n_765),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1111),
.Y(n_1125)
);

XOR2x1_ASAP7_75t_L g1126 ( 
.A(n_1125),
.B(n_1111),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_SL g1127 ( 
.A1(n_1119),
.A2(n_1118),
.B(n_773),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1120),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1126),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_1129),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1130),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1131),
.A2(n_1128),
.B(n_1121),
.C(n_1127),
.Y(n_1132)
);

BUFx2_ASAP7_75t_SL g1133 ( 
.A(n_1131),
.Y(n_1133)
);

INVx3_ASAP7_75t_SL g1134 ( 
.A(n_1131),
.Y(n_1134)
);

AOI222xp33_ASAP7_75t_L g1135 ( 
.A1(n_1134),
.A2(n_1123),
.B1(n_1124),
.B2(n_1122),
.C1(n_773),
.C2(n_771),
.Y(n_1135)
);

AOI222xp33_ASAP7_75t_L g1136 ( 
.A1(n_1133),
.A2(n_773),
.B1(n_771),
.B2(n_765),
.C1(n_762),
.C2(n_755),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1132),
.A2(n_196),
.B(n_197),
.Y(n_1137)
);

OAI222xp33_ASAP7_75t_L g1138 ( 
.A1(n_1132),
.A2(n_920),
.B1(n_910),
.B2(n_907),
.C1(n_206),
.C2(n_208),
.Y(n_1138)
);

AOI222xp33_ASAP7_75t_L g1139 ( 
.A1(n_1138),
.A2(n_755),
.B1(n_771),
.B2(n_765),
.C1(n_762),
.C2(n_210),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1137),
.A2(n_762),
.B1(n_771),
.B2(n_765),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1135),
.A2(n_897),
.B1(n_904),
.B2(n_901),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_SL g1142 ( 
.A1(n_1136),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1139),
.B(n_209),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1140),
.A2(n_221),
.B(n_893),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1141),
.A2(n_904),
.B1(n_901),
.B2(n_893),
.Y(n_1145)
);

AOI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1143),
.A2(n_1142),
.B1(n_1145),
.B2(n_1144),
.C(n_882),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1146),
.A2(n_904),
.B1(n_891),
.B2(n_906),
.Y(n_1147)
);


endmodule