module fake_jpeg_31035_n_117 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_117);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_53),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_56),
.Y(n_67)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_62),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_73),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_41),
.B1(n_40),
.B2(n_37),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_1),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_19),
.B1(n_35),
.B2(n_34),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_18),
.B1(n_32),
.B2(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_82),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_2),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_17),
.B1(n_30),
.B2(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_84),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_3),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_70),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_4),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_6),
.C(n_7),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_5),
.Y(n_99)
);

MAJx2_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_98),
.C(n_92),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_85),
.B(n_95),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_5),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_90),
.C(n_102),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_107),
.A2(n_90),
.B1(n_87),
.B2(n_86),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_109),
.C(n_110),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_106),
.C(n_102),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_101),
.C(n_103),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_111),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_100),
.C(n_10),
.Y(n_115)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_8),
.A3(n_12),
.B1(n_15),
.B2(n_16),
.C1(n_20),
.C2(n_21),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_22),
.Y(n_117)
);


endmodule