module fake_aes_2626_n_578 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_578);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_578;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g70 ( .A(n_60), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_42), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_27), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_29), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_3), .Y(n_74) );
CKINVDCx16_ASAP7_75t_R g75 ( .A(n_56), .Y(n_75) );
INVx1_ASAP7_75t_SL g76 ( .A(n_10), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_28), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_14), .Y(n_78) );
INVxp33_ASAP7_75t_L g79 ( .A(n_13), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_9), .Y(n_80) );
OR2x2_ASAP7_75t_L g81 ( .A(n_26), .B(n_11), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_31), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_13), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_51), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_69), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_30), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_19), .Y(n_87) );
CKINVDCx14_ASAP7_75t_R g88 ( .A(n_45), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_23), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_36), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_17), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_64), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_62), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_35), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_40), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_50), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_38), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_9), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_43), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_66), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_59), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_25), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_3), .Y(n_103) );
INVxp33_ASAP7_75t_SL g104 ( .A(n_12), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_67), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_0), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_11), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_14), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_32), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_16), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_10), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_34), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_110), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_72), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_72), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_102), .Y(n_116) );
INVx3_ASAP7_75t_L g117 ( .A(n_110), .Y(n_117) );
INVx3_ASAP7_75t_L g118 ( .A(n_83), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_73), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_73), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_70), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_91), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_77), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_91), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_102), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_77), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_85), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_90), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_75), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_82), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_82), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_79), .B(n_0), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_84), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_74), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_105), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_83), .B(n_1), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_96), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_105), .B(n_1), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_109), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_109), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_88), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_93), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_74), .B(n_2), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_71), .B(n_2), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_78), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_93), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_78), .B(n_4), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_146), .B(n_95), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_113), .B(n_108), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_117), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_116), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_126), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_117), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_116), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_126), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_116), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_126), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_129), .A2(n_111), .B1(n_87), .B2(n_108), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_126), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_113), .B(n_112), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_126), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_116), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_145), .B(n_112), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_116), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_122), .A2(n_107), .B1(n_106), .B2(n_87), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_126), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_146), .B(n_81), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_117), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_149), .B(n_99), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_132), .A2(n_104), .B1(n_103), .B2(n_98), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_114), .B(n_115), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_114), .B(n_94), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_116), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
INVx1_ASAP7_75t_SL g183 ( .A(n_124), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_139), .B(n_146), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_142), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
OR2x6_ASAP7_75t_L g190 ( .A(n_132), .B(n_81), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_142), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_134), .B(n_148), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_143), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_143), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_121), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_139), .B(n_107), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_139), .B(n_106), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_143), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_166), .B(n_134), .Y(n_199) );
NOR3xp33_ASAP7_75t_SL g200 ( .A(n_195), .B(n_128), .C(n_127), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_167), .Y(n_201) );
BUFx12f_ASAP7_75t_L g202 ( .A(n_167), .Y(n_202) );
NOR3xp33_ASAP7_75t_SL g203 ( .A(n_172), .B(n_140), .C(n_164), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_155), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_192), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_162), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_192), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_184), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_188), .B(n_148), .Y(n_209) );
NOR3xp33_ASAP7_75t_SL g210 ( .A(n_170), .B(n_177), .C(n_147), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_183), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_184), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_162), .Y(n_213) );
OR2x6_ASAP7_75t_L g214 ( .A(n_190), .B(n_139), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_153), .B(n_139), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_153), .B(n_190), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_162), .B(n_144), .Y(n_217) );
NOR2xp33_ASAP7_75t_R g218 ( .A(n_151), .B(n_117), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_155), .Y(n_219) );
OAI22xp5_ASAP7_75t_SL g220 ( .A1(n_178), .A2(n_76), .B1(n_150), .B2(n_80), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_196), .B(n_115), .Y(n_221) );
INVxp67_ASAP7_75t_L g222 ( .A(n_190), .Y(n_222) );
INVxp67_ASAP7_75t_L g223 ( .A(n_190), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_162), .Y(n_224) );
BUFx4f_ASAP7_75t_L g225 ( .A(n_175), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_190), .Y(n_226) );
INVx4_ASAP7_75t_L g227 ( .A(n_184), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_155), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_196), .B(n_135), .Y(n_229) );
BUFx8_ASAP7_75t_L g230 ( .A(n_151), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_196), .B(n_135), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_178), .A2(n_123), .B1(n_119), .B2(n_130), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_197), .B(n_123), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_158), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_197), .B(n_136), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_181), .Y(n_236) );
NOR2xp33_ASAP7_75t_R g237 ( .A(n_151), .B(n_119), .Y(n_237) );
BUFx3_ASAP7_75t_L g238 ( .A(n_158), .Y(n_238) );
BUFx5_ASAP7_75t_L g239 ( .A(n_151), .Y(n_239) );
INVxp67_ASAP7_75t_SL g240 ( .A(n_175), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_197), .B(n_120), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_158), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_181), .Y(n_243) );
INVxp67_ASAP7_75t_L g244 ( .A(n_180), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_197), .B(n_120), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_151), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_184), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_175), .B(n_130), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_151), .B(n_137), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_176), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_176), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_176), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_194), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_151), .A2(n_137), .B1(n_136), .B2(n_133), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_208), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_206), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_212), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_244), .B(n_179), .Y(n_258) );
INVxp67_ASAP7_75t_L g259 ( .A(n_201), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_199), .B(n_133), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_212), .Y(n_261) );
INVxp67_ASAP7_75t_L g262 ( .A(n_201), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_225), .B(n_150), .Y(n_263) );
BUFx12f_ASAP7_75t_L g264 ( .A(n_202), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_206), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_247), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_248), .B(n_141), .Y(n_267) );
NAND3xp33_ASAP7_75t_L g268 ( .A(n_210), .B(n_131), .C(n_138), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_202), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_247), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_225), .B(n_131), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_214), .A2(n_138), .B1(n_131), .B2(n_125), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_216), .B(n_138), .Y(n_273) );
INVxp67_ASAP7_75t_SL g274 ( .A(n_240), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_206), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_214), .A2(n_143), .B1(n_80), .B2(n_125), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_216), .B(n_118), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_211), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_208), .B(n_118), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_225), .B(n_118), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_246), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_224), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_230), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_211), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_224), .Y(n_285) );
OR2x6_ASAP7_75t_L g286 ( .A(n_214), .B(n_118), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_214), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_224), .Y(n_288) );
BUFx2_ASAP7_75t_SL g289 ( .A(n_239), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_237), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_207), .B(n_125), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_254), .A2(n_143), .B1(n_97), .B2(n_100), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_230), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_207), .A2(n_143), .B1(n_89), .B2(n_101), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_200), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_208), .Y(n_296) );
CKINVDCx16_ASAP7_75t_R g297 ( .A(n_226), .Y(n_297) );
BUFx12f_ASAP7_75t_L g298 ( .A(n_230), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_204), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_209), .B(n_92), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_227), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_254), .B(n_185), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_233), .A2(n_157), .B1(n_165), .B2(n_193), .Y(n_303) );
INVx6_ASAP7_75t_L g304 ( .A(n_281), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_277), .A2(n_220), .B1(n_205), .B2(n_222), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_277), .A2(n_223), .B1(n_227), .B2(n_215), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_293), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_293), .B(n_227), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_272), .A2(n_235), .B1(n_231), .B2(n_229), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_257), .Y(n_310) );
INVx4_ASAP7_75t_L g311 ( .A(n_286), .Y(n_311) );
AOI22xp33_ASAP7_75t_SL g312 ( .A1(n_278), .A2(n_217), .B1(n_218), .B2(n_215), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_272), .A2(n_221), .B1(n_245), .B2(n_241), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_293), .B(n_246), .Y(n_314) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_259), .A2(n_203), .B1(n_232), .B2(n_249), .C(n_213), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_286), .B(n_213), .Y(n_316) );
BUFx12f_ASAP7_75t_L g317 ( .A(n_264), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_298), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_286), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_281), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_257), .B(n_239), .Y(n_321) );
INVx1_ASAP7_75t_SL g322 ( .A(n_280), .Y(n_322) );
INVx4_ASAP7_75t_SL g323 ( .A(n_298), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_277), .A2(n_239), .B1(n_252), .B2(n_238), .Y(n_324) );
OA21x2_ASAP7_75t_L g325 ( .A1(n_268), .A2(n_161), .B(n_171), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_260), .A2(n_252), .B(n_204), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_299), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_273), .B(n_280), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_286), .B(n_238), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_277), .A2(n_239), .B1(n_251), .B2(n_250), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_262), .A2(n_239), .B1(n_251), .B2(n_250), .Y(n_331) );
NAND2x1_ASAP7_75t_L g332 ( .A(n_299), .B(n_219), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_287), .A2(n_239), .B1(n_219), .B2(n_242), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_261), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_261), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_273), .B(n_239), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_299), .Y(n_337) );
OAI211xp5_ASAP7_75t_L g338 ( .A1(n_305), .A2(n_300), .B(n_284), .C(n_295), .Y(n_338) );
OA21x2_ASAP7_75t_L g339 ( .A1(n_326), .A2(n_268), .B(n_302), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_328), .B(n_258), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_304), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_320), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_327), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_315), .A2(n_309), .B1(n_274), .B2(n_322), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_328), .B(n_266), .Y(n_345) );
INVx5_ASAP7_75t_L g346 ( .A(n_320), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_313), .A2(n_258), .B1(n_291), .B2(n_269), .C(n_266), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_313), .A2(n_279), .B1(n_291), .B2(n_264), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_310), .A2(n_270), .B1(n_279), .B2(n_267), .C(n_294), .Y(n_349) );
OAI211xp5_ASAP7_75t_L g350 ( .A1(n_312), .A2(n_292), .B(n_263), .C(n_276), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_322), .A2(n_279), .B1(n_283), .B2(n_270), .Y(n_351) );
NAND3xp33_ASAP7_75t_L g352 ( .A(n_331), .B(n_292), .C(n_303), .Y(n_352) );
NAND3xp33_ASAP7_75t_L g353 ( .A(n_310), .B(n_303), .C(n_271), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_334), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_334), .B(n_297), .Y(n_355) );
NAND3xp33_ASAP7_75t_L g356 ( .A(n_335), .B(n_185), .C(n_189), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_335), .B(n_297), .Y(n_357) );
A2O1A1Ixp33_ASAP7_75t_L g358 ( .A1(n_327), .A2(n_275), .B(n_265), .C(n_256), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_327), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_337), .B(n_301), .Y(n_360) );
OAI211xp5_ASAP7_75t_SL g361 ( .A1(n_306), .A2(n_255), .B(n_154), .C(n_187), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_343), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_359), .B(n_337), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_345), .B(n_337), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_346), .B(n_345), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_355), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g367 ( .A1(n_347), .A2(n_307), .B(n_319), .C(n_316), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_346), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_344), .A2(n_311), .B1(n_329), .B2(n_319), .Y(n_369) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_338), .A2(n_311), .B1(n_318), .B2(n_307), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_354), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_357), .A2(n_311), .B1(n_318), .B2(n_317), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_343), .B(n_336), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_360), .B(n_336), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_360), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_340), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_358), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_358), .Y(n_378) );
NAND2xp33_ASAP7_75t_R g379 ( .A(n_341), .B(n_323), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_348), .A2(n_308), .B1(n_323), .B2(n_318), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_351), .A2(n_324), .B1(n_330), .B2(n_255), .C(n_333), .Y(n_381) );
A2O1A1Ixp33_ASAP7_75t_L g382 ( .A1(n_350), .A2(n_316), .B(n_308), .C(n_314), .Y(n_382) );
OAI33xp33_ASAP7_75t_L g383 ( .A1(n_361), .A2(n_160), .A3(n_154), .B1(n_157), .B2(n_163), .B3(n_165), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_342), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_346), .Y(n_385) );
AO21x1_ASAP7_75t_SL g386 ( .A1(n_346), .A2(n_321), .B(n_323), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_353), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_342), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_342), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g390 ( .A1(n_349), .A2(n_255), .B1(n_296), .B2(n_329), .C(n_285), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_352), .B(n_308), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_388), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_375), .B(n_341), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_371), .B(n_341), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_371), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_374), .B(n_342), .Y(n_396) );
OAI33xp33_ASAP7_75t_L g397 ( .A1(n_376), .A2(n_163), .A3(n_191), .B1(n_187), .B2(n_186), .B3(n_182), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_364), .B(n_346), .Y(n_398) );
OAI31xp33_ASAP7_75t_L g399 ( .A1(n_372), .A2(n_316), .A3(n_314), .B(n_296), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_362), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_366), .A2(n_316), .B1(n_329), .B2(n_314), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_384), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_368), .Y(n_403) );
INVx4_ASAP7_75t_L g404 ( .A(n_368), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_374), .B(n_342), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_380), .A2(n_329), .B1(n_317), .B2(n_304), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_373), .B(n_339), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_373), .B(n_320), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_387), .B(n_181), .C(n_169), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_365), .B(n_320), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_365), .B(n_320), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_368), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_365), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_385), .Y(n_414) );
OR2x6_ASAP7_75t_L g415 ( .A(n_369), .B(n_304), .Y(n_415) );
NAND4xp25_ASAP7_75t_L g416 ( .A(n_382), .B(n_168), .C(n_173), .D(n_174), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_363), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_377), .B(n_325), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_377), .Y(n_419) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_370), .A2(n_288), .B1(n_332), .B2(n_356), .C(n_290), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_378), .B(n_325), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_379), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_378), .B(n_325), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_390), .A2(n_304), .B1(n_332), .B2(n_281), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_391), .B(n_325), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_367), .B(n_181), .C(n_169), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_389), .Y(n_427) );
OA21x2_ASAP7_75t_L g428 ( .A1(n_389), .A2(n_152), .B(n_156), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_381), .B(n_169), .C(n_185), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_395), .B(n_4), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_407), .B(n_388), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_407), .B(n_388), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_404), .B(n_388), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_425), .B(n_388), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_414), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_413), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_425), .B(n_386), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_393), .B(n_383), .Y(n_438) );
OAI221xp5_ASAP7_75t_L g439 ( .A1(n_401), .A2(n_275), .B1(n_256), .B2(n_282), .C(n_265), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_394), .Y(n_440) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_404), .B(n_386), .Y(n_441) );
AOI32xp33_ASAP7_75t_L g442 ( .A1(n_406), .A2(n_5), .A3(n_6), .B1(n_7), .B2(n_8), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_400), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_396), .B(n_5), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_414), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_396), .B(n_6), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_394), .Y(n_447) );
OAI33xp33_ASAP7_75t_L g448 ( .A1(n_393), .A2(n_7), .A3(n_8), .B1(n_12), .B2(n_15), .B3(n_16), .Y(n_448) );
NOR3xp33_ASAP7_75t_L g449 ( .A(n_416), .B(n_397), .C(n_420), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_413), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_398), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_408), .B(n_15), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_417), .B(n_17), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_398), .B(n_18), .Y(n_454) );
NOR2x1_ASAP7_75t_L g455 ( .A(n_404), .B(n_289), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_404), .B(n_18), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g457 ( .A(n_429), .B(n_152), .C(n_156), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_415), .B(n_63), .Y(n_458) );
NAND4xp25_ASAP7_75t_L g459 ( .A(n_399), .B(n_159), .C(n_161), .D(n_171), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_415), .B(n_411), .Y(n_460) );
INVx5_ASAP7_75t_L g461 ( .A(n_403), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_408), .B(n_20), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_419), .B(n_20), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_422), .B(n_21), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_405), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_402), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_402), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_427), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_464), .A2(n_429), .B(n_424), .C(n_426), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_451), .B(n_410), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_441), .B(n_412), .Y(n_471) );
NOR4xp25_ASAP7_75t_L g472 ( .A(n_464), .B(n_411), .C(n_418), .D(n_423), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_449), .A2(n_415), .B1(n_403), .B2(n_412), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_437), .B(n_412), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_437), .B(n_415), .Y(n_475) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_455), .B(n_409), .Y(n_476) );
AOI32xp33_ASAP7_75t_L g477 ( .A1(n_456), .A2(n_418), .A3(n_421), .B1(n_423), .B2(n_392), .Y(n_477) );
INVxp67_ASAP7_75t_L g478 ( .A(n_456), .Y(n_478) );
OAI21xp33_ASAP7_75t_L g479 ( .A1(n_442), .A2(n_415), .B(n_421), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_454), .B(n_22), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_468), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_440), .B(n_402), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_447), .B(n_392), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_461), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_465), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_450), .B(n_428), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g487 ( .A(n_458), .B(n_281), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_436), .B(n_428), .Y(n_488) );
O2A1O1Ixp5_ASAP7_75t_SL g489 ( .A1(n_430), .A2(n_191), .B(n_182), .C(n_173), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_443), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_444), .B(n_428), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_458), .A2(n_446), .B1(n_444), .B2(n_461), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_438), .B(n_169), .Y(n_493) );
AND2x4_ASAP7_75t_L g494 ( .A(n_460), .B(n_24), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_457), .A2(n_282), .B(n_275), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_453), .B(n_33), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_448), .A2(n_281), .B1(n_239), .B2(n_234), .Y(n_497) );
INVxp67_ASAP7_75t_L g498 ( .A(n_452), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_446), .Y(n_499) );
OAI332xp33_ASAP7_75t_L g500 ( .A1(n_463), .A2(n_198), .A3(n_194), .B1(n_242), .B2(n_234), .B3(n_228), .C1(n_253), .C2(n_47), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_435), .B(n_37), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_458), .A2(n_281), .B1(n_185), .B2(n_189), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_452), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_462), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_460), .A2(n_189), .B1(n_198), .B2(n_228), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_445), .B(n_39), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_431), .B(n_41), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_472), .B(n_431), .Y(n_508) );
NAND2xp33_ASAP7_75t_R g509 ( .A(n_471), .B(n_433), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_474), .B(n_432), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_485), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_478), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_490), .Y(n_513) );
AND2x2_ASAP7_75t_SL g514 ( .A(n_471), .B(n_433), .Y(n_514) );
NOR3xp33_ASAP7_75t_SL g515 ( .A(n_479), .B(n_439), .C(n_459), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_475), .B(n_461), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_499), .B(n_432), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_470), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_503), .B(n_434), .Y(n_519) );
AOI211xp5_ASAP7_75t_L g520 ( .A1(n_492), .A2(n_433), .B(n_434), .C(n_467), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_493), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_498), .B(n_461), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_504), .B(n_467), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_484), .B(n_461), .Y(n_524) );
NOR2x1p5_ASAP7_75t_SL g525 ( .A(n_486), .B(n_466), .Y(n_525) );
NAND2x1_ASAP7_75t_L g526 ( .A(n_476), .B(n_443), .Y(n_526) );
AOI21xp5_ASAP7_75t_SL g527 ( .A1(n_469), .A2(n_44), .B(n_46), .Y(n_527) );
OAI21xp5_ASAP7_75t_SL g528 ( .A1(n_473), .A2(n_48), .B(n_49), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_473), .Y(n_529) );
OAI21xp5_ASAP7_75t_SL g530 ( .A1(n_477), .A2(n_52), .B(n_53), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_491), .B(n_54), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_481), .Y(n_532) );
NOR2xp33_ASAP7_75t_R g533 ( .A(n_494), .B(n_55), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_487), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_482), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_512), .B(n_480), .Y(n_536) );
NAND3x2_ASAP7_75t_L g537 ( .A(n_516), .B(n_488), .C(n_500), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_515), .B(n_505), .C(n_496), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_529), .A2(n_483), .B1(n_507), .B2(n_501), .Y(n_539) );
XNOR2x1_ASAP7_75t_L g540 ( .A(n_518), .B(n_476), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_508), .B(n_502), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_530), .A2(n_506), .B(n_495), .Y(n_542) );
AOI21xp33_ASAP7_75t_SL g543 ( .A1(n_509), .A2(n_497), .B(n_58), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_535), .B(n_489), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_511), .B(n_57), .Y(n_545) );
OAI221xp5_ASAP7_75t_L g546 ( .A1(n_515), .A2(n_61), .B1(n_65), .B2(n_68), .C(n_236), .Y(n_546) );
NOR2x1p5_ASAP7_75t_L g547 ( .A(n_509), .B(n_236), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_513), .Y(n_548) );
AOI211xp5_ASAP7_75t_SL g549 ( .A1(n_527), .A2(n_528), .B(n_533), .C(n_531), .Y(n_549) );
XNOR2x1_ASAP7_75t_L g550 ( .A(n_522), .B(n_236), .Y(n_550) );
O2A1O1Ixp5_ASAP7_75t_L g551 ( .A1(n_524), .A2(n_243), .B(n_526), .C(n_532), .Y(n_551) );
INVxp67_ASAP7_75t_L g552 ( .A(n_540), .Y(n_552) );
AOI211xp5_ASAP7_75t_L g553 ( .A1(n_543), .A2(n_533), .B(n_521), .C(n_534), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_548), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_551), .B(n_514), .Y(n_555) );
NOR2xp67_ASAP7_75t_L g556 ( .A(n_546), .B(n_510), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_537), .A2(n_517), .B1(n_519), .B2(n_523), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_541), .Y(n_558) );
AND2x2_ASAP7_75t_SL g559 ( .A(n_549), .B(n_525), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_544), .B(n_513), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_544), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_547), .A2(n_550), .B1(n_539), .B2(n_542), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_536), .Y(n_563) );
AOI321xp33_ASAP7_75t_L g564 ( .A1(n_545), .A2(n_472), .A3(n_508), .B1(n_549), .B2(n_520), .C(n_541), .Y(n_564) );
OAI221xp5_ASAP7_75t_L g565 ( .A1(n_540), .A2(n_538), .B1(n_508), .B2(n_541), .C(n_530), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_552), .B(n_563), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_557), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_554), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_559), .A2(n_555), .B1(n_565), .B2(n_556), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_566), .B(n_558), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_568), .Y(n_571) );
NAND3xp33_ASAP7_75t_SL g572 ( .A(n_569), .B(n_564), .C(n_555), .Y(n_572) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_572), .A2(n_567), .B1(n_562), .B2(n_553), .C(n_561), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_571), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_573), .A2(n_567), .B1(n_570), .B2(n_559), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_574), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_576), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_577), .A2(n_575), .B(n_560), .Y(n_578) );
endmodule