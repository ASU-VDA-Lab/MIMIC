module fake_jpeg_548_n_22 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_22);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_22;

wire n_13;
wire n_21;
wire n_10;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

AND2x2_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_5),
.Y(n_7)
);

INVx1_ASAP7_75t_SL g8 ( 
.A(n_1),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_7),
.Y(n_13)
);

NAND2xp33_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_0),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_16),
.A2(n_9),
.B(n_7),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_13),
.Y(n_20)
);

AOI322xp5_ASAP7_75t_L g22 ( 
.A1(n_20),
.A2(n_21),
.A3(n_15),
.B1(n_12),
.B2(n_17),
.C1(n_0),
.C2(n_6),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_11),
.C(n_15),
.Y(n_21)
);


endmodule