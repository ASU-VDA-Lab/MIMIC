module fake_aes_12459_n_681 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_39, n_681);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_39;
output n_681;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_15), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_52), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_63), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_22), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_91), .Y(n_99) );
HB1xp67_ASAP7_75t_L g100 ( .A(n_1), .Y(n_100) );
CKINVDCx14_ASAP7_75t_R g101 ( .A(n_32), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_78), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_25), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_79), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_92), .Y(n_105) );
BUFx5_ASAP7_75t_L g106 ( .A(n_26), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_70), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_35), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_85), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_76), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_20), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_55), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_53), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_24), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_50), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_14), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_60), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_36), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_46), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_45), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_37), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_88), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_6), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_44), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_33), .Y(n_125) );
INVx1_ASAP7_75t_SL g126 ( .A(n_17), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_30), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_68), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_62), .Y(n_129) );
NOR2xp67_ASAP7_75t_L g130 ( .A(n_49), .B(n_23), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_5), .Y(n_131) );
INVxp67_ASAP7_75t_L g132 ( .A(n_0), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_89), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_59), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
OR2x2_ASAP7_75t_L g136 ( .A(n_94), .B(n_73), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_14), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_11), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_123), .B(n_0), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_111), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_128), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_112), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_116), .B(n_1), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_137), .B(n_2), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_98), .B(n_2), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_124), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_111), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_96), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_111), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_106), .Y(n_151) );
BUFx12f_ASAP7_75t_L g152 ( .A(n_103), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_106), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_138), .B(n_3), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_124), .B(n_3), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_97), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_140), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_149), .B(n_157), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_151), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_149), .B(n_98), .Y(n_162) );
NAND3xp33_ASAP7_75t_L g163 ( .A(n_156), .B(n_127), .C(n_135), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_143), .A2(n_118), .B1(n_133), .B2(n_112), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_151), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_156), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_140), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_157), .B(n_105), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_147), .B(n_125), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_156), .B(n_101), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_156), .A2(n_100), .B1(n_105), .B2(n_132), .Y(n_171) );
NAND3xp33_ASAP7_75t_L g172 ( .A(n_143), .B(n_108), .C(n_99), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_143), .B(n_101), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_143), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_153), .Y(n_177) );
OR2x6_ASAP7_75t_L g178 ( .A(n_139), .B(n_136), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_140), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_146), .A2(n_95), .B1(n_131), .B2(n_126), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_147), .Y(n_181) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_147), .Y(n_182) );
NOR2xp33_ASAP7_75t_SL g183 ( .A(n_178), .B(n_118), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_176), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_178), .A2(n_155), .B1(n_139), .B2(n_144), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_162), .B(n_152), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_178), .A2(n_155), .B1(n_144), .B2(n_133), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_166), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_160), .A2(n_145), .B(n_147), .C(n_110), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_168), .B(n_141), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_178), .B(n_145), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_162), .B(n_152), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_178), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_170), .B(n_152), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_177), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_176), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_170), .B(n_107), .Y(n_197) );
INVxp67_ASAP7_75t_L g198 ( .A(n_164), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_178), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_170), .B(n_109), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_160), .B(n_142), .Y(n_201) );
OAI22xp5_ASAP7_75t_SL g202 ( .A1(n_164), .A2(n_102), .B1(n_104), .B2(n_129), .Y(n_202) );
NOR2xp33_ASAP7_75t_SL g203 ( .A(n_166), .B(n_113), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_166), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_182), .B(n_114), .Y(n_205) );
O2A1O1Ixp5_ASAP7_75t_L g206 ( .A1(n_182), .A2(n_115), .B(n_119), .C(n_121), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_177), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_171), .B(n_117), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_163), .A2(n_134), .B1(n_122), .B2(n_125), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_173), .B(n_106), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_173), .B(n_106), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_176), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_176), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_159), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_188), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_195), .A2(n_207), .B(n_210), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_187), .A2(n_172), .B1(n_163), .B2(n_169), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_184), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_191), .B(n_172), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_198), .A2(n_169), .B(n_181), .C(n_180), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_184), .Y(n_221) );
AO31x2_ASAP7_75t_L g222 ( .A1(n_211), .A2(n_159), .A3(n_161), .B(n_165), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_191), .B(n_181), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_192), .B(n_181), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_195), .A2(n_177), .B(n_161), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_195), .A2(n_165), .B(n_175), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_188), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_196), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_196), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_187), .A2(n_175), .B1(n_174), .B2(n_130), .Y(n_230) );
INVx2_ASAP7_75t_SL g231 ( .A(n_191), .Y(n_231) );
O2A1O1Ixp5_ASAP7_75t_L g232 ( .A1(n_206), .A2(n_174), .B(n_179), .C(n_167), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_208), .B(n_4), .Y(n_233) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_207), .A2(n_179), .B(n_167), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_203), .B(n_106), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_188), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_191), .B(n_106), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_189), .A2(n_179), .B(n_167), .C(n_158), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_185), .A2(n_120), .B1(n_154), .B2(n_150), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_205), .B(n_106), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_207), .A2(n_158), .B(n_120), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_194), .B(n_4), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_186), .B(n_5), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_193), .A2(n_120), .B1(n_154), .B2(n_150), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_230), .B(n_193), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_234), .A2(n_214), .B(n_204), .Y(n_246) );
AOI21x1_ASAP7_75t_L g247 ( .A1(n_239), .A2(n_158), .B(n_214), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_230), .B(n_199), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_240), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_220), .A2(n_213), .B(n_199), .C(n_183), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_231), .B(n_201), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_218), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_216), .A2(n_213), .B(n_205), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_SL g254 ( .A1(n_235), .A2(n_200), .B(n_197), .C(n_204), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_225), .A2(n_203), .B(n_204), .Y(n_255) );
NAND2x1p5_ASAP7_75t_L g256 ( .A(n_215), .B(n_212), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_226), .A2(n_204), .B(n_212), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_221), .Y(n_258) );
NAND2x1p5_ASAP7_75t_L g259 ( .A(n_215), .B(n_212), .Y(n_259) );
NAND3xp33_ASAP7_75t_L g260 ( .A(n_242), .B(n_183), .C(n_201), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_219), .A2(n_188), .B(n_190), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_217), .A2(n_209), .B(n_202), .C(n_188), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_224), .A2(n_188), .B(n_202), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_228), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_217), .A2(n_154), .B(n_150), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_215), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_243), .B(n_6), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_222), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_251), .B(n_229), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_246), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_266), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_259), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_265), .A2(n_239), .B(n_238), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_251), .B(n_222), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_252), .Y(n_275) );
OA21x2_ASAP7_75t_L g276 ( .A1(n_250), .A2(n_232), .B(n_237), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_246), .Y(n_277) );
OR2x6_ASAP7_75t_L g278 ( .A(n_268), .B(n_227), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g279 ( .A(n_268), .B(n_227), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_259), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_260), .A2(n_233), .B1(n_223), .B2(n_236), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_245), .B(n_222), .Y(n_282) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_250), .A2(n_241), .B(n_244), .Y(n_283) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_247), .A2(n_154), .B(n_150), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_258), .B(n_227), .Y(n_285) );
INVx4_ASAP7_75t_L g286 ( .A(n_259), .Y(n_286) );
NAND2x1_ASAP7_75t_L g287 ( .A(n_255), .B(n_120), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_264), .B(n_61), .Y(n_288) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_247), .A2(n_154), .B(n_150), .Y(n_289) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_270), .A2(n_263), .B(n_248), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_274), .B(n_267), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_284), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_274), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_274), .B(n_253), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_284), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_279), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_284), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_279), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_282), .B(n_249), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_284), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_279), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_269), .A2(n_261), .B1(n_257), .B2(n_254), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_278), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_278), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_275), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_278), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_286), .B(n_266), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_286), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_279), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_287), .A2(n_256), .B(n_262), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_275), .B(n_256), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_282), .B(n_7), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_278), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_282), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_301), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_305), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_293), .B(n_278), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_296), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_305), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_293), .B(n_278), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_292), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_294), .B(n_278), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_292), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_292), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_295), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_296), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_315), .B(n_288), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_294), .B(n_270), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_313), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_295), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_294), .B(n_270), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_315), .B(n_288), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_299), .B(n_288), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_313), .B(n_277), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_295), .Y(n_336) );
AND2x4_ASAP7_75t_SL g337 ( .A(n_309), .B(n_286), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_297), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_297), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_297), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_301), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_313), .B(n_277), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_300), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_300), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_296), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_291), .B(n_277), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_291), .B(n_285), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_299), .B(n_280), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_300), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_306), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_306), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_309), .B(n_280), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_290), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_312), .B(n_288), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_310), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_298), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_290), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_324), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_317), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_329), .B(n_307), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_317), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_324), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_348), .B(n_312), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_329), .B(n_303), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_332), .B(n_303), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_348), .B(n_309), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_347), .B(n_309), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_330), .B(n_304), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_347), .B(n_304), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_346), .B(n_314), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_332), .B(n_318), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_320), .B(n_314), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_320), .Y(n_374) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_349), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_335), .B(n_310), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_335), .B(n_307), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_342), .B(n_290), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_318), .B(n_290), .Y(n_379) );
BUFx4f_ASAP7_75t_L g380 ( .A(n_337), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_321), .B(n_298), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_342), .B(n_298), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_323), .B(n_302), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_349), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_349), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_324), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_321), .A2(n_288), .B1(n_308), .B2(n_281), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_323), .B(n_302), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_322), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_322), .B(n_308), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_325), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_325), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_331), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_349), .B(n_289), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_331), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_338), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_338), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_340), .B(n_308), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_340), .B(n_343), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_343), .B(n_311), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_344), .B(n_289), .Y(n_401) );
OAI21xp5_ASAP7_75t_L g402 ( .A1(n_344), .A2(n_281), .B(n_311), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_351), .B(n_289), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_351), .B(n_289), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_352), .B(n_308), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_356), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_356), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_352), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_346), .B(n_269), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_325), .B(n_289), .Y(n_410) );
AOI33xp33_ASAP7_75t_L g411 ( .A1(n_354), .A2(n_254), .A3(n_8), .B1(n_9), .B2(n_10), .B3(n_11), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_353), .B(n_285), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_326), .B(n_311), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_326), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_327), .B(n_286), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_326), .B(n_284), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_345), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_319), .B(n_7), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_336), .B(n_276), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_336), .B(n_276), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_336), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_339), .B(n_276), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_337), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_372), .B(n_339), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_396), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
NOR2xp67_ASAP7_75t_L g427 ( .A(n_423), .B(n_339), .Y(n_427) );
INVx3_ASAP7_75t_SL g428 ( .A(n_423), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_408), .B(n_350), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_372), .B(n_350), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_372), .B(n_350), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_365), .B(n_353), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_359), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_360), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_359), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_360), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_370), .B(n_334), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_362), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_365), .B(n_327), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_371), .B(n_334), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_362), .B(n_328), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_384), .Y(n_442) );
OAI21xp5_ASAP7_75t_SL g443 ( .A1(n_418), .A2(n_337), .B(n_355), .Y(n_443) );
INVxp33_ASAP7_75t_SL g444 ( .A(n_380), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_374), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_379), .B(n_354), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_374), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_366), .B(n_328), .Y(n_448) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_387), .B(n_355), .C(n_333), .D(n_358), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_389), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_389), .Y(n_451) );
HB1xp67_ASAP7_75t_SL g452 ( .A(n_380), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_380), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_371), .B(n_333), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_364), .B(n_327), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_411), .B(n_358), .C(n_140), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_393), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_393), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_366), .B(n_357), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_395), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_395), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_368), .B(n_357), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_417), .B(n_357), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_399), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_367), .B(n_316), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_373), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_359), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_417), .B(n_316), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_390), .B(n_341), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_398), .B(n_341), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_363), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_416), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_363), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_363), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_391), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_369), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_391), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_409), .B(n_319), .Y(n_478) );
NOR2x1_ASAP7_75t_L g479 ( .A(n_415), .B(n_319), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_379), .B(n_286), .Y(n_480) );
NAND2x1p5_ASAP7_75t_L g481 ( .A(n_385), .B(n_271), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_379), .B(n_283), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_406), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_391), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_416), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_378), .B(n_276), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_378), .B(n_276), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_379), .B(n_283), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_383), .B(n_283), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_382), .B(n_272), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_377), .B(n_272), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_369), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_377), .B(n_272), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_405), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_381), .B(n_271), .Y(n_495) );
NOR2x1_ASAP7_75t_R g496 ( .A(n_406), .B(n_271), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_414), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_383), .B(n_276), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_388), .B(n_8), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_400), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_381), .B(n_271), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_388), .B(n_9), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_427), .B(n_361), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_425), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_464), .B(n_414), .Y(n_505) );
OR2x6_ASAP7_75t_L g506 ( .A(n_453), .B(n_407), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_425), .Y(n_507) );
OAI31xp67_ASAP7_75t_L g508 ( .A1(n_443), .A2(n_392), .A3(n_386), .B(n_13), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_500), .B(n_361), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_426), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_452), .A2(n_361), .B1(n_375), .B2(n_407), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_424), .B(n_431), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_426), .Y(n_513) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_479), .B(n_410), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_476), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_492), .Y(n_516) );
NOR2xp67_ASAP7_75t_L g517 ( .A(n_500), .B(n_410), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_472), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_466), .B(n_421), .Y(n_519) );
AND3x2_ASAP7_75t_L g520 ( .A(n_502), .B(n_394), .C(n_400), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_502), .A2(n_381), .B1(n_412), .B2(n_400), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_494), .B(n_421), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_431), .B(n_381), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_434), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_432), .B(n_376), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_436), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_438), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_445), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_444), .A2(n_402), .B(n_400), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_439), .B(n_413), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_459), .B(n_413), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_447), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_450), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_451), .Y(n_534) );
INVxp67_ASAP7_75t_L g535 ( .A(n_468), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_428), .B(n_10), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_457), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_472), .B(n_385), .Y(n_538) );
OR2x6_ASAP7_75t_L g539 ( .A(n_463), .B(n_401), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_485), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_428), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_446), .B(n_419), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_458), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_460), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_446), .B(n_422), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_SL g546 ( .A1(n_444), .A2(n_386), .B(n_392), .C(n_287), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_485), .B(n_420), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_461), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_497), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_430), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_429), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_478), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_L g553 ( .A1(n_499), .A2(n_404), .B(n_403), .C(n_401), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_489), .B(n_420), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_440), .B(n_403), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_437), .B(n_404), .Y(n_556) );
INVxp67_ASAP7_75t_SL g557 ( .A(n_442), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_455), .B(n_12), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_495), .B(n_422), .Y(n_559) );
INVxp67_ASAP7_75t_SL g560 ( .A(n_442), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_483), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_454), .Y(n_562) );
XNOR2x1_ASAP7_75t_L g563 ( .A(n_490), .B(n_12), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_501), .B(n_394), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_469), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_480), .B(n_271), .Y(n_566) );
NOR3xp33_ASAP7_75t_L g567 ( .A(n_456), .B(n_273), .C(n_15), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_470), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_448), .B(n_154), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_489), .B(n_283), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_441), .B(n_283), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_500), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_465), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_455), .A2(n_271), .B1(n_283), .B2(n_17), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_504), .B(n_433), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_519), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_569), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_541), .B(n_463), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_541), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_507), .B(n_482), .Y(n_581) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_539), .A2(n_449), .B1(n_462), .B2(n_498), .Y(n_582) );
NOR2xp67_ASAP7_75t_L g583 ( .A(n_511), .B(n_468), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_523), .B(n_488), .Y(n_584) );
OAI211xp5_ASAP7_75t_L g585 ( .A1(n_536), .A2(n_462), .B(n_488), .C(n_487), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_521), .A2(n_493), .B1(n_491), .B2(n_480), .Y(n_586) );
AOI21xp33_ASAP7_75t_L g587 ( .A1(n_558), .A2(n_496), .B(n_16), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_521), .A2(n_480), .B1(n_486), .B2(n_471), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_505), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_510), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_512), .B(n_484), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_513), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_506), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_551), .B(n_484), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_535), .A2(n_435), .B1(n_477), .B2(n_475), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_522), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_518), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_561), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_552), .A2(n_435), .B1(n_477), .B2(n_475), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_562), .B(n_563), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_522), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_567), .B(n_433), .C(n_474), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_508), .A2(n_474), .B(n_473), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_553), .B(n_473), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_550), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g606 ( .A1(n_529), .A2(n_471), .B1(n_467), .B2(n_481), .C(n_150), .Y(n_606) );
AOI322xp5_ASAP7_75t_L g607 ( .A1(n_554), .A2(n_467), .A3(n_148), .B1(n_140), .B2(n_19), .C1(n_13), .C2(n_16), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_549), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_515), .A2(n_148), .B1(n_140), .B2(n_481), .C(n_271), .Y(n_609) );
INVxp67_ASAP7_75t_SL g610 ( .A(n_557), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_565), .B(n_148), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_524), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_526), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_527), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_528), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_506), .Y(n_616) );
AOI222xp33_ASAP7_75t_L g617 ( .A1(n_511), .A2(n_148), .B1(n_18), .B2(n_19), .C1(n_273), .C2(n_271), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_556), .B(n_148), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_532), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_516), .B(n_18), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_582), .A2(n_520), .B1(n_539), .B2(n_509), .Y(n_621) );
AOI21xp33_ASAP7_75t_L g622 ( .A1(n_580), .A2(n_514), .B(n_506), .Y(n_622) );
OAI322xp33_ASAP7_75t_L g623 ( .A1(n_598), .A2(n_568), .A3(n_573), .B1(n_560), .B2(n_555), .C1(n_570), .C2(n_534), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_611), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_603), .A2(n_574), .B1(n_537), .B2(n_548), .C(n_543), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_593), .B(n_616), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_604), .A2(n_574), .B1(n_533), .B2(n_544), .C(n_572), .Y(n_627) );
AOI211xp5_ASAP7_75t_L g628 ( .A1(n_587), .A2(n_517), .B(n_503), .C(n_546), .Y(n_628) );
AOI222xp33_ASAP7_75t_L g629 ( .A1(n_583), .A2(n_572), .B1(n_538), .B2(n_503), .C1(n_509), .C2(n_571), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_576), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_587), .A2(n_539), .B(n_571), .Y(n_631) );
O2A1O1Ixp33_ASAP7_75t_L g632 ( .A1(n_600), .A2(n_540), .B(n_547), .C(n_525), .Y(n_632) );
AOI21xp33_ASAP7_75t_SL g633 ( .A1(n_578), .A2(n_566), .B(n_531), .Y(n_633) );
AOI222xp33_ASAP7_75t_L g634 ( .A1(n_593), .A2(n_545), .B1(n_542), .B2(n_564), .C1(n_559), .C2(n_530), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_606), .A2(n_273), .B(n_148), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_616), .A2(n_21), .B1(n_27), .B2(n_28), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_610), .A2(n_29), .B(n_31), .C(n_34), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_585), .A2(n_38), .B(n_39), .C(n_40), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_618), .Y(n_639) );
OAI211xp5_ASAP7_75t_SL g640 ( .A1(n_607), .A2(n_41), .B(n_42), .C(n_43), .Y(n_640) );
O2A1O1Ixp33_ASAP7_75t_L g641 ( .A1(n_620), .A2(n_617), .B(n_592), .C(n_590), .Y(n_641) );
OAI21xp33_ASAP7_75t_L g642 ( .A1(n_588), .A2(n_47), .B(n_48), .Y(n_642) );
AOI21xp33_ASAP7_75t_L g643 ( .A1(n_617), .A2(n_51), .B(n_54), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_581), .B(n_56), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_586), .A2(n_57), .B(n_58), .Y(n_645) );
A2O1A1Ixp33_ASAP7_75t_L g646 ( .A1(n_602), .A2(n_64), .B(n_65), .C(n_66), .Y(n_646) );
NAND3xp33_ASAP7_75t_SL g647 ( .A(n_609), .B(n_67), .C(n_69), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_579), .B(n_71), .Y(n_648) );
NAND3xp33_ASAP7_75t_SL g649 ( .A(n_595), .B(n_93), .C(n_74), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_594), .A2(n_72), .B(n_75), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_605), .B(n_77), .Y(n_651) );
AOI21xp33_ASAP7_75t_SL g652 ( .A1(n_608), .A2(n_80), .B(n_81), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g653 ( .A(n_577), .B(n_82), .C(n_83), .D(n_84), .Y(n_653) );
OAI211xp5_ASAP7_75t_L g654 ( .A1(n_599), .A2(n_87), .B(n_90), .C(n_601), .Y(n_654) );
AOI22xp33_ASAP7_75t_SL g655 ( .A1(n_589), .A2(n_596), .B1(n_584), .B2(n_591), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_575), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_612), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_657) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_619), .A2(n_583), .B(n_541), .C(n_587), .Y(n_658) );
NOR4xp25_ASAP7_75t_L g659 ( .A(n_632), .B(n_623), .C(n_641), .D(n_658), .Y(n_659) );
NAND3xp33_ASAP7_75t_SL g660 ( .A(n_628), .B(n_625), .C(n_631), .Y(n_660) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_627), .A2(n_626), .B1(n_621), .B2(n_624), .C1(n_639), .C2(n_656), .Y(n_661) );
OAI211xp5_ASAP7_75t_SL g662 ( .A1(n_629), .A2(n_631), .B(n_622), .C(n_643), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_657), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_633), .A2(n_646), .B(n_654), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_634), .B(n_630), .Y(n_665) );
NOR3xp33_ASAP7_75t_L g666 ( .A(n_660), .B(n_636), .C(n_637), .Y(n_666) );
NAND4xp75_ASAP7_75t_L g667 ( .A(n_664), .B(n_650), .C(n_635), .D(n_651), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_663), .B(n_655), .Y(n_668) );
NAND3x1_ASAP7_75t_L g669 ( .A(n_665), .B(n_635), .C(n_648), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_668), .B(n_662), .Y(n_670) );
XNOR2xp5_ASAP7_75t_L g671 ( .A(n_667), .B(n_659), .Y(n_671) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_666), .B(n_661), .C(n_645), .D(n_653), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_671), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_670), .Y(n_674) );
AO22x2_ASAP7_75t_L g675 ( .A1(n_673), .A2(n_672), .B1(n_669), .B2(n_638), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_674), .Y(n_676) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_676), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_677), .A2(n_673), .B(n_675), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_678), .A2(n_649), .B1(n_640), .B2(n_652), .C(n_642), .Y(n_679) );
OR2x6_ASAP7_75t_L g680 ( .A(n_679), .B(n_644), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_680), .A2(n_647), .B1(n_575), .B2(n_597), .Y(n_681) );
endmodule