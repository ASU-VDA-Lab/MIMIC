module fake_jpeg_12655_n_584 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_584);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_584;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_548;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_60),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_62),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_64),
.Y(n_191)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_67),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_68),
.Y(n_193)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_71),
.Y(n_180)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_10),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_80),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_75),
.Y(n_140)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_78),
.Y(n_188)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g194 ( 
.A(n_79),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_17),
.B(n_11),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_17),
.B(n_11),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_85),
.B(n_98),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_86),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_55),
.Y(n_89)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_90),
.Y(n_181)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_92),
.Y(n_175)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_93),
.Y(n_195)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_29),
.B(n_11),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_29),
.A2(n_5),
.B(n_15),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_99),
.B(n_109),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_30),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_38),
.B(n_12),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_101),
.B(n_13),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_42),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_115),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_103),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_38),
.B(n_12),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_31),
.Y(n_113)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_30),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_116),
.A2(n_30),
.B1(n_42),
.B2(n_40),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_118),
.Y(n_134)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_120),
.Y(n_146)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_52),
.C(n_53),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_124),
.B(n_159),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_81),
.A2(n_34),
.B1(n_46),
.B2(n_48),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_126),
.A2(n_167),
.B1(n_171),
.B2(n_179),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_85),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_130),
.B(n_14),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_30),
.B1(n_46),
.B2(n_34),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_131),
.A2(n_158),
.B(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_98),
.A2(n_46),
.B1(n_34),
.B2(n_30),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_150),
.A2(n_187),
.B1(n_192),
.B2(n_1),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_13),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_113),
.A2(n_42),
.B1(n_51),
.B2(n_53),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_157),
.A2(n_89),
.B(n_75),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_61),
.A2(n_42),
.B1(n_35),
.B2(n_51),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_102),
.B(n_35),
.C(n_39),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_82),
.A2(n_18),
.B1(n_48),
.B2(n_45),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_111),
.A3(n_106),
.B1(n_104),
.B2(n_107),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_87),
.A2(n_43),
.B1(n_28),
.B2(n_45),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_88),
.A2(n_18),
.B1(n_28),
.B2(n_44),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_86),
.A2(n_39),
.B1(n_19),
.B2(n_44),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_90),
.A2(n_19),
.B1(n_43),
.B2(n_49),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_109),
.B(n_50),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_185),
.B(n_186),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_92),
.B(n_50),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g187 ( 
.A1(n_95),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_73),
.B(n_12),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_189),
.B(n_14),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_96),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_192)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_198),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_201),
.B(n_233),
.Y(n_279)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_151),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_202),
.Y(n_275)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_203),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_204),
.B(n_213),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_205),
.A2(n_138),
.B1(n_195),
.B2(n_149),
.Y(n_292)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_206),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_SL g207 ( 
.A(n_145),
.Y(n_207)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_207),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_208),
.Y(n_310)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_209),
.Y(n_283)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_210),
.Y(n_312)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_211),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_130),
.B(n_16),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_132),
.Y(n_214)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_153),
.Y(n_215)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_216),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_133),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_217),
.B(n_236),
.Y(n_296)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_134),
.Y(n_218)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_218),
.Y(n_300)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_219),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_165),
.A2(n_112),
.B1(n_59),
.B2(n_78),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_221),
.A2(n_247),
.B1(n_254),
.B2(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_223),
.Y(n_298)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_142),
.Y(n_224)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_224),
.Y(n_305)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_225),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_152),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_228),
.Y(n_268)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_142),
.Y(n_227)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_227),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_152),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_123),
.A2(n_116),
.B1(n_56),
.B2(n_62),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_229),
.Y(n_288)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_129),
.Y(n_230)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_230),
.Y(n_281)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_144),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_231),
.Y(n_289)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_232),
.Y(n_294)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_235),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_177),
.A2(n_70),
.B1(n_68),
.B2(n_64),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_237),
.A2(n_188),
.B1(n_193),
.B2(n_191),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_146),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_238),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_121),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_259),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_140),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_165),
.B(n_0),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_244),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_140),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_245),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_167),
.B(n_171),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_172),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_246),
.B(n_249),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_126),
.A2(n_63),
.B1(n_164),
.B2(n_169),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_181),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_248),
.A2(n_250),
.B1(n_255),
.B2(n_195),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_169),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_176),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_168),
.Y(n_251)
);

INVx13_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_164),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_253),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_137),
.B(n_1),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_181),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_155),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_258),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_187),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_166),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_141),
.Y(n_259)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_178),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_260),
.B(n_262),
.Y(n_318)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_141),
.Y(n_261)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_139),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_143),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_263),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_174),
.A2(n_4),
.B(n_179),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_264),
.A2(n_4),
.B(n_147),
.C(n_175),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_182),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_265),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_272),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_199),
.B(n_242),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_301),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_205),
.A2(n_158),
.B1(n_131),
.B2(n_127),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_290),
.A2(n_309),
.B1(n_197),
.B2(n_263),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_292),
.A2(n_311),
.B1(n_317),
.B2(n_232),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_199),
.B(n_238),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_244),
.B(n_149),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_304),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_200),
.B(n_135),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_254),
.A2(n_196),
.B1(n_160),
.B2(n_135),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_212),
.A2(n_161),
.B1(n_136),
.B2(n_128),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_315),
.Y(n_354)
);

XNOR2x1_ASAP7_75t_SL g349 ( 
.A(n_316),
.B(n_4),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_212),
.A2(n_188),
.B1(n_136),
.B2(n_196),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_304),
.A2(n_197),
.B1(n_257),
.B2(n_201),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_321),
.A2(n_328),
.B1(n_335),
.B2(n_347),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_287),
.B(n_220),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_322),
.B(n_348),
.Y(n_376)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_275),
.Y(n_323)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_323),
.Y(n_363)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_275),
.Y(n_325)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_325),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_326),
.A2(n_330),
.B1(n_341),
.B2(n_351),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_292),
.A2(n_261),
.B1(n_259),
.B2(n_191),
.Y(n_328)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_308),
.Y(n_329)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_329),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_274),
.A2(n_263),
.B1(n_215),
.B2(n_219),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_231),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_333),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_273),
.B(n_230),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_275),
.Y(n_334)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_280),
.Y(n_336)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_251),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_279),
.A2(n_240),
.B(n_239),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_339),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_340),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_274),
.A2(n_239),
.B1(n_211),
.B2(n_203),
.Y(n_341)
);

AO21x1_ASAP7_75t_L g342 ( 
.A1(n_279),
.A2(n_240),
.B(n_233),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_342),
.Y(n_397)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_305),
.Y(n_343)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_343),
.Y(n_394)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_344),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_288),
.A2(n_240),
.B1(n_209),
.B2(n_210),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_345),
.A2(n_308),
.B1(n_284),
.B2(n_267),
.Y(n_388)
);

OA22x2_ASAP7_75t_L g346 ( 
.A1(n_311),
.A2(n_216),
.B1(n_198),
.B2(n_227),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_357),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_273),
.A2(n_302),
.B1(n_301),
.B2(n_288),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_206),
.Y(n_348)
);

OAI21xp33_ASAP7_75t_L g375 ( 
.A1(n_349),
.A2(n_360),
.B(n_296),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_276),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_353),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_309),
.A2(n_260),
.B1(n_234),
.B2(n_224),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_268),
.A2(n_178),
.B1(n_193),
.B2(n_223),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_352),
.A2(n_358),
.B1(n_284),
.B2(n_280),
.Y(n_392)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_286),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_359),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_279),
.A2(n_303),
.B1(n_270),
.B2(n_313),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_356),
.A2(n_278),
.B1(n_313),
.B2(n_306),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_214),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_299),
.A2(n_250),
.B1(n_297),
.B2(n_318),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_277),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_307),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_362),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_278),
.B(n_306),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_333),
.B(n_296),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_366),
.B(n_370),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_326),
.A2(n_270),
.B1(n_300),
.B2(n_293),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_368),
.A2(n_379),
.B1(n_386),
.B2(n_328),
.Y(n_405)
);

OAI21xp33_ASAP7_75t_L g412 ( 
.A1(n_375),
.A2(n_366),
.B(n_369),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_332),
.B(n_282),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_384),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_291),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_382),
.C(n_383),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_327),
.A2(n_293),
.B1(n_283),
.B2(n_312),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_324),
.B(n_291),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_310),
.C(n_320),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_282),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_327),
.A2(n_312),
.B1(n_298),
.B2(n_319),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_358),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_396),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_388),
.A2(n_308),
.B1(n_294),
.B2(n_289),
.Y(n_431)
);

OAI21x1_ASAP7_75t_SL g403 ( 
.A1(n_392),
.A2(n_330),
.B(n_341),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_271),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_320),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_334),
.Y(n_419)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_399),
.Y(n_435)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_363),
.Y(n_400)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_400),
.Y(n_436)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_363),
.Y(n_402)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_402),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_403),
.A2(n_414),
.B(n_394),
.Y(n_454)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_372),
.Y(n_404)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_404),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_405),
.A2(n_422),
.B1(n_423),
.B2(n_425),
.Y(n_433)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_372),
.Y(n_406)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_406),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_339),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_407),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_385),
.A2(n_354),
.B(n_331),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_408),
.A2(n_412),
.B(n_380),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_398),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_409),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_369),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_410),
.B(n_416),
.Y(n_447)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_413),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_367),
.A2(n_354),
.B(n_331),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_389),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_381),
.A2(n_367),
.B1(n_387),
.B2(n_397),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_417),
.A2(n_420),
.B1(n_421),
.B2(n_426),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_396),
.A2(n_321),
.B(n_337),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_418),
.A2(n_371),
.B(n_295),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_419),
.B(n_429),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_381),
.A2(n_342),
.B1(n_351),
.B2(n_353),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_364),
.A2(n_342),
.B1(n_355),
.B2(n_349),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_368),
.A2(n_361),
.B1(n_346),
.B2(n_323),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_365),
.A2(n_346),
.B1(n_343),
.B2(n_359),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_424),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_365),
.A2(n_346),
.B1(n_325),
.B2(n_322),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_364),
.A2(n_340),
.B1(n_305),
.B2(n_319),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_379),
.A2(n_340),
.B1(n_336),
.B2(n_298),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_428),
.A2(n_430),
.B1(n_431),
.B2(n_393),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_376),
.B(n_289),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_386),
.A2(n_267),
.B1(n_344),
.B2(n_329),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_434),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_425),
.A2(n_376),
.B1(n_392),
.B2(n_373),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_437),
.A2(n_442),
.B1(n_446),
.B2(n_454),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_419),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_459),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_417),
.A2(n_416),
.B1(n_413),
.B2(n_420),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_R g471 ( 
.A(n_443),
.B(n_414),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_383),
.C(n_378),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_456),
.C(n_427),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_418),
.A2(n_390),
.B1(n_377),
.B2(n_394),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_415),
.B(n_382),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_450),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_411),
.B(n_390),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_391),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_451),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_410),
.B(n_374),
.Y(n_453)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_453),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_395),
.Y(n_455)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_455),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_399),
.B(n_374),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_411),
.A2(n_371),
.B1(n_395),
.B2(n_294),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_458),
.A2(n_426),
.B1(n_402),
.B2(n_400),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_407),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_460),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_407),
.B(n_295),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_421),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_465),
.B(n_451),
.C(n_408),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_461),
.Y(n_466)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_466),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_447),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_478),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_470),
.B(n_441),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_471),
.B(n_484),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_427),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_485),
.Y(n_490)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_447),
.Y(n_474)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_474),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_401),
.Y(n_475)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_475),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_401),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_476),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_409),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_477),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_406),
.Y(n_478)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_438),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_479),
.B(n_480),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_450),
.B(n_404),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_436),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_481),
.A2(n_488),
.B1(n_444),
.B2(n_449),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_443),
.B(n_422),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_423),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_487),
.Y(n_511)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_436),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_446),
.B(n_281),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_489),
.B(n_452),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_442),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_491),
.B(n_495),
.Y(n_519)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_493),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_469),
.B(n_465),
.C(n_473),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_505),
.C(n_512),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_470),
.B(n_462),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_497),
.B(n_498),
.Y(n_529)
);

FAx1_ASAP7_75t_SL g498 ( 
.A(n_476),
.B(n_438),
.CI(n_452),
.CON(n_498),
.SN(n_498)
);

A2O1A1Ixp33_ASAP7_75t_SL g500 ( 
.A1(n_474),
.A2(n_454),
.B(n_432),
.C(n_433),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_500),
.A2(n_487),
.B1(n_486),
.B2(n_463),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_441),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_504),
.B(n_405),
.C(n_481),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_468),
.B(n_460),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_472),
.A2(n_435),
.B1(n_457),
.B2(n_444),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_506),
.A2(n_510),
.B1(n_483),
.B2(n_486),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_464),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_472),
.A2(n_435),
.B1(n_432),
.B2(n_451),
.Y(n_510)
);

NOR2x1_ASAP7_75t_L g513 ( 
.A(n_503),
.B(n_475),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_513),
.A2(n_523),
.B(n_488),
.Y(n_539)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_516),
.Y(n_531)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_501),
.Y(n_517)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_517),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_499),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_518),
.B(n_520),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_510),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_521),
.A2(n_524),
.B1(n_431),
.B2(n_430),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_498),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_522),
.B(n_491),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_502),
.A2(n_485),
.B(n_477),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_512),
.A2(n_511),
.B1(n_509),
.B2(n_471),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_507),
.Y(n_525)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_525),
.Y(n_545)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_505),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_528),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_463),
.C(n_484),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_527),
.B(n_490),
.C(n_495),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_500),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_524),
.A2(n_496),
.B1(n_492),
.B2(n_500),
.Y(n_533)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_533),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_534),
.B(n_538),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_490),
.C(n_504),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_536),
.Y(n_556)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_537),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_528),
.B(n_502),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_539),
.A2(n_543),
.B(n_449),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_515),
.B(n_500),
.C(n_497),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_541),
.B(n_515),
.C(n_519),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_542),
.B(n_457),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_521),
.A2(n_530),
.B1(n_514),
.B2(n_529),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_544),
.A2(n_526),
.B1(n_514),
.B2(n_523),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_546),
.B(n_534),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_547),
.B(n_552),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_536),
.B(n_519),
.C(n_525),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_549),
.B(n_551),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_531),
.A2(n_513),
.B1(n_517),
.B2(n_428),
.Y(n_551)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_553),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_531),
.A2(n_403),
.B1(n_439),
.B2(n_424),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_554),
.B(n_543),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_539),
.A2(n_535),
.B(n_538),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_557),
.A2(n_541),
.B1(n_540),
.B2(n_532),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_551),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_558),
.B(n_563),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_555),
.B(n_532),
.Y(n_560)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_560),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_562),
.B(n_565),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_549),
.B(n_540),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_566),
.B(n_557),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_564),
.B(n_548),
.Y(n_570)
);

AOI21x1_ASAP7_75t_L g575 ( 
.A1(n_570),
.A2(n_553),
.B(n_561),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_571),
.B(n_572),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_560),
.A2(n_556),
.B(n_546),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_567),
.B(n_550),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_573),
.B(n_574),
.C(n_575),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_569),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_576),
.B(n_568),
.C(n_559),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_559),
.C(n_547),
.Y(n_579)
);

AOI322xp5_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_544),
.A3(n_577),
.B1(n_554),
.B2(n_545),
.C1(n_552),
.C2(n_542),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_580),
.A2(n_545),
.B(n_439),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_581),
.B(n_269),
.C(n_266),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_582),
.B(n_269),
.C(n_266),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_583),
.B(n_281),
.Y(n_584)
);


endmodule