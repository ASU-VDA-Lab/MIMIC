module fake_jpeg_17617_n_21 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_21);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_21;

wire n_13;
wire n_10;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

BUFx24_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

OR2x2_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_L g13 ( 
.A1(n_6),
.A2(n_0),
.B1(n_5),
.B2(n_4),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_13),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_17),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_3),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_10),
.B(n_4),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_11),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

AOI322xp5_ASAP7_75t_L g21 ( 
.A1(n_20),
.A2(n_9),
.A3(n_11),
.B1(n_14),
.B2(n_18),
.C1(n_17),
.C2(n_15),
.Y(n_21)
);


endmodule