module fake_jpeg_26314_n_322 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_7),
.B(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_18),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_38),
.B(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_55),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_25),
.B1(n_29),
.B2(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_61),
.B1(n_68),
.B2(n_77),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_62),
.Y(n_86)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_25),
.B1(n_34),
.B2(n_29),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_20),
.B1(n_23),
.B2(n_31),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_25),
.B1(n_29),
.B2(n_21),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_69),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_17),
.B1(n_30),
.B2(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_22),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_0),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_21),
.B1(n_18),
.B2(n_27),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_28),
.B(n_35),
.C(n_32),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_79),
.A2(n_33),
.B(n_9),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_81),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_48),
.B1(n_39),
.B2(n_21),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_75),
.B1(n_65),
.B2(n_50),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_32),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_84),
.B(n_9),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_47),
.C(n_41),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_22),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_92),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_22),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_111),
.B1(n_33),
.B2(n_1),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_107),
.Y(n_141)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_20),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_20),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_49),
.A2(n_36),
.B1(n_30),
.B2(n_31),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_23),
.B(n_33),
.C(n_35),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_0),
.B(n_1),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_23),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_110),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_75),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_67),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_57),
.A2(n_33),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_58),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_2),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_119),
.B1(n_136),
.B2(n_111),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_118),
.A2(n_125),
.B(n_129),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_78),
.A2(n_65),
.B1(n_50),
.B2(n_57),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_144),
.B1(n_112),
.B2(n_110),
.Y(n_155)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_2),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_132),
.B(n_145),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_88),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_139),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_101),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_115),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_84),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_91),
.A2(n_9),
.B1(n_13),
.B2(n_11),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_133),
.A2(n_104),
.B1(n_89),
.B2(n_113),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_90),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_148),
.B(n_149),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_92),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_153),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_161),
.B1(n_174),
.B2(n_176),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_123),
.A2(n_79),
.B1(n_106),
.B2(n_97),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_102),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_157),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_93),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_160),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_87),
.B1(n_80),
.B2(n_82),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_87),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_166),
.Y(n_203)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_99),
.Y(n_165)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_98),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_95),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_168),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_100),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_100),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_98),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_126),
.A2(n_82),
.B1(n_107),
.B2(n_109),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_143),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_126),
.A2(n_96),
.B1(n_81),
.B2(n_104),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_126),
.A2(n_10),
.B1(n_13),
.B2(n_6),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_129),
.B1(n_118),
.B2(n_120),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_131),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_180),
.B(n_185),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_142),
.C(n_135),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_182),
.C(n_207),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_149),
.C(n_159),
.Y(n_182)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_187),
.Y(n_228)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_118),
.Y(n_189)
);

A2O1A1O1Ixp25_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_193),
.B(n_154),
.C(n_147),
.D(n_171),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_152),
.A2(n_129),
.B1(n_119),
.B2(n_117),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_201),
.B1(n_161),
.B2(n_155),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_142),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_202),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_127),
.B1(n_125),
.B2(n_137),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_173),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_204),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_150),
.B(n_136),
.CI(n_145),
.CON(n_206),
.SN(n_206)
);

XOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_137),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_127),
.C(n_143),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_192),
.B1(n_202),
.B2(n_184),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_200),
.B(n_147),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_195),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_158),
.B1(n_157),
.B2(n_175),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_213),
.A2(n_191),
.B1(n_185),
.B2(n_189),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_196),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_216),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_177),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_170),
.B(n_178),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_217),
.A2(n_221),
.B(n_222),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_201),
.B(n_170),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_188),
.A2(n_137),
.B(n_130),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_224),
.B(n_230),
.Y(n_242)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_10),
.B(n_6),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_229),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_130),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_194),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_232),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_184),
.A2(n_173),
.B1(n_6),
.B2(n_8),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_190),
.B1(n_187),
.B2(n_206),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_188),
.A2(n_4),
.B(n_5),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_234),
.A2(n_224),
.B(n_207),
.C(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_182),
.C(n_181),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_245),
.C(n_231),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_248),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_217),
.B(n_234),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_192),
.C(n_197),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_249),
.B1(n_210),
.B2(n_233),
.Y(n_265)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_190),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_255),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_213),
.B(n_193),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_223),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_256),
.Y(n_259)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_242),
.B(n_230),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_263),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_261),
.A2(n_244),
.B(n_241),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_222),
.C(n_215),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_269),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_242),
.B(n_221),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_271),
.C(n_244),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_273),
.B1(n_252),
.B2(n_243),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_216),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_225),
.C(n_199),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

AO22x1_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_206),
.B1(n_199),
.B2(n_220),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_280),
.C(n_285),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_239),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_283),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_239),
.B(n_243),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_278),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_253),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_284),
.B(n_274),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_244),
.C(n_257),
.Y(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_265),
.A2(n_251),
.B1(n_246),
.B2(n_253),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_240),
.C(n_248),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_267),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_279),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_289),
.B(n_291),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_259),
.Y(n_291)
);

AO221x1_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_229),
.B1(n_232),
.B2(n_211),
.C(n_273),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_294),
.B(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_228),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_295),
.B1(n_290),
.B2(n_179),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_290),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_297),
.A2(n_299),
.B(n_296),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_300),
.B(n_301),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_276),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_280),
.B1(n_273),
.B2(n_263),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_262),
.C(n_281),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_275),
.C(n_11),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_179),
.B1(n_269),
.B2(n_277),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_310),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_4),
.A3(n_5),
.B1(n_11),
.B2(n_16),
.C1(n_275),
.C2(n_305),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_313),
.B(n_302),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_312),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_311),
.B(n_303),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_301),
.C(n_308),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_318),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_308),
.B(n_5),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_5),
.Y(n_322)
);


endmodule