module real_aes_5650_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_552;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_922;
wire n_482;
wire n_520;
wire n_633;
wire n_926;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_0), .A2(n_225), .B1(n_305), .B2(n_311), .Y(n_614) );
AO22x2_ASAP7_75t_L g595 ( .A1(n_1), .A2(n_596), .B1(n_616), .B2(n_617), .Y(n_595) );
INVxp67_ASAP7_75t_SL g616 ( .A(n_1), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_2), .A2(n_56), .B1(n_360), .B2(n_370), .Y(n_634) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_3), .Y(n_644) );
AND2x4_ASAP7_75t_L g658 ( .A(n_3), .B(n_659), .Y(n_658) );
AND2x4_ASAP7_75t_L g667 ( .A(n_3), .B(n_241), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_4), .A2(n_110), .B1(n_670), .B2(n_683), .Y(n_701) );
INVx1_ASAP7_75t_L g515 ( .A(n_5), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_6), .A2(n_187), .B1(n_370), .B2(n_372), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_7), .A2(n_213), .B1(n_366), .B2(n_368), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_8), .A2(n_84), .B1(n_305), .B2(n_311), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_9), .A2(n_13), .B1(n_491), .B2(n_492), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_10), .A2(n_15), .B1(n_353), .B2(n_355), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_11), .A2(n_194), .B1(n_353), .B2(n_503), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_12), .A2(n_70), .B1(n_462), .B2(n_500), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_14), .A2(n_103), .B1(n_457), .B2(n_459), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_16), .A2(n_73), .B1(n_362), .B2(n_470), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_17), .A2(n_202), .B1(n_428), .B2(n_429), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_18), .A2(n_111), .B1(n_491), .B2(n_492), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_19), .A2(n_106), .B1(n_585), .B2(n_586), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_20), .Y(n_668) );
AO22x2_ASAP7_75t_L g682 ( .A1(n_21), .A2(n_66), .B1(n_670), .B2(n_683), .Y(n_682) );
AO22x1_ASAP7_75t_L g684 ( .A1(n_22), .A2(n_248), .B1(n_685), .B2(n_687), .Y(n_684) );
INVxp33_ASAP7_75t_SL g719 ( .A(n_23), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_24), .A2(n_102), .B1(n_888), .B2(n_890), .Y(n_887) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_25), .A2(n_30), .B1(n_509), .B2(n_510), .C(n_513), .Y(n_508) );
INVx1_ASAP7_75t_L g528 ( .A(n_26), .Y(n_528) );
INVx1_ASAP7_75t_L g909 ( .A(n_27), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_28), .A2(n_95), .B1(n_387), .B2(n_435), .Y(n_917) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_29), .A2(n_328), .B(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_31), .A2(n_125), .B1(n_328), .B2(n_330), .Y(n_327) );
XNOR2x1_ASAP7_75t_L g520 ( .A(n_32), .B(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_32), .A2(n_105), .B1(n_666), .B2(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_33), .A2(n_156), .B1(n_461), .B2(n_463), .Y(n_460) );
INVx1_ASAP7_75t_L g628 ( .A(n_34), .Y(n_628) );
INVx1_ASAP7_75t_L g280 ( .A(n_35), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_35), .B(n_183), .Y(n_295) );
INVxp67_ASAP7_75t_L g339 ( .A(n_35), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_36), .A2(n_137), .B1(n_409), .B2(n_470), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_37), .A2(n_75), .B1(n_424), .B2(n_429), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_38), .A2(n_196), .B1(n_660), .B2(n_670), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_39), .A2(n_91), .B1(n_360), .B2(n_362), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_40), .A2(n_113), .B1(n_414), .B2(n_466), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_41), .A2(n_109), .B1(n_685), .B2(n_692), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_42), .A2(n_128), .B1(n_362), .B2(n_462), .Y(n_879) );
XNOR2x1_ASAP7_75t_L g430 ( .A(n_43), .B(n_431), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_44), .A2(n_67), .B1(n_324), .B2(n_325), .Y(n_323) );
XNOR2x1_ASAP7_75t_L g400 ( .A(n_45), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_46), .B(n_265), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_47), .A2(n_79), .B1(n_576), .B2(n_577), .Y(n_575) );
AOI21xp33_ASAP7_75t_SL g598 ( .A1(n_48), .A2(n_550), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g288 ( .A(n_49), .Y(n_288) );
INVx1_ASAP7_75t_L g564 ( .A(n_50), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_51), .A2(n_233), .B1(n_330), .B2(n_333), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_52), .A2(n_148), .B1(n_424), .B2(n_590), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_53), .A2(n_206), .B1(n_411), .B2(n_412), .Y(n_410) );
BUFx2_ASAP7_75t_L g604 ( .A(n_54), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_55), .A2(n_89), .B1(n_491), .B2(n_492), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_57), .A2(n_216), .B1(n_683), .B2(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g514 ( .A(n_58), .Y(n_514) );
INVx2_ASAP7_75t_L g642 ( .A(n_59), .Y(n_642) );
INVxp33_ASAP7_75t_SL g671 ( .A(n_60), .Y(n_671) );
XNOR2x1_ASAP7_75t_L g872 ( .A(n_60), .B(n_873), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_60), .A2(n_901), .B1(n_922), .B2(n_924), .Y(n_900) );
INVx1_ASAP7_75t_L g657 ( .A(n_61), .Y(n_657) );
AND2x4_ASAP7_75t_L g663 ( .A(n_61), .B(n_642), .Y(n_663) );
INVx1_ASAP7_75t_SL g686 ( .A(n_61), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_62), .A2(n_217), .B1(n_424), .B2(n_550), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_63), .A2(n_902), .B1(n_903), .B2(n_904), .Y(n_901) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_63), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_64), .A2(n_135), .B1(n_424), .B2(n_585), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_65), .A2(n_165), .B1(n_316), .B2(n_320), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_68), .B(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_69), .A2(n_145), .B1(n_378), .B2(n_552), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g369 ( .A1(n_71), .A2(n_228), .B1(n_370), .B2(n_372), .Y(n_369) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_72), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_74), .A2(n_185), .B1(n_341), .B2(n_342), .Y(n_493) );
INVx1_ASAP7_75t_L g543 ( .A(n_76), .Y(n_543) );
INVx1_ASAP7_75t_L g560 ( .A(n_77), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_78), .A2(n_161), .B1(n_467), .B2(n_579), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_80), .A2(n_626), .B(n_627), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_81), .A2(n_119), .B1(n_370), .B2(n_876), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_82), .A2(n_112), .B1(n_893), .B2(n_894), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_83), .A2(n_195), .B1(n_384), .B2(n_387), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_85), .A2(n_133), .B1(n_429), .B2(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g266 ( .A(n_86), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_86), .B(n_182), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_87), .A2(n_132), .B1(n_372), .B2(n_404), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_88), .A2(n_152), .B1(n_404), .B2(n_405), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_90), .A2(n_126), .B1(n_670), .B2(n_683), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_92), .A2(n_192), .B1(n_328), .B2(n_332), .Y(n_483) );
AO221x2_ASAP7_75t_L g652 ( .A1(n_93), .A2(n_94), .B1(n_653), .B2(n_660), .C(n_664), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_96), .A2(n_244), .B1(n_655), .B2(n_683), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_97), .A2(n_160), .B1(n_392), .B2(n_395), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_98), .B(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g349 ( .A(n_99), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_100), .A2(n_188), .B1(n_368), .B2(n_372), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_101), .A2(n_243), .B1(n_324), .B2(n_325), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_104), .A2(n_116), .B1(n_434), .B2(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g451 ( .A(n_107), .Y(n_451) );
INVx1_ASAP7_75t_L g600 ( .A(n_108), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_114), .A2(n_229), .B1(n_305), .B2(n_311), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_115), .A2(n_214), .B1(n_341), .B2(n_342), .Y(n_554) );
INVx1_ASAP7_75t_L g530 ( .A(n_117), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_118), .A2(n_175), .B1(n_405), .B2(n_539), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_120), .A2(n_138), .B1(n_408), .B2(n_409), .Y(n_407) );
XOR2x2_ASAP7_75t_L g256 ( .A(n_121), .B(n_257), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_121), .A2(n_186), .B1(n_685), .B2(n_692), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_122), .A2(n_212), .B1(n_330), .B2(n_423), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_123), .A2(n_124), .B1(n_429), .B2(n_916), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_127), .A2(n_129), .B1(n_412), .B2(n_470), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_130), .A2(n_155), .B1(n_525), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_131), .A2(n_169), .B1(n_423), .B2(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g419 ( .A(n_134), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_136), .A2(n_164), .B1(n_469), .B2(n_471), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_139), .A2(n_220), .B1(n_408), .B2(n_458), .Y(n_877) );
INVx1_ASAP7_75t_L g478 ( .A(n_140), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_141), .A2(n_231), .B1(n_414), .B2(n_415), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_142), .A2(n_191), .B1(n_411), .B2(n_464), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_143), .B(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_144), .A2(n_172), .B1(n_655), .B2(n_666), .Y(n_679) );
XOR2xp5_ASAP7_75t_L g618 ( .A(n_146), .B(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_147), .A2(n_167), .B1(n_438), .B2(n_440), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g913 ( .A1(n_149), .A2(n_222), .B1(n_370), .B2(n_462), .Y(n_913) );
INVx1_ASAP7_75t_L g884 ( .A(n_150), .Y(n_884) );
OA22x2_ASAP7_75t_L g270 ( .A1(n_151), .A2(n_183), .B1(n_265), .B2(n_269), .Y(n_270) );
INVx1_ASAP7_75t_L g302 ( .A(n_151), .Y(n_302) );
AOI21xp33_ASAP7_75t_L g442 ( .A1(n_153), .A2(n_443), .B(n_448), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_154), .A2(n_246), .B1(n_372), .B2(n_539), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_157), .A2(n_205), .B1(n_414), .B2(n_503), .Y(n_502) );
XOR2x2_ASAP7_75t_L g570 ( .A(n_158), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g454 ( .A(n_159), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_162), .A2(n_239), .B1(n_414), .B2(n_503), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_163), .A2(n_166), .B1(n_341), .B2(n_342), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_168), .A2(n_230), .B1(n_305), .B2(n_311), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_170), .A2(n_207), .B1(n_439), .B2(n_450), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_171), .A2(n_181), .B1(n_324), .B2(n_325), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_173), .A2(n_204), .B1(n_332), .B2(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g714 ( .A(n_174), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_176), .A2(n_235), .B1(n_470), .B2(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g565 ( .A(n_177), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_177), .A2(n_197), .B1(n_655), .B2(n_687), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_178), .B(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g608 ( .A(n_179), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_180), .A2(n_211), .B1(n_341), .B2(n_342), .Y(n_615) );
INVx1_ASAP7_75t_L g282 ( .A(n_182), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_182), .B(n_299), .Y(n_298) );
OAI21xp33_ASAP7_75t_L g313 ( .A1(n_183), .A2(n_201), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_184), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g526 ( .A(n_189), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_190), .A2(n_232), .B1(n_324), .B2(n_325), .Y(n_489) );
INVx1_ASAP7_75t_L g381 ( .A(n_193), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_198), .A2(n_242), .B1(n_259), .B2(n_283), .C(n_287), .Y(n_258) );
INVx1_ASAP7_75t_SL g715 ( .A(n_199), .Y(n_715) );
AOI221x1_ASAP7_75t_SL g906 ( .A1(n_200), .A2(n_210), .B1(n_378), .B2(n_907), .C(n_908), .Y(n_906) );
INVx1_ASAP7_75t_L g268 ( .A(n_201), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_201), .B(n_234), .Y(n_296) );
AOI21xp33_ASAP7_75t_L g377 ( .A1(n_203), .A2(n_378), .B(n_380), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g540 ( .A1(n_208), .A2(n_238), .B1(n_509), .B2(n_541), .C(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_209), .A2(n_512), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g487 ( .A(n_215), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g881 ( .A1(n_218), .A2(n_882), .B(n_883), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_219), .A2(n_237), .B1(n_414), .B2(n_503), .Y(n_919) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_221), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g485 ( .A1(n_223), .A2(n_284), .B(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_224), .A2(n_227), .B1(n_366), .B2(n_458), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_226), .A2(n_588), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_234), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_236), .B(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_240), .B(n_450), .Y(n_532) );
INVx1_ASAP7_75t_L g659 ( .A(n_241), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_245), .A2(n_247), .B1(n_353), .B2(n_503), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_645), .B(n_648), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_473), .B(n_637), .Y(n_250) );
INVx1_ASAP7_75t_L g647 ( .A(n_251), .Y(n_647) );
XNOR2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_343), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND3x1_ASAP7_75t_L g257 ( .A(n_258), .B(n_303), .C(n_322), .Y(n_257) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_259), .Y(n_390) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g426 ( .A(n_260), .Y(n_426) );
INVx2_ASAP7_75t_L g882 ( .A(n_260), .Y(n_882) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g447 ( .A(n_261), .Y(n_447) );
BUFx3_ASAP7_75t_L g588 ( .A(n_261), .Y(n_588) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_271), .Y(n_261) );
AND2x4_ASAP7_75t_L g317 ( .A(n_262), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g321 ( .A(n_262), .B(n_308), .Y(n_321) );
AND2x4_ASAP7_75t_L g332 ( .A(n_262), .B(n_329), .Y(n_332) );
AND2x2_ASAP7_75t_L g367 ( .A(n_262), .B(n_308), .Y(n_367) );
AND2x2_ASAP7_75t_L g398 ( .A(n_262), .B(n_329), .Y(n_398) );
AND2x4_ASAP7_75t_L g491 ( .A(n_262), .B(n_308), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_262), .B(n_326), .Y(n_492) );
AND2x2_ASAP7_75t_L g512 ( .A(n_262), .B(n_271), .Y(n_512) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_270), .Y(n_262) );
INVx1_ASAP7_75t_L g286 ( .A(n_263), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
NAND2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g269 ( .A(n_265), .Y(n_269) );
INVx3_ASAP7_75t_L g275 ( .A(n_265), .Y(n_275) );
NAND2xp33_ASAP7_75t_L g281 ( .A(n_265), .B(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_265), .Y(n_293) );
INVx1_ASAP7_75t_L g314 ( .A(n_265), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_266), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g338 ( .A1(n_268), .A2(n_314), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g285 ( .A(n_270), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g307 ( .A(n_270), .Y(n_307) );
AND2x2_ASAP7_75t_L g337 ( .A(n_270), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g284 ( .A(n_271), .B(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g330 ( .A(n_271), .B(n_312), .Y(n_330) );
AND2x4_ASAP7_75t_L g342 ( .A(n_271), .B(n_306), .Y(n_342) );
AND2x2_ASAP7_75t_L g358 ( .A(n_271), .B(n_306), .Y(n_358) );
AND2x4_ASAP7_75t_L g386 ( .A(n_271), .B(n_285), .Y(n_386) );
AND2x4_ASAP7_75t_L g388 ( .A(n_271), .B(n_312), .Y(n_388) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_277), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_L g308 ( .A(n_273), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g319 ( .A(n_273), .B(n_310), .Y(n_319) );
AND2x4_ASAP7_75t_L g329 ( .A(n_273), .B(n_277), .Y(n_329) );
AND2x2_ASAP7_75t_L g334 ( .A(n_273), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_275), .B(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_L g299 ( .A(n_275), .Y(n_299) );
NAND3xp33_ASAP7_75t_L g297 ( .A(n_276), .B(n_298), .C(n_300), .Y(n_297) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g310 ( .A(n_278), .Y(n_310) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g328 ( .A(n_285), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g379 ( .A(n_285), .B(n_329), .Y(n_379) );
AND2x4_ASAP7_75t_L g306 ( .A(n_286), .B(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_289), .B(n_487), .Y(n_486) );
INVx4_ASAP7_75t_L g545 ( .A(n_289), .Y(n_545) );
INVx4_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx3_ASAP7_75t_L g382 ( .A(n_290), .Y(n_382) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_291), .Y(n_421) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_294), .B(n_297), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_293), .B(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_294), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_299), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g312 ( .A(n_300), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_315), .Y(n_303) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
AND2x4_ASAP7_75t_L g324 ( .A(n_306), .B(n_318), .Y(n_324) );
AND2x4_ASAP7_75t_L g341 ( .A(n_306), .B(n_329), .Y(n_341) );
AND2x4_ASAP7_75t_L g354 ( .A(n_306), .B(n_329), .Y(n_354) );
AND2x4_ASAP7_75t_L g361 ( .A(n_306), .B(n_308), .Y(n_361) );
AND2x4_ASAP7_75t_L g371 ( .A(n_306), .B(n_326), .Y(n_371) );
AND2x4_ASAP7_75t_L g311 ( .A(n_308), .B(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g364 ( .A(n_308), .B(n_312), .Y(n_364) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g325 ( .A(n_312), .B(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g373 ( .A(n_312), .B(n_326), .Y(n_373) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx3_ASAP7_75t_L g368 ( .A(n_317), .Y(n_368) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_317), .Y(n_409) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_317), .Y(n_458) );
BUFx12f_ASAP7_75t_L g539 ( .A(n_317), .Y(n_539) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g326 ( .A(n_319), .Y(n_326) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx4f_ASAP7_75t_L g408 ( .A(n_321), .Y(n_408) );
AND4x1_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .C(n_331), .D(n_340), .Y(n_322) );
INVx2_ASAP7_75t_L g609 ( .A(n_332), .Y(n_609) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_337), .Y(n_333) );
AND2x4_ASAP7_75t_L g394 ( .A(n_334), .B(n_337), .Y(n_394) );
AND2x4_ASAP7_75t_L g606 ( .A(n_334), .B(n_337), .Y(n_606) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
XNOR2x1_ASAP7_75t_L g345 ( .A(n_346), .B(n_430), .Y(n_345) );
AO22x2_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_399), .B2(n_400), .Y(n_346) );
INVx2_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
XNOR2x1_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
NOR2x1_ASAP7_75t_L g350 ( .A(n_351), .B(n_374), .Y(n_350) );
NAND4xp25_ASAP7_75t_L g351 ( .A(n_352), .B(n_359), .C(n_365), .D(n_369), .Y(n_351) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx12f_ASAP7_75t_L g414 ( .A(n_354), .Y(n_414) );
INVx3_ASAP7_75t_L g581 ( .A(n_354), .Y(n_581) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx3_ASAP7_75t_L g415 ( .A(n_358), .Y(n_415) );
BUFx5_ASAP7_75t_L g467 ( .A(n_358), .Y(n_467) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_358), .Y(n_503) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx12f_ASAP7_75t_L g411 ( .A(n_361), .Y(n_411) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_361), .Y(n_462) );
INVx4_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g412 ( .A(n_363), .Y(n_412) );
INVx1_ASAP7_75t_L g472 ( .A(n_363), .Y(n_472) );
INVx4_ASAP7_75t_L g500 ( .A(n_363), .Y(n_500) );
INVx1_ASAP7_75t_L g577 ( .A(n_363), .Y(n_577) );
INVx2_ASAP7_75t_L g921 ( .A(n_363), .Y(n_921) );
INVx8_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx8_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_367), .Y(n_470) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_371), .Y(n_404) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_371), .Y(n_464) );
BUFx3_ASAP7_75t_L g459 ( .A(n_372), .Y(n_459) );
BUFx12f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx6_ASAP7_75t_L g406 ( .A(n_373), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_389), .C(n_391), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_383), .Y(n_376) );
INVx4_ASAP7_75t_L g531 ( .A(n_378), .Y(n_531) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx3_ASAP7_75t_L g439 ( .A(n_379), .Y(n_439) );
BUFx3_ASAP7_75t_L g550 ( .A(n_379), .Y(n_550) );
INVx1_ASAP7_75t_L g623 ( .A(n_379), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx4_ASAP7_75t_L g453 ( .A(n_382), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_382), .B(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_382), .B(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_382), .B(n_600), .Y(n_599) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g585 ( .A(n_385), .Y(n_585) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
BUFx8_ASAP7_75t_SL g435 ( .A(n_386), .Y(n_435) );
BUFx3_ASAP7_75t_L g509 ( .A(n_386), .Y(n_509) );
INVx2_ASAP7_75t_L g889 ( .A(n_386), .Y(n_889) );
BUFx3_ASAP7_75t_L g436 ( .A(n_387), .Y(n_436) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_388), .Y(n_424) );
INVx3_ASAP7_75t_L g891 ( .A(n_388), .Y(n_891) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g552 ( .A(n_393), .Y(n_552) );
INVx2_ASAP7_75t_L g916 ( .A(n_393), .Y(n_916) );
INVx5_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
BUFx4f_ASAP7_75t_L g450 ( .A(n_394), .Y(n_450) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g590 ( .A(n_396), .Y(n_590) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g894 ( .A(n_397), .Y(n_894) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx3_ASAP7_75t_L g429 ( .A(n_398), .Y(n_429) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_398), .Y(n_525) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
NOR2x1_ASAP7_75t_L g401 ( .A(n_402), .B(n_416), .Y(n_401) );
NAND4xp25_ASAP7_75t_L g402 ( .A(n_403), .B(n_407), .C(n_410), .D(n_413), .Y(n_402) );
INVx5_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g876 ( .A(n_406), .Y(n_876) );
BUFx12f_ASAP7_75t_L g576 ( .A(n_411), .Y(n_576) );
NAND4xp25_ASAP7_75t_SL g416 ( .A(n_417), .B(n_422), .C(n_425), .D(n_427), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_SL g592 ( .A(n_421), .Y(n_592) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_421), .Y(n_631) );
INVx3_ASAP7_75t_L g527 ( .A(n_424), .Y(n_527) );
INVx2_ASAP7_75t_L g441 ( .A(n_429), .Y(n_441) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_455), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_437), .C(n_442), .Y(n_432) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g561 ( .A(n_435), .Y(n_561) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g541 ( .A(n_446), .Y(n_541) );
INVx1_ASAP7_75t_L g907 ( .A(n_446), .Y(n_907) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g482 ( .A(n_447), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_451), .B1(n_452), .B2(n_454), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND4xp25_ASAP7_75t_SL g455 ( .A(n_456), .B(n_460), .C(n_465), .D(n_468), .Y(n_455) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g646 ( .A(n_473), .Y(n_646) );
XNOR2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_567), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_516), .B1(n_517), .B2(n_566), .Y(n_474) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_475), .Y(n_566) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
XNOR2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_495), .Y(n_476) );
XNOR2x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
OR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_488), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g480 ( .A(n_481), .B(n_483), .C(n_484), .D(n_485), .Y(n_480) );
BUFx3_ASAP7_75t_L g626 ( .A(n_482), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .C(n_493), .D(n_494), .Y(n_488) );
XNOR2x1_ASAP7_75t_L g495 ( .A(n_496), .B(n_515), .Y(n_495) );
NAND4xp75_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .C(n_505), .D(n_508), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
XNOR2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_546), .Y(n_519) );
NAND4xp75_ASAP7_75t_L g521 ( .A(n_522), .B(n_533), .C(n_536), .D(n_540), .Y(n_521) );
NOR2xp67_ASAP7_75t_L g522 ( .A(n_523), .B(n_529), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_526), .B1(n_527), .B2(n_528), .Y(n_523) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_532), .Y(n_529) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
XOR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_565), .Y(n_546) );
NOR4xp75_ASAP7_75t_L g547 ( .A(n_548), .B(n_553), .C(n_556), .D(n_559), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OAI21x1_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_561), .B(n_562), .Y(n_559) );
XOR2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_593), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_572), .B(n_582), .Y(n_571) );
NAND4xp25_ASAP7_75t_SL g572 ( .A(n_573), .B(n_574), .C(n_575), .D(n_578), .Y(n_572) );
BUFx4f_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND4xp25_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .C(n_589), .D(n_591), .Y(n_582) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_SL g910 ( .A(n_592), .Y(n_910) );
BUFx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
XNOR2xp5_ASAP7_75t_SL g594 ( .A(n_595), .B(n_618), .Y(n_594) );
INVx1_ASAP7_75t_L g617 ( .A(n_596), .Y(n_617) );
NOR2x1_ASAP7_75t_L g596 ( .A(n_597), .B(n_611), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .C(n_610), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_605), .B1(n_607), .B2(n_609), .Y(n_602) );
CKINVDCx16_ASAP7_75t_R g603 ( .A(n_604), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g627 ( .A1(n_605), .A2(n_628), .B(n_629), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g883 ( .A1(n_605), .A2(n_884), .B(n_885), .Y(n_883) );
INVx4_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
CKINVDCx9p33_ASAP7_75t_R g607 ( .A(n_608), .Y(n_607) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .C(n_614), .D(n_615), .Y(n_611) );
NOR2x1_ASAP7_75t_SL g619 ( .A(n_620), .B(n_632), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .C(n_625), .Y(n_620) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g893 ( .A(n_623), .Y(n_893) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g886 ( .A(n_631), .Y(n_886) );
NAND4xp25_ASAP7_75t_SL g632 ( .A(n_633), .B(n_634), .C(n_635), .D(n_636), .Y(n_632) );
BUFx10_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_643), .C(n_644), .Y(n_639) );
AND2x2_ASAP7_75t_L g897 ( .A(n_640), .B(n_898), .Y(n_897) );
AND2x2_ASAP7_75t_L g923 ( .A(n_640), .B(n_899), .Y(n_923) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OA21x2_ASAP7_75t_L g925 ( .A1(n_641), .A2(n_686), .B(n_926), .Y(n_925) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g656 ( .A(n_642), .B(n_657), .Y(n_656) );
AND3x4_ASAP7_75t_L g685 ( .A(n_642), .B(n_658), .C(n_686), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_643), .B(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_644), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
OAI221xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_868), .B1(n_870), .B2(n_895), .C(n_900), .Y(n_648) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_828), .C(n_844), .Y(n_649) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_672), .B(n_775), .C(n_801), .Y(n_650) );
HB1xp67_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_652), .B(n_785), .Y(n_784) );
AOI211xp5_ASAP7_75t_L g801 ( .A1(n_652), .A2(n_802), .B(n_806), .C(n_818), .Y(n_801) );
INVx2_ASAP7_75t_L g829 ( .A(n_652), .Y(n_829) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_654), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_716) );
INVx3_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
AND2x4_ASAP7_75t_L g666 ( .A(n_656), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g687 ( .A(n_656), .B(n_667), .Y(n_687) );
AND2x2_ASAP7_75t_L g692 ( .A(n_656), .B(n_667), .Y(n_692) );
AND2x4_ASAP7_75t_L g662 ( .A(n_658), .B(n_663), .Y(n_662) );
AND2x4_ASAP7_75t_L g683 ( .A(n_658), .B(n_663), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_658), .B(n_663), .Y(n_718) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_L g670 ( .A(n_663), .B(n_667), .Y(n_670) );
AND2x2_ASAP7_75t_L g690 ( .A(n_663), .B(n_667), .Y(n_690) );
AND2x2_ASAP7_75t_L g707 ( .A(n_663), .B(n_667), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B1(n_669), .B2(n_671), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_665), .A2(n_669), .B1(n_714), .B2(n_715), .Y(n_713) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_667), .Y(n_926) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g869 ( .A(n_670), .Y(n_869) );
NOR4xp25_ASAP7_75t_SL g672 ( .A(n_673), .B(n_729), .C(n_737), .D(n_755), .Y(n_672) );
OAI322xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_693), .A3(n_703), .B1(n_709), .B2(n_722), .C1(n_723), .C2(n_725), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_680), .Y(n_674) );
INVx5_ASAP7_75t_L g730 ( .A(n_675), .Y(n_730) );
INVx3_ASAP7_75t_L g740 ( .A(n_675), .Y(n_740) );
AOI32xp33_ASAP7_75t_L g766 ( .A1(n_675), .A2(n_767), .A3(n_769), .B1(n_771), .B2(n_773), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_675), .B(n_711), .Y(n_817) );
INVx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g758 ( .A(n_676), .B(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g774 ( .A(n_676), .B(n_681), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_676), .B(n_722), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_676), .B(n_756), .Y(n_835) );
AND2x2_ASAP7_75t_L g862 ( .A(n_676), .B(n_727), .Y(n_862) );
INVx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g726 ( .A(n_677), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g754 ( .A(n_677), .B(n_747), .Y(n_754) );
OR2x2_ASAP7_75t_L g796 ( .A(n_677), .B(n_797), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx2_ASAP7_75t_L g797 ( .A(n_680), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_680), .B(n_712), .Y(n_867) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_688), .Y(n_680) );
CKINVDCx6p67_ASAP7_75t_R g722 ( .A(n_681), .Y(n_722) );
INVx1_ASAP7_75t_L g728 ( .A(n_681), .Y(n_728) );
OR2x2_ASAP7_75t_L g747 ( .A(n_681), .B(n_688), .Y(n_747) );
AND2x2_ASAP7_75t_L g810 ( .A(n_681), .B(n_743), .Y(n_810) );
OR2x6_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g743 ( .A(n_688), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_688), .B(n_733), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_688), .B(n_712), .Y(n_772) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_688), .Y(n_780) );
BUFx2_ASAP7_75t_L g786 ( .A(n_688), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_688), .B(n_712), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_688), .B(n_774), .Y(n_838) );
AND2x4_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_702), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_694), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g724 ( .A(n_695), .B(n_703), .Y(n_724) );
AND2x2_ASAP7_75t_L g856 ( .A(n_695), .B(n_735), .Y(n_856) );
AND2x2_ASAP7_75t_L g858 ( .A(n_695), .B(n_859), .Y(n_858) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_699), .Y(n_695) );
OR2x2_ASAP7_75t_L g702 ( .A(n_696), .B(n_699), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_696), .Y(n_721) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
OR2x2_ASAP7_75t_L g720 ( .A(n_699), .B(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_699), .B(n_703), .Y(n_748) );
OR2x2_ASAP7_75t_L g770 ( .A(n_699), .B(n_705), .Y(n_770) );
AND2x2_ASAP7_75t_L g790 ( .A(n_699), .B(n_721), .Y(n_790) );
INVx1_ASAP7_75t_L g805 ( .A(n_699), .Y(n_805) );
AND2x2_ASAP7_75t_L g815 ( .A(n_699), .B(n_789), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_699), .B(n_735), .Y(n_865) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g736 ( .A(n_702), .Y(n_736) );
OR2x2_ASAP7_75t_L g756 ( .A(n_702), .B(n_735), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_702), .B(n_782), .Y(n_781) );
OAI322xp33_ASAP7_75t_L g833 ( .A1(n_702), .A2(n_711), .A3(n_725), .B1(n_742), .B2(n_751), .C1(n_774), .C2(n_834), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_702), .B(n_733), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_703), .B(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_703), .B(n_721), .Y(n_765) );
AND2x2_ASAP7_75t_L g794 ( .A(n_703), .B(n_790), .Y(n_794) );
INVx3_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx3_ASAP7_75t_L g735 ( .A(n_705), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_705), .B(n_733), .Y(n_782) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_720), .Y(n_710) );
INVx1_ASAP7_75t_L g792 ( .A(n_711), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g803 ( .A(n_711), .B(n_785), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_711), .B(n_770), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_711), .B(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx3_ASAP7_75t_L g733 ( .A(n_712), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_712), .B(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_712), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_712), .B(n_735), .Y(n_821) );
OR2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g752 ( .A(n_720), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_720), .B(n_735), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_720), .B(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_721), .B(n_827), .Y(n_834) );
AOI221xp5_ASAP7_75t_L g852 ( .A1(n_721), .A2(n_741), .B1(n_752), .B2(n_810), .C(n_853), .Y(n_852) );
AND2x2_ASAP7_75t_L g785 ( .A(n_722), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g851 ( .A(n_722), .Y(n_851) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g791 ( .A(n_724), .B(n_726), .C(n_792), .Y(n_791) );
OAI21xp5_ASAP7_75t_SL g824 ( .A1(n_724), .A2(n_734), .B(n_825), .Y(n_824) );
AOI221xp5_ASAP7_75t_L g845 ( .A1(n_724), .A2(n_734), .B1(n_841), .B2(n_846), .C(n_847), .Y(n_845) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_726), .B(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_727), .B(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
CKINVDCx14_ASAP7_75t_R g854 ( .A(n_730), .Y(n_854) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
AND2x2_ASAP7_75t_L g745 ( .A(n_733), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g800 ( .A(n_733), .B(n_790), .Y(n_800) );
INVx1_ASAP7_75t_SL g849 ( .A(n_733), .Y(n_849) );
AND2x2_ASAP7_75t_L g808 ( .A(n_734), .B(n_792), .Y(n_808) );
AOI211xp5_ASAP7_75t_L g839 ( .A1(n_734), .A2(n_767), .B(n_840), .C(n_843), .Y(n_839) );
AND2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_735), .B(n_752), .Y(n_751) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_735), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_735), .B(n_800), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_744), .B(n_748), .C(n_749), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI311xp33_ASAP7_75t_L g783 ( .A1(n_740), .A2(n_784), .A3(n_787), .B1(n_791), .C1(n_793), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_740), .B(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AOI21xp33_ASAP7_75t_L g836 ( .A1(n_742), .A2(n_764), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g760 ( .A(n_743), .Y(n_760) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_747), .A2(n_748), .B1(n_803), .B2(n_804), .Y(n_802) );
OAI221xp5_ASAP7_75t_L g818 ( .A1(n_747), .A2(n_757), .B1(n_819), .B2(n_822), .C(n_824), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_748), .B(n_867), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_753), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OAI221xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B1(n_761), .B2(n_764), .C(n_766), .Y(n_755) );
INVx1_ASAP7_75t_L g814 ( .A(n_756), .Y(n_814) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g841 ( .A(n_760), .Y(n_841) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_765), .B(n_849), .Y(n_848) );
AND2x2_ASAP7_75t_L g843 ( .A(n_767), .B(n_794), .Y(n_843) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g846 ( .A(n_772), .Y(n_846) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_774), .A2(n_829), .B1(n_830), .B2(n_839), .Y(n_828) );
AOI211xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_778), .B(n_783), .C(n_798), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AOI21xp33_ASAP7_75t_L g798 ( .A1(n_777), .A2(n_797), .B(n_799), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g806 ( .A1(n_777), .A2(n_807), .B1(n_809), .B2(n_811), .C(n_813), .Y(n_806) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_780), .B(n_814), .Y(n_832) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_792), .B(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_792), .B(n_814), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_797), .B(n_817), .Y(n_816) );
OAI221xp5_ASAP7_75t_L g847 ( .A1(n_803), .A2(n_805), .B1(n_848), .B2(n_850), .C(n_852), .Y(n_847) );
INVxp67_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
AOI211xp5_ASAP7_75t_L g857 ( .A1(n_810), .A2(n_858), .B(n_860), .C(n_866), .Y(n_857) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OAI21xp33_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B(n_816), .Y(n_813) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g859 ( .A(n_821), .Y(n_859) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
OAI321xp33_ASAP7_75t_L g844 ( .A1(n_829), .A2(n_837), .A3(n_845), .B1(n_854), .B2(n_855), .C(n_857), .Y(n_844) );
NOR4xp25_ASAP7_75t_SL g830 ( .A(n_831), .B(n_833), .C(n_835), .D(n_836), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_849), .B(n_865), .Y(n_864) );
CKINVDCx14_ASAP7_75t_R g850 ( .A(n_851), .Y(n_850) );
INVxp67_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
CKINVDCx5p33_ASAP7_75t_R g868 ( .A(n_869), .Y(n_868) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
OR2x2_ASAP7_75t_L g873 ( .A(n_874), .B(n_880), .Y(n_873) );
NAND4xp25_ASAP7_75t_L g874 ( .A(n_875), .B(n_877), .C(n_878), .D(n_879), .Y(n_874) );
NAND3xp33_ASAP7_75t_SL g880 ( .A(n_881), .B(n_887), .C(n_892), .Y(n_880) );
INVx2_ASAP7_75t_SL g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVxp33_ASAP7_75t_SL g904 ( .A(n_905), .Y(n_904) );
NAND4xp75_ASAP7_75t_L g905 ( .A(n_906), .B(n_911), .C(n_914), .D(n_918), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_910), .Y(n_908) );
AND2x2_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .Y(n_911) );
AND2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_917), .Y(n_914) );
AND2x2_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .Y(n_918) );
BUFx3_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
BUFx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
endmodule