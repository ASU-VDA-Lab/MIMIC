module real_aes_1668_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_789;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_0), .B(n_502), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_1), .A2(n_504), .B(n_505), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_2), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_3), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_4), .B(n_269), .Y(n_537) );
INVx1_ASAP7_75t_L g155 ( .A(n_5), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_6), .B(n_174), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_7), .B(n_269), .Y(n_564) );
INVx1_ASAP7_75t_L g238 ( .A(n_8), .Y(n_238) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_9), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_10), .Y(n_203) );
NAND2xp33_ASAP7_75t_L g526 ( .A(n_11), .B(n_266), .Y(n_526) );
INVx2_ASAP7_75t_L g144 ( .A(n_12), .Y(n_144) );
AOI221x1_ASAP7_75t_L g570 ( .A1(n_13), .A2(n_25), .B1(n_502), .B2(n_504), .C(n_571), .Y(n_570) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_14), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_15), .B(n_502), .Y(n_522) );
INVx1_ASAP7_75t_L g267 ( .A(n_16), .Y(n_267) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_17), .A2(n_219), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_18), .B(n_178), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_19), .B(n_269), .Y(n_514) );
AO21x1_ASAP7_75t_L g532 ( .A1(n_20), .A2(n_502), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g109 ( .A(n_21), .Y(n_109) );
INVx1_ASAP7_75t_L g264 ( .A(n_22), .Y(n_264) );
INVx1_ASAP7_75t_SL g184 ( .A(n_23), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_24), .B(n_161), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_26), .Y(n_787) );
AOI33xp33_ASAP7_75t_L g224 ( .A1(n_27), .A2(n_53), .A3(n_150), .B1(n_159), .B2(n_225), .B3(n_226), .Y(n_224) );
NAND2x1_ASAP7_75t_L g545 ( .A(n_28), .B(n_269), .Y(n_545) );
NAND2x1_ASAP7_75t_L g563 ( .A(n_29), .B(n_266), .Y(n_563) );
INVx1_ASAP7_75t_L g195 ( .A(n_30), .Y(n_195) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_31), .A2(n_85), .B(n_144), .Y(n_143) );
OR2x2_ASAP7_75t_L g175 ( .A(n_31), .B(n_85), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_32), .B(n_169), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_33), .B(n_266), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_34), .B(n_269), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_35), .B(n_266), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_36), .A2(n_504), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g149 ( .A(n_37), .Y(n_149) );
AND2x2_ASAP7_75t_L g167 ( .A(n_37), .B(n_155), .Y(n_167) );
AND2x2_ASAP7_75t_L g173 ( .A(n_37), .B(n_152), .Y(n_173) );
OR2x6_ASAP7_75t_L g107 ( .A(n_38), .B(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_39), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_40), .B(n_502), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_41), .B(n_169), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_42), .A2(n_142), .B1(n_174), .B2(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_43), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_44), .B(n_161), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_45), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_46), .B(n_266), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_47), .B(n_219), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_48), .B(n_161), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_49), .A2(n_504), .B(n_562), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_50), .Y(n_251) );
OAI222xp33_ASAP7_75t_L g127 ( .A1(n_51), .A2(n_128), .B1(n_785), .B2(n_786), .C1(n_787), .C2(n_788), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_51), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_52), .B(n_266), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_54), .B(n_161), .Y(n_214) );
INVx1_ASAP7_75t_L g154 ( .A(n_55), .Y(n_154) );
INVx1_ASAP7_75t_L g163 ( .A(n_55), .Y(n_163) );
AND2x2_ASAP7_75t_L g215 ( .A(n_56), .B(n_178), .Y(n_215) );
AOI221xp5_ASAP7_75t_L g236 ( .A1(n_57), .A2(n_73), .B1(n_147), .B2(n_169), .C(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_58), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_59), .B(n_269), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_60), .B(n_142), .Y(n_205) );
AOI21xp5_ASAP7_75t_SL g146 ( .A1(n_61), .A2(n_147), .B(n_156), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_62), .A2(n_504), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g261 ( .A(n_63), .Y(n_261) );
AO21x1_ASAP7_75t_L g534 ( .A1(n_64), .A2(n_504), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_65), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g213 ( .A(n_66), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_67), .B(n_502), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_68), .A2(n_147), .B(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g556 ( .A(n_69), .B(n_179), .Y(n_556) );
INVx1_ASAP7_75t_L g152 ( .A(n_70), .Y(n_152) );
INVx1_ASAP7_75t_L g165 ( .A(n_70), .Y(n_165) );
AND2x2_ASAP7_75t_L g566 ( .A(n_71), .B(n_141), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_72), .B(n_169), .Y(n_227) );
AND2x2_ASAP7_75t_L g186 ( .A(n_74), .B(n_141), .Y(n_186) );
INVx1_ASAP7_75t_L g262 ( .A(n_75), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_76), .A2(n_147), .B(n_183), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_77), .A2(n_147), .B(n_218), .C(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g110 ( .A(n_78), .Y(n_110) );
AND2x2_ASAP7_75t_L g499 ( .A(n_79), .B(n_141), .Y(n_499) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_80), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_81), .B(n_502), .Y(n_516) );
OAI22xp5_ASAP7_75t_SL g798 ( .A1(n_82), .A2(n_490), .B1(n_799), .B2(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_82), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_83), .A2(n_147), .B1(n_222), .B2(n_223), .Y(n_221) );
AND2x2_ASAP7_75t_L g533 ( .A(n_84), .B(n_174), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_86), .B(n_266), .Y(n_515) );
AND2x2_ASAP7_75t_L g548 ( .A(n_87), .B(n_141), .Y(n_548) );
INVx1_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_89), .B(n_269), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_90), .A2(n_504), .B(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_91), .B(n_266), .Y(n_572) );
AND2x2_ASAP7_75t_L g228 ( .A(n_92), .B(n_141), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_93), .B(n_269), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_94), .A2(n_193), .B(n_194), .C(n_197), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_95), .Y(n_803) );
INVx1_ASAP7_75t_SL g117 ( .A(n_96), .Y(n_117) );
BUFx2_ASAP7_75t_SL g796 ( .A(n_96), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_97), .A2(n_504), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_98), .B(n_161), .Y(n_160) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_114), .B(n_802), .Y(n_99) );
INVx2_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g804 ( .A(n_101), .Y(n_804) );
INVx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g103 ( .A(n_104), .B(n_111), .Y(n_103) );
INVx1_ASAP7_75t_L g786 ( .A(n_104), .Y(n_786) );
INVx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_106), .B(n_125), .Y(n_124) );
OR2x6_ASAP7_75t_SL g489 ( .A(n_106), .B(n_125), .Y(n_489) );
AND2x6_ASAP7_75t_SL g784 ( .A(n_106), .B(n_107), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_107), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_127), .B(n_792), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_118), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_119), .A2(n_798), .B(n_801), .Y(n_797) );
NOR2xp33_ASAP7_75t_SL g119 ( .A(n_120), .B(n_126), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_123), .Y(n_801) );
BUFx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_487), .B1(n_490), .B2(n_783), .Y(n_129) );
AOI22x1_ASAP7_75t_L g788 ( .A1(n_130), .A2(n_488), .B1(n_789), .B2(n_791), .Y(n_788) );
INVx1_ASAP7_75t_SL g130 ( .A(n_131), .Y(n_130) );
AND3x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_377), .C(n_440), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_341), .Y(n_133) );
NOR3xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_282), .C(n_311), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_136), .B(n_271), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_187), .B1(n_229), .B2(n_241), .Y(n_136) );
NAND2x1_ASAP7_75t_L g426 ( .A(n_137), .B(n_272), .Y(n_426) );
INVx2_ASAP7_75t_SL g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_176), .Y(n_138) );
INVx2_ASAP7_75t_L g243 ( .A(n_139), .Y(n_243) );
INVx4_ASAP7_75t_L g287 ( .A(n_139), .Y(n_287) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_139), .Y(n_307) );
AND2x4_ASAP7_75t_L g318 ( .A(n_139), .B(n_286), .Y(n_318) );
AND2x2_ASAP7_75t_L g324 ( .A(n_139), .B(n_246), .Y(n_324) );
NOR2x1_ASAP7_75t_SL g454 ( .A(n_139), .B(n_257), .Y(n_454) );
OR2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_145), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_141), .A2(n_192), .B1(n_198), .B2(n_199), .Y(n_191) );
INVx3_ASAP7_75t_L g199 ( .A(n_141), .Y(n_199) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_142), .B(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx4f_ASAP7_75t_L g219 ( .A(n_143), .Y(n_219) );
AND2x4_ASAP7_75t_L g174 ( .A(n_144), .B(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_SL g179 ( .A(n_144), .B(n_175), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_168), .B(n_174), .Y(n_145) );
INVxp67_ASAP7_75t_L g204 ( .A(n_147), .Y(n_204) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_153), .Y(n_147) );
NOR2x1p5_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
INVx1_ASAP7_75t_L g226 ( .A(n_150), .Y(n_226) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OR2x6_ASAP7_75t_L g158 ( .A(n_151), .B(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x6_ASAP7_75t_L g266 ( .A(n_152), .B(n_162), .Y(n_266) );
AND2x6_ASAP7_75t_L g504 ( .A(n_153), .B(n_173), .Y(n_504) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
INVx2_ASAP7_75t_L g159 ( .A(n_154), .Y(n_159) );
AND2x4_ASAP7_75t_L g269 ( .A(n_154), .B(n_164), .Y(n_269) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_155), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_160), .C(n_166), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_SL g183 ( .A1(n_158), .A2(n_166), .B(n_184), .C(n_185), .Y(n_183) );
INVxp67_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_158), .A2(n_166), .B(n_213), .C(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_SL g237 ( .A1(n_158), .A2(n_166), .B(n_238), .C(n_239), .Y(n_237) );
INVx2_ASAP7_75t_L g256 ( .A(n_158), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_158), .A2(n_196), .B1(n_261), .B2(n_262), .Y(n_260) );
AND2x2_ASAP7_75t_L g170 ( .A(n_159), .B(n_171), .Y(n_170) );
INVxp33_ASAP7_75t_L g225 ( .A(n_159), .Y(n_225) );
INVx1_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
AND2x4_ASAP7_75t_L g502 ( .A(n_161), .B(n_167), .Y(n_502) );
AND2x4_ASAP7_75t_L g161 ( .A(n_162), .B(n_164), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g222 ( .A(n_166), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_166), .A2(n_254), .B(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_166), .B(n_174), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_166), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_166), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_166), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_166), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_166), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_166), .A2(n_553), .B(n_554), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_166), .A2(n_563), .B(n_564), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_166), .A2(n_572), .B(n_573), .Y(n_571) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_167), .Y(n_197) );
INVx1_ASAP7_75t_L g206 ( .A(n_169), .Y(n_206) );
AND2x4_ASAP7_75t_L g169 ( .A(n_170), .B(n_172), .Y(n_169) );
INVx1_ASAP7_75t_L g249 ( .A(n_170), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_172), .Y(n_250) );
BUFx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_SL g510 ( .A(n_174), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_174), .A2(n_522), .B(n_523), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_174), .B(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g290 ( .A(n_176), .Y(n_290) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_176), .Y(n_304) );
INVx1_ASAP7_75t_L g315 ( .A(n_176), .Y(n_315) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_176), .Y(n_327) );
AND2x2_ASAP7_75t_L g359 ( .A(n_176), .B(n_257), .Y(n_359) );
AND2x2_ASAP7_75t_L g391 ( .A(n_176), .B(n_275), .Y(n_391) );
INVx1_ASAP7_75t_L g398 ( .A(n_176), .Y(n_398) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_180), .B(n_186), .Y(n_176) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_177), .A2(n_560), .B(n_566), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_178), .A2(n_501), .B(n_503), .Y(n_500) );
OA21x2_ASAP7_75t_L g569 ( .A1(n_178), .A2(n_570), .B(n_574), .Y(n_569) );
OA21x2_ASAP7_75t_L g609 ( .A1(n_178), .A2(n_570), .B(n_574), .Y(n_609) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_207), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g340 ( .A(n_189), .B(n_279), .Y(n_340) );
INVx2_ASAP7_75t_L g414 ( .A(n_189), .Y(n_414) );
AND2x2_ASAP7_75t_L g437 ( .A(n_189), .B(n_207), .Y(n_437) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_190), .B(n_232), .Y(n_278) );
INVx2_ASAP7_75t_L g299 ( .A(n_190), .Y(n_299) );
AND2x4_ASAP7_75t_L g321 ( .A(n_190), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g356 ( .A(n_190), .Y(n_356) );
AND2x2_ASAP7_75t_L g433 ( .A(n_190), .B(n_235), .Y(n_433) );
OR2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_200), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_199), .A2(n_209), .B(n_215), .Y(n_208) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_199), .A2(n_209), .B(n_215), .Y(n_232) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_199), .A2(n_542), .B(n_548), .Y(n_541) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_199), .A2(n_550), .B(n_556), .Y(n_549) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_199), .A2(n_542), .B(n_548), .Y(n_577) );
AO21x2_ASAP7_75t_L g595 ( .A1(n_199), .A2(n_550), .B(n_556), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_204), .B1(n_205), .B2(n_206), .Y(n_200) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g404 ( .A(n_207), .Y(n_404) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_216), .Y(n_207) );
NOR2xp67_ASAP7_75t_L g329 ( .A(n_208), .B(n_299), .Y(n_329) );
AND2x2_ASAP7_75t_L g334 ( .A(n_208), .B(n_299), .Y(n_334) );
INVx2_ASAP7_75t_L g347 ( .A(n_208), .Y(n_347) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_208), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
AND2x4_ASAP7_75t_L g320 ( .A(n_216), .B(n_231), .Y(n_320) );
AND2x2_ASAP7_75t_L g335 ( .A(n_216), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g388 ( .A(n_216), .Y(n_388) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_217), .B(n_235), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_217), .B(n_232), .Y(n_392) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_220), .B(n_228), .Y(n_217) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_218), .A2(n_220), .B(n_228), .Y(n_281) );
INVx2_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_219), .A2(n_236), .B(n_240), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_221), .B(n_227), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVxp33_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2x1p5_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
INVx3_ASAP7_75t_L g296 ( .A(n_231), .Y(n_296) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_232), .Y(n_294) );
AND2x2_ASAP7_75t_L g463 ( .A(n_232), .B(n_464), .Y(n_463) );
INVx3_ASAP7_75t_L g351 ( .A(n_233), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_233), .B(n_388), .Y(n_483) );
BUFx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g298 ( .A(n_234), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x4_ASAP7_75t_L g279 ( .A(n_235), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g322 ( .A(n_235), .Y(n_322) );
INVxp67_ASAP7_75t_L g336 ( .A(n_235), .Y(n_336) );
INVx1_ASAP7_75t_L g396 ( .A(n_235), .Y(n_396) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_235), .Y(n_464) );
INVx1_ASAP7_75t_L g448 ( .A(n_241), .Y(n_448) );
NOR2x1_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
NOR2x1_ASAP7_75t_L g368 ( .A(n_242), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g402 ( .A(n_243), .B(n_274), .Y(n_402) );
OR2x2_ASAP7_75t_L g438 ( .A(n_244), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g420 ( .A(n_245), .B(n_398), .Y(n_420) );
AND2x2_ASAP7_75t_L g472 ( .A(n_245), .B(n_307), .Y(n_472) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_257), .Y(n_245) );
AND2x4_ASAP7_75t_L g274 ( .A(n_246), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g286 ( .A(n_246), .Y(n_286) );
INVx2_ASAP7_75t_L g303 ( .A(n_246), .Y(n_303) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_246), .Y(n_481) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_252), .Y(n_246) );
NOR3xp33_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .C(n_251), .Y(n_248) );
INVx3_ASAP7_75t_L g275 ( .A(n_257), .Y(n_275) );
INVx2_ASAP7_75t_L g369 ( .A(n_257), .Y(n_369) );
AND2x4_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_263), .B(n_270), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B1(n_267), .B2(n_268), .Y(n_263) );
INVxp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVxp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_276), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_273), .B(n_349), .Y(n_366) );
NOR2x1_ASAP7_75t_L g408 ( .A(n_273), .B(n_287), .Y(n_408) );
INVx4_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_274), .B(n_349), .Y(n_486) );
AND2x2_ASAP7_75t_L g302 ( .A(n_275), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g316 ( .A(n_275), .Y(n_316) );
AOI22xp5_ASAP7_75t_SL g364 ( .A1(n_276), .A2(n_365), .B1(n_366), .B2(n_367), .Y(n_364) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
NAND2x1p5_ASAP7_75t_L g361 ( .A(n_277), .B(n_335), .Y(n_361) );
INVx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g422 ( .A(n_278), .B(n_310), .Y(n_422) );
AND2x2_ASAP7_75t_L g292 ( .A(n_279), .B(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g328 ( .A(n_279), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g424 ( .A(n_279), .B(n_414), .Y(n_424) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g346 ( .A(n_281), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g372 ( .A(n_281), .Y(n_372) );
AND2x2_ASAP7_75t_L g462 ( .A(n_281), .B(n_299), .Y(n_462) );
OAI221xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_291), .B1(n_295), .B2(n_300), .C(n_305), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
INVx1_ASAP7_75t_L g363 ( .A(n_285), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_285), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_285), .B(n_359), .Y(n_478) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NOR2xp67_ASAP7_75t_SL g331 ( .A(n_287), .B(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_287), .Y(n_344) );
OR2x2_ASAP7_75t_L g428 ( .A(n_287), .B(n_429), .Y(n_428) );
AND2x4_ASAP7_75t_SL g480 ( .A(n_287), .B(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g349 ( .A(n_289), .Y(n_349) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_290), .Y(n_439) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AOI221x1_ASAP7_75t_L g379 ( .A1(n_292), .A2(n_380), .B1(n_382), .B2(n_385), .C(n_389), .Y(n_379) );
AND2x2_ASAP7_75t_L g365 ( .A(n_293), .B(n_321), .Y(n_365) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x2_ASAP7_75t_L g308 ( .A(n_296), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_296), .B(n_298), .Y(n_435) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
AND2x2_ASAP7_75t_SL g306 ( .A(n_302), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_302), .B(n_315), .Y(n_332) );
INVx2_ASAP7_75t_L g339 ( .A(n_302), .Y(n_339) );
INVx1_ASAP7_75t_L g384 ( .A(n_303), .Y(n_384) );
BUFx2_ASAP7_75t_L g473 ( .A(n_304), .Y(n_473) );
NAND2xp33_ASAP7_75t_SL g305 ( .A(n_306), .B(n_308), .Y(n_305) );
OR2x6_ASAP7_75t_L g338 ( .A(n_307), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g419 ( .A(n_307), .B(n_359), .Y(n_419) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_330), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_319), .B1(n_323), .B2(n_328), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_317), .Y(n_313) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_314), .B(n_318), .Y(n_376) );
AND2x4_ASAP7_75t_L g382 ( .A(n_314), .B(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_SL g314 ( .A(n_315), .B(n_316), .Y(n_314) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_315), .Y(n_407) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_318), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_318), .B(n_349), .Y(n_381) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_318), .Y(n_465) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g412 ( .A(n_320), .B(n_413), .Y(n_412) );
INVx3_ASAP7_75t_L g373 ( .A(n_321), .Y(n_373) );
NAND2x1_ASAP7_75t_SL g417 ( .A(n_321), .B(n_372), .Y(n_417) );
AND2x2_ASAP7_75t_L g451 ( .A(n_321), .B(n_346), .Y(n_451) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B1(n_337), .B2(n_340), .Y(n_330) );
BUFx2_ASAP7_75t_L g446 ( .A(n_332), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_333), .A2(n_402), .B1(n_476), .B2(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2x1p5_ASAP7_75t_L g387 ( .A(n_334), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g354 ( .A(n_335), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_339), .B(n_471), .C(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
AOI211x1_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_350), .B(n_352), .C(n_370), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_345), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
AND2x2_ASAP7_75t_L g432 ( .A(n_346), .B(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_346), .B(n_413), .Y(n_444) );
AND2x2_ASAP7_75t_L g476 ( .A(n_346), .B(n_414), .Y(n_476) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g457 ( .A(n_349), .Y(n_457) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g386 ( .A(n_351), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_364), .Y(n_352) );
AOI22xp5_ASAP7_75t_SL g353 ( .A1(n_354), .A2(n_357), .B1(n_360), .B2(n_362), .Y(n_353) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g394 ( .A(n_356), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g409 ( .A(n_356), .Y(n_409) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_359), .B(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g415 ( .A(n_368), .B(n_398), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_374), .B(n_375), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_372), .B(n_394), .Y(n_469) );
OR2x2_ASAP7_75t_L g447 ( .A(n_373), .B(n_392), .Y(n_447) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND3x1_ASAP7_75t_L g378 ( .A(n_379), .B(n_399), .C(n_423), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_382), .A2(n_412), .B1(n_415), .B2(n_416), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_383), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_SL g456 ( .A(n_383), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_383), .B(n_457), .Y(n_460) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI222xp33_ASAP7_75t_L g443 ( .A1(n_387), .A2(n_444), .B1(n_445), .B2(n_446), .C1(n_447), .C2(n_448), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B1(n_393), .B2(n_397), .Y(n_389) );
INVx1_ASAP7_75t_SL g429 ( .A(n_391), .Y(n_429) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g466 ( .A(n_395), .B(n_462), .Y(n_466) );
NOR2x1_ASAP7_75t_L g399 ( .A(n_400), .B(n_410), .Y(n_399) );
AOI21xp5_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_403), .B(n_409), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_418), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_417), .B(n_431), .Y(n_430) );
OAI21xp5_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_420), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g445 ( .A(n_420), .Y(n_445) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_427), .B2(n_430), .C(n_434), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B(n_438), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
NAND3x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_467), .C(n_474), .Y(n_441) );
NOR2x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_449), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_458), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_451), .B(n_452), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_453), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_461), .B1(n_465), .B2(n_466), .Y(n_458) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_468), .B(n_470), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
AOI22xp5_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_477), .B1(n_479), .B2(n_482), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVxp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
CKINVDCx11_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g800 ( .A(n_490), .Y(n_800) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g791 ( .A(n_491), .Y(n_791) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_692), .Y(n_491) );
NOR4xp25_ASAP7_75t_L g492 ( .A(n_493), .B(n_610), .C(n_636), .D(n_676), .Y(n_492) );
OAI211xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_527), .B(n_557), .C(n_596), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_508), .Y(n_495) );
AND2x2_ASAP7_75t_L g763 ( .A(n_496), .B(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_497), .B(n_508), .Y(n_630) );
BUFx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g558 ( .A(n_498), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_498), .B(n_583), .Y(n_582) );
INVx5_ASAP7_75t_L g616 ( .A(n_498), .Y(n_616) );
NOR2x1_ASAP7_75t_SL g658 ( .A(n_498), .B(n_509), .Y(n_658) );
AND2x2_ASAP7_75t_L g714 ( .A(n_498), .B(n_520), .Y(n_714) );
OR2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_519), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_509), .B(n_520), .Y(n_586) );
AND2x2_ASAP7_75t_L g647 ( .A(n_509), .B(n_616), .Y(n_647) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_517), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_510), .B(n_518), .Y(n_517) );
AO21x2_ASAP7_75t_L g600 ( .A1(n_510), .A2(n_511), .B(n_517), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_516), .Y(n_511) );
AND2x2_ASAP7_75t_L g659 ( .A(n_519), .B(n_583), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_519), .B(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g703 ( .A(n_519), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g736 ( .A(n_519), .B(n_558), .Y(n_736) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g580 ( .A(n_520), .Y(n_580) );
AND2x2_ASAP7_75t_L g613 ( .A(n_520), .B(n_614), .Y(n_613) );
BUFx3_ASAP7_75t_L g648 ( .A(n_520), .Y(n_648) );
OR2x2_ASAP7_75t_L g724 ( .A(n_520), .B(n_583), .Y(n_724) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_540), .Y(n_528) );
AOI211x1_ASAP7_75t_SL g653 ( .A1(n_529), .A2(n_645), .B(n_654), .C(n_656), .Y(n_653) );
AND2x2_ASAP7_75t_SL g698 ( .A(n_529), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_529), .B(n_696), .Y(n_743) );
BUFx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g593 ( .A(n_530), .Y(n_593) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g568 ( .A(n_531), .Y(n_568) );
OAI21x1_ASAP7_75t_SL g531 ( .A1(n_532), .A2(n_534), .B(n_538), .Y(n_531) );
INVx1_ASAP7_75t_L g539 ( .A(n_533), .Y(n_539) );
AOI322xp5_ASAP7_75t_L g557 ( .A1(n_540), .A2(n_558), .A3(n_567), .B1(n_575), .B2(n_578), .C1(n_584), .C2(n_587), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_540), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_549), .Y(n_540) );
INVx2_ASAP7_75t_L g591 ( .A(n_541), .Y(n_591) );
INVxp67_ASAP7_75t_L g633 ( .A(n_541), .Y(n_633) );
BUFx3_ASAP7_75t_L g697 ( .A(n_541), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .Y(n_542) );
INVx2_ASAP7_75t_L g606 ( .A(n_549), .Y(n_606) );
AND2x2_ASAP7_75t_L g655 ( .A(n_549), .B(n_569), .Y(n_655) );
AND2x2_ASAP7_75t_L g699 ( .A(n_549), .B(n_608), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_551), .B(n_555), .Y(n_550) );
AND2x2_ASAP7_75t_L g584 ( .A(n_558), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_558), .B(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_SL g778 ( .A(n_558), .B(n_613), .Y(n_778) );
INVx4_ASAP7_75t_L g583 ( .A(n_559), .Y(n_583) );
AND2x2_ASAP7_75t_L g615 ( .A(n_559), .B(n_616), .Y(n_615) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_559), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_565), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_567), .B(n_652), .Y(n_677) );
INVx1_ASAP7_75t_SL g716 ( .A(n_567), .Y(n_716) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x4_ASAP7_75t_L g607 ( .A(n_568), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_568), .B(n_606), .Y(n_675) );
AND2x2_ASAP7_75t_L g727 ( .A(n_568), .B(n_577), .Y(n_727) );
OR2x2_ASAP7_75t_L g751 ( .A(n_568), .B(n_569), .Y(n_751) );
AND2x2_ASAP7_75t_L g575 ( .A(n_569), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g625 ( .A(n_569), .B(n_606), .Y(n_625) );
AND2x2_ASAP7_75t_SL g681 ( .A(n_569), .B(n_593), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_575), .B(n_688), .Y(n_705) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
BUFx2_ASAP7_75t_L g640 ( .A(n_577), .Y(n_640) );
AND2x4_ASAP7_75t_SL g680 ( .A(n_577), .B(n_594), .Y(n_680) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
OR2x2_ASAP7_75t_L g628 ( .A(n_579), .B(n_582), .Y(n_628) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g597 ( .A(n_580), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g745 ( .A(n_580), .B(n_658), .Y(n_745) );
AND2x2_ASAP7_75t_L g761 ( .A(n_580), .B(n_615), .Y(n_761) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI311xp33_ASAP7_75t_L g731 ( .A1(n_582), .A2(n_670), .A3(n_732), .B(n_734), .C(n_741), .Y(n_731) );
AND2x4_ASAP7_75t_L g598 ( .A(n_583), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g602 ( .A(n_583), .Y(n_602) );
NAND2x1p5_ASAP7_75t_L g672 ( .A(n_583), .B(n_616), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_583), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g715 ( .A(n_583), .B(n_702), .Y(n_715) );
AND2x2_ASAP7_75t_L g601 ( .A(n_585), .B(n_602), .Y(n_601) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_586), .Y(n_619) );
OR2x2_ASAP7_75t_L g708 ( .A(n_586), .B(n_672), .Y(n_708) );
INVx1_ASAP7_75t_L g764 ( .A(n_586), .Y(n_764) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g673 ( .A(n_590), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g687 ( .A(n_590), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g762 ( .A(n_590), .B(n_635), .Y(n_762) );
BUFx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g605 ( .A(n_591), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g624 ( .A(n_591), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g686 ( .A(n_592), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_592), .A2(n_742), .B1(n_743), .B2(n_744), .Y(n_741) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g635 ( .A(n_593), .B(n_606), .Y(n_635) );
AND2x4_ASAP7_75t_L g688 ( .A(n_593), .B(n_595), .Y(n_688) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI21xp33_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_601), .B(n_603), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_597), .A2(n_683), .B1(n_687), .B2(n_689), .Y(n_682) );
AND2x2_ASAP7_75t_SL g642 ( .A(n_598), .B(n_616), .Y(n_642) );
INVx2_ASAP7_75t_L g704 ( .A(n_598), .Y(n_704) );
AND2x2_ASAP7_75t_L g718 ( .A(n_598), .B(n_714), .Y(n_718) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g614 ( .A(n_600), .Y(n_614) );
INVx1_ASAP7_75t_L g667 ( .A(n_600), .Y(n_667) );
INVx1_ASAP7_75t_L g618 ( .A(n_602), .Y(n_618) );
AND3x2_ASAP7_75t_L g646 ( .A(n_602), .B(n_647), .C(n_648), .Y(n_646) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g710 ( .A(n_605), .Y(n_710) );
AND2x2_ASAP7_75t_L g638 ( .A(n_607), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g709 ( .A(n_607), .B(n_710), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_607), .A2(n_721), .B1(n_725), .B2(n_728), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_607), .B(n_755), .Y(n_759) );
BUFx2_ASAP7_75t_L g650 ( .A(n_608), .Y(n_650) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g621 ( .A(n_609), .Y(n_621) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_609), .Y(n_740) );
OAI221xp5_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_620), .B1(n_622), .B2(n_623), .C(n_626), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_617), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g702 ( .A(n_614), .Y(n_702) );
INVx2_ASAP7_75t_SL g691 ( .A(n_615), .Y(n_691) );
AND2x2_ASAP7_75t_L g773 ( .A(n_615), .B(n_640), .Y(n_773) );
INVx4_ASAP7_75t_L g664 ( .A(n_616), .Y(n_664) );
INVx1_ASAP7_75t_L g622 ( .A(n_617), .Y(n_622) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x4_ASAP7_75t_L g733 ( .A(n_621), .B(n_688), .Y(n_733) );
INVx1_ASAP7_75t_SL g772 ( .A(n_621), .Y(n_772) );
AND2x2_ASAP7_75t_L g777 ( .A(n_621), .B(n_680), .Y(n_777) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g719 ( .A(n_625), .Y(n_719) );
OAI21xp5_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_629), .B(n_631), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g652 ( .A(n_633), .Y(n_652) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g649 ( .A(n_635), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g739 ( .A(n_635), .B(n_740), .Y(n_739) );
OAI211xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_641), .B(n_643), .C(n_660), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g732 ( .A(n_639), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_640), .B(n_655), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_640), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g765 ( .A(n_640), .B(n_688), .Y(n_765) );
OAI221xp5_ASAP7_75t_SL g676 ( .A1(n_641), .A2(n_665), .B1(n_677), .B2(n_678), .C(n_682), .Y(n_676) );
INVx3_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g747 ( .A(n_642), .B(n_648), .Y(n_747) );
OAI32xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_649), .A3(n_651), .B1(n_653), .B2(n_657), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_647), .Y(n_737) );
INVx2_ASAP7_75t_L g670 ( .A(n_648), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_L g779 ( .A1(n_648), .A2(n_700), .B(n_780), .C(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g685 ( .A(n_650), .Y(n_685) );
OR2x2_ASAP7_75t_L g781 ( .A(n_650), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_654), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g742 ( .A(n_657), .Y(n_742) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g723 ( .A(n_658), .Y(n_723) );
OAI21xp33_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_669), .B(n_673), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
OR2x2_ASAP7_75t_L g700 ( .A(n_663), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_664), .B(n_667), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_666), .A2(n_698), .B1(n_767), .B2(n_770), .C(n_774), .Y(n_766) );
INVx2_ASAP7_75t_L g769 ( .A(n_666), .Y(n_769) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
OR2x2_ASAP7_75t_L g690 ( .A(n_670), .B(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g757 ( .A(n_670), .B(n_715), .Y(n_757) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g755 ( .A(n_680), .Y(n_755) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_688), .B(n_718), .Y(n_775) );
INVx2_ASAP7_75t_L g782 ( .A(n_688), .Y(n_782) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g752 ( .A1(n_690), .A2(n_753), .B1(n_756), .B2(n_758), .C(n_760), .Y(n_752) );
AND5x1_ASAP7_75t_L g692 ( .A(n_693), .B(n_731), .C(n_746), .D(n_766), .E(n_776), .Y(n_692) );
NOR2xp33_ASAP7_75t_SL g693 ( .A(n_694), .B(n_711), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_700), .B1(n_703), .B2(n_705), .C(n_706), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_696), .B(n_698), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI221xp5_ASAP7_75t_SL g711 ( .A1(n_712), .A2(n_716), .B1(n_717), .B2(n_719), .C(n_720), .Y(n_711) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_716), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
OR2x2_ASAP7_75t_L g729 ( .A(n_724), .B(n_730), .Y(n_729) );
CKINVDCx16_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_737), .B(n_738), .Y(n_734) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B(n_752), .Y(n_746) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVxp67_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVxp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B1(n_763), .B2(n_765), .Y(n_760) );
O2A1O1Ixp33_ASAP7_75t_L g776 ( .A1(n_762), .A2(n_777), .B(n_778), .C(n_779), .Y(n_776) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g780 ( .A(n_773), .Y(n_780) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
CKINVDCx11_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_784), .Y(n_790) );
INVx3_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_797), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
CKINVDCx11_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
CKINVDCx8_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
endmodule