module fake_jpeg_31919_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_14),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_9),
.B(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_16),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_60),
.Y(n_65)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_63),
.B1(n_4),
.B2(n_5),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_70),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_42),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_45),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_75),
.B1(n_45),
.B2(n_6),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_5),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_78),
.B(n_81),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_54),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_8),
.C(n_9),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_70),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_7),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_88),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_35),
.B1(n_22),
.B2(n_23),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_6),
.B(n_7),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_90),
.B(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_19),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_100),
.B(n_101),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_83),
.C(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_10),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_86),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_13),
.B1(n_18),
.B2(n_24),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_11),
.C(n_12),
.Y(n_108)
);

OAI31xp33_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_29),
.A3(n_30),
.B(n_31),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_113),
.A2(n_114),
.B1(n_108),
.B2(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_118),
.B1(n_113),
.B2(n_94),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_119),
.A2(n_120),
.B1(n_112),
.B2(n_110),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_116),
.A2(n_104),
.B1(n_97),
.B2(n_95),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_120),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_123),
.A2(n_114),
.B(n_109),
.Y(n_124)
);

AOI221xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_32),
.B1(n_33),
.B2(n_103),
.C(n_98),
.Y(n_125)
);


endmodule