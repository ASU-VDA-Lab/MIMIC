module fake_ariane_345_n_1881 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1881);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1881;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g195 ( 
.A(n_59),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_144),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_7),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_151),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_110),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_55),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_8),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_80),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_60),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_69),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_92),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_44),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_93),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_98),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_28),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_36),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_51),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_139),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_116),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_70),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_101),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_105),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_24),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_45),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_26),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_24),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_57),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_178),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_20),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_85),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_39),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_114),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_20),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_19),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_115),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_108),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_26),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_77),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_60),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_81),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_84),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_120),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_155),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_19),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_40),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_157),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_57),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_148),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_5),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_83),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_27),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_37),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_142),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_140),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_67),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_75),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_86),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_103),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_56),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_152),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_177),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_182),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_194),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_47),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_168),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_169),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_162),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_5),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_94),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_125),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_52),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_72),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_62),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_192),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_106),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_43),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_14),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_136),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_16),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_25),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_4),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_12),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_78),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_117),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_159),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_36),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_167),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_122),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_113),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_100),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_102),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_130),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_49),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_173),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_12),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_31),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_50),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_118),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_13),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_150),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_32),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_4),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_18),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_37),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_54),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_56),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_87),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_107),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_47),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_65),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_147),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_50),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_31),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_97),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_18),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_165),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_73),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_35),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_76),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_52),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_66),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_45),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_10),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_7),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_119),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_149),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_79),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_0),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_41),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_181),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_44),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_145),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_134),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_158),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_23),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_166),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_186),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_59),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_175),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_129),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_143),
.Y(n_347)
);

BUFx8_ASAP7_75t_SL g348 ( 
.A(n_3),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_29),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_95),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_22),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_6),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_58),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_63),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_74),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_176),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_124),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_156),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_15),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_1),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_34),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_41),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_43),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_9),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_55),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_123),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_0),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_138),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_132),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_90),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_38),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_172),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_27),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_71),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_88),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_89),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_40),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_126),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_35),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_25),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_49),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_10),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_54),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_14),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_64),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_170),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_48),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_127),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_227),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_348),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_300),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_308),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_331),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_262),
.B(n_1),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_353),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_346),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_218),
.B(n_2),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_356),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_203),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_308),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_308),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_231),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_233),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_308),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_384),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_250),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_258),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_235),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_238),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_292),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_258),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_315),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_242),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_384),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_309),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_309),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_251),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_209),
.B(n_2),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_255),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_318),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_265),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_319),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_209),
.B(n_3),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_221),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_379),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_379),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_274),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_195),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_196),
.B(n_6),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_205),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_364),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_381),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_311),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_311),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_341),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_197),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_279),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_387),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_299),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_337),
.B(n_380),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_245),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_R g448 ( 
.A(n_241),
.B(n_137),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_245),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_269),
.B(n_8),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_216),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_207),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_301),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_197),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_302),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_207),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_202),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_202),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_307),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_261),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_321),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_325),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_207),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_324),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_325),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_358),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_214),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_326),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_329),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_303),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_358),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_214),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_214),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_330),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_376),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_376),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_269),
.B(n_9),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_263),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_237),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_253),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_334),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_257),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_263),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_200),
.B(n_11),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_446),
.B(n_337),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_SL g488 ( 
.A(n_448),
.B(n_303),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_405),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_392),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g491 ( 
.A(n_450),
.B(n_269),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_415),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_392),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_403),
.B(n_263),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_399),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_429),
.B(n_221),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_391),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_407),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_389),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_393),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_400),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_413),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_400),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_398),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_401),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_457),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_402),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_446),
.B(n_337),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_406),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_404),
.B(n_272),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_429),
.B(n_297),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_406),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_396),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_394),
.A2(n_367),
.B1(n_312),
.B2(n_277),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_411),
.B(n_412),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_409),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_410),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_424),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_410),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_416),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_416),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_408),
.B(n_217),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_390),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_418),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_417),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_418),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_433),
.A2(n_388),
.B(n_230),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_447),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_429),
.B(n_297),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_447),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_449),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_449),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_421),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_423),
.B(n_272),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_414),
.B(n_430),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_460),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_460),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_R g542 ( 
.A(n_425),
.B(n_232),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_457),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_462),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_431),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_426),
.A2(n_228),
.B1(n_383),
.B2(n_382),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_442),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_428),
.B(n_451),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_462),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_465),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_445),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_428),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_435),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_436),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_465),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_440),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_453),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_455),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_452),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_459),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_466),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_466),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_456),
.Y(n_563)
);

BUFx4f_ASAP7_75t_L g564 ( 
.A(n_531),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_529),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_494),
.B(n_461),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_504),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_542),
.B(n_464),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_491),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_497),
.B(n_468),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_513),
.B(n_538),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_492),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_552),
.Y(n_573)
);

AND2x2_ASAP7_75t_SL g574 ( 
.A(n_500),
.B(n_478),
.Y(n_574)
);

NOR2x1p5_ASAP7_75t_L g575 ( 
.A(n_537),
.B(n_545),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_552),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_491),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_497),
.B(n_469),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_532),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_547),
.B(n_474),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_550),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_491),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_557),
.B(n_483),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_560),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_487),
.B(n_223),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_487),
.B(n_236),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_491),
.A2(n_397),
.B1(n_395),
.B2(n_422),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_506),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_532),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_535),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_551),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_511),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_504),
.Y(n_593)
);

NOR3xp33_ASAP7_75t_L g594 ( 
.A(n_546),
.B(n_486),
.C(n_244),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_556),
.B(n_519),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_551),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_491),
.Y(n_597)
);

AND2x2_ASAP7_75t_SL g598 ( 
.A(n_500),
.B(n_270),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_550),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_535),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_508),
.B(n_454),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_511),
.B(n_239),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_506),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_543),
.B(n_458),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_515),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_548),
.B(n_470),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_R g607 ( 
.A(n_498),
.B(n_463),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_497),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_501),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_491),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_497),
.B(n_471),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_491),
.A2(n_427),
.B1(n_282),
.B2(n_377),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_550),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_546),
.B(n_481),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_550),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_526),
.B(n_467),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_514),
.B(n_240),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_514),
.B(n_471),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_514),
.B(n_246),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_540),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_558),
.B(n_198),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_515),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_495),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_540),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_539),
.B(n_472),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_550),
.Y(n_626)
);

OAI22xp33_ASAP7_75t_L g627 ( 
.A1(n_518),
.A2(n_229),
.B1(n_328),
.B2(n_383),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_536),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_514),
.B(n_247),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_505),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_533),
.B(n_475),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_499),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_539),
.B(n_488),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_541),
.Y(n_634)
);

CKINVDCx11_ASAP7_75t_R g635 ( 
.A(n_503),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_533),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_518),
.B(n_473),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_536),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_533),
.B(n_475),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_522),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_541),
.Y(n_641)
);

OR2x6_ASAP7_75t_L g642 ( 
.A(n_533),
.B(n_481),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_504),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_536),
.B(n_562),
.Y(n_644)
);

AND2x6_ASAP7_75t_L g645 ( 
.A(n_536),
.B(n_256),
.Y(n_645)
);

AND3x1_ASAP7_75t_L g646 ( 
.A(n_562),
.B(n_285),
.C(n_283),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_520),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_553),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_544),
.B(n_482),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_531),
.A2(n_360),
.B1(n_286),
.B2(n_287),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_562),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_527),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_531),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_549),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_562),
.B(n_476),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_555),
.B(n_268),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_555),
.B(n_276),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_490),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_531),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_524),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_SL g661 ( 
.A(n_534),
.B(n_485),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_534),
.A2(n_226),
.B1(n_359),
.B2(n_228),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_561),
.B(n_484),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_504),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_524),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_561),
.B(n_479),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_490),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_504),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_509),
.B(n_293),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_493),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_493),
.B(n_304),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_525),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_489),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_502),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_502),
.A2(n_362),
.B1(n_305),
.B2(n_310),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_525),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_517),
.B(n_432),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_509),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_509),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_507),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_510),
.B(n_476),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_SL g682 ( 
.A(n_559),
.B(n_272),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_563),
.B(n_434),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_509),
.B(n_306),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_510),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_512),
.B(n_482),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_554),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_496),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_509),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_512),
.B(n_477),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_489),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_496),
.Y(n_692)
);

OR2x6_ASAP7_75t_L g693 ( 
.A(n_516),
.B(n_484),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_489),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_516),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_521),
.B(n_477),
.Y(n_696)
);

INVxp33_ASAP7_75t_L g697 ( 
.A(n_489),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_489),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_521),
.B(n_419),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_523),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_523),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_528),
.Y(n_702)
);

BUFx4f_ASAP7_75t_L g703 ( 
.A(n_528),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_530),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_506),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_542),
.B(n_314),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_606),
.B(n_480),
.Y(n_707)
);

OR2x6_ASAP7_75t_L g708 ( 
.A(n_584),
.B(n_419),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_602),
.B(n_248),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_592),
.B(n_335),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_602),
.B(n_290),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_581),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_584),
.B(n_420),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_644),
.A2(n_249),
.B(n_243),
.Y(n_714)
);

OR2x6_ASAP7_75t_L g715 ( 
.A(n_572),
.B(n_420),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_602),
.B(n_633),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_592),
.B(n_199),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_602),
.B(n_296),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_570),
.B(n_213),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_602),
.B(n_323),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_602),
.B(n_336),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_604),
.B(n_380),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_704),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_702),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_648),
.B(n_219),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_591),
.B(n_380),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_608),
.B(n_355),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_703),
.A2(n_369),
.B(n_342),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_569),
.B(n_199),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_608),
.B(n_201),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_565),
.B(n_437),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_569),
.B(n_201),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_699),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_578),
.B(n_219),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_595),
.B(n_226),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_686),
.B(n_204),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_649),
.Y(n_737)
);

NOR3xp33_ASAP7_75t_L g738 ( 
.A(n_580),
.B(n_344),
.C(n_288),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_686),
.B(n_204),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_686),
.B(n_206),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_616),
.B(n_206),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_658),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_582),
.B(n_208),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_571),
.A2(n_361),
.B(n_371),
.C(n_354),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_649),
.B(n_628),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_612),
.A2(n_352),
.B1(n_349),
.B2(n_363),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_649),
.B(n_208),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_649),
.B(n_211),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_628),
.B(n_211),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_703),
.A2(n_369),
.B(n_338),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_688),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_667),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_628),
.B(n_212),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_638),
.B(n_651),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_670),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_688),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_621),
.A2(n_225),
.B1(n_386),
.B2(n_224),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_566),
.A2(n_372),
.B(n_347),
.C(n_374),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_601),
.B(n_351),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_564),
.A2(n_700),
.B(n_695),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_632),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_692),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_638),
.B(n_212),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_692),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_582),
.B(n_597),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_674),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_597),
.B(n_215),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_597),
.B(n_215),
.Y(n_768)
);

AND2x6_ASAP7_75t_SL g769 ( 
.A(n_614),
.B(n_683),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_680),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_581),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_638),
.B(n_651),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_621),
.A2(n_375),
.B(n_351),
.C(n_359),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_585),
.B(n_365),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_587),
.B(n_365),
.C(n_373),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_695),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_610),
.B(n_220),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_701),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_596),
.B(n_437),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_651),
.B(n_220),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_685),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_610),
.B(n_222),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_596),
.B(n_677),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_663),
.B(n_222),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_701),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_663),
.B(n_224),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_663),
.B(n_225),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_573),
.B(n_284),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_610),
.B(n_284),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_576),
.B(n_291),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_585),
.B(n_291),
.Y(n_791)
);

NOR2x1p5_ASAP7_75t_L g792 ( 
.A(n_630),
.B(n_373),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_588),
.Y(n_793)
);

AND2x6_ASAP7_75t_SL g794 ( 
.A(n_614),
.B(n_438),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_586),
.B(n_340),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_586),
.B(n_340),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_577),
.B(n_343),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_611),
.B(n_343),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_588),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_L g800 ( 
.A(n_625),
.B(n_382),
.C(n_350),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_L g801 ( 
.A(n_580),
.B(n_583),
.C(n_594),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_681),
.A2(n_378),
.B(n_350),
.C(n_357),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_583),
.B(n_378),
.C(n_357),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_SL g804 ( 
.A(n_630),
.B(n_345),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_618),
.B(n_345),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_631),
.B(n_366),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_690),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_603),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_574),
.B(n_366),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_639),
.B(n_368),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_603),
.Y(n_811)
);

BUFx8_ASAP7_75t_L g812 ( 
.A(n_640),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_605),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_574),
.B(n_368),
.Y(n_814)
);

NAND3xp33_ASAP7_75t_L g815 ( 
.A(n_666),
.B(n_370),
.C(n_386),
.Y(n_815)
);

OR2x6_ASAP7_75t_L g816 ( 
.A(n_575),
.B(n_438),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_605),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_579),
.B(n_370),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_589),
.B(n_234),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_590),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_600),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_577),
.B(n_198),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_694),
.A2(n_294),
.B(n_252),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_620),
.B(n_254),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_636),
.B(n_259),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_642),
.B(n_11),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_624),
.B(n_260),
.Y(n_827)
);

NOR2x1p5_ASAP7_75t_L g828 ( 
.A(n_652),
.B(n_439),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_634),
.B(n_264),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_577),
.B(n_198),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_622),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_642),
.B(n_13),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_L g833 ( 
.A(n_577),
.B(n_198),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_641),
.B(n_266),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_622),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_696),
.A2(n_654),
.B(n_700),
.C(n_564),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_636),
.B(n_267),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_700),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_642),
.B(n_15),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_636),
.B(n_271),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_642),
.B(n_16),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_693),
.B(n_617),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_617),
.B(n_17),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_693),
.B(n_273),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_693),
.B(n_275),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_655),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_619),
.B(n_17),
.Y(n_847)
);

AOI221xp5_ASAP7_75t_L g848 ( 
.A1(n_627),
.A2(n_444),
.B1(n_443),
.B2(n_441),
.C(n_439),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_619),
.B(n_278),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_629),
.B(n_21),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_629),
.B(n_21),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_577),
.B(n_198),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_568),
.B(n_22),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_706),
.B(n_317),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_614),
.A2(n_444),
.B1(n_443),
.B2(n_441),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_647),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_568),
.B(n_23),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_660),
.Y(n_858)
);

NAND3xp33_ASAP7_75t_L g859 ( 
.A(n_706),
.B(n_320),
.C(n_339),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_656),
.B(n_313),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_697),
.B(n_28),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_564),
.A2(n_280),
.B(n_281),
.C(n_289),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_660),
.Y(n_863)
);

AOI221xp5_ASAP7_75t_L g864 ( 
.A1(n_662),
.A2(n_295),
.B1(n_298),
.B2(n_316),
.C(n_322),
.Y(n_864)
);

NOR2x1_ASAP7_75t_L g865 ( 
.A(n_731),
.B(n_614),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_846),
.B(n_653),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_735),
.B(n_650),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_836),
.A2(n_653),
.B(n_659),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_742),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_735),
.B(n_637),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_809),
.A2(n_598),
.B1(n_646),
.B2(n_609),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_754),
.A2(n_659),
.B(n_697),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_772),
.A2(n_567),
.B(n_664),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_778),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_741),
.A2(n_656),
.B(n_657),
.C(n_669),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_752),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_785),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_755),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_809),
.A2(n_657),
.B(n_669),
.C(n_684),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_783),
.B(n_722),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_751),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_729),
.A2(n_593),
.B(n_668),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_761),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_826),
.A2(n_598),
.B1(n_675),
.B2(n_652),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_729),
.A2(n_679),
.B(n_668),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_732),
.A2(n_679),
.B(n_593),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_737),
.B(n_623),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_737),
.B(n_623),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_707),
.B(n_645),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_732),
.A2(n_664),
.B(n_678),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_743),
.A2(n_664),
.B(n_678),
.Y(n_891)
);

AOI21x1_ASAP7_75t_L g892 ( 
.A1(n_822),
.A2(n_705),
.B(n_665),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_767),
.A2(n_567),
.B(n_689),
.Y(n_893)
);

OAI21xp33_ASAP7_75t_L g894 ( 
.A1(n_804),
.A2(n_682),
.B(n_687),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_768),
.A2(n_782),
.B(n_777),
.Y(n_895)
);

AO21x1_ASAP7_75t_L g896 ( 
.A1(n_716),
.A2(n_684),
.B(n_665),
.Y(n_896)
);

NOR2xp67_ASAP7_75t_L g897 ( 
.A(n_815),
.B(n_609),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_801),
.B(n_745),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_777),
.A2(n_698),
.B(n_673),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_719),
.B(n_645),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_756),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_782),
.A2(n_613),
.B(n_581),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_766),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_812),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_814),
.A2(n_609),
.B1(n_645),
.B2(n_607),
.Y(n_905)
);

O2A1O1Ixp5_ASAP7_75t_L g906 ( 
.A1(n_789),
.A2(n_705),
.B(n_672),
.C(n_676),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_719),
.B(n_734),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_789),
.A2(n_613),
.B(n_581),
.Y(n_908)
);

NAND3xp33_ASAP7_75t_SL g909 ( 
.A(n_814),
.B(n_661),
.C(n_635),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_712),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_838),
.A2(n_645),
.B(n_671),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_765),
.A2(n_671),
.B(n_643),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_749),
.A2(n_613),
.B(n_599),
.Y(n_913)
);

NAND2x1p5_ASAP7_75t_L g914 ( 
.A(n_724),
.B(n_643),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_753),
.A2(n_613),
.B(n_599),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_712),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_763),
.A2(n_599),
.B(n_615),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_762),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_780),
.A2(n_599),
.B(n_615),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_715),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_715),
.Y(n_921)
);

AO21x1_ASAP7_75t_L g922 ( 
.A1(n_853),
.A2(n_671),
.B(n_615),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_770),
.B(n_671),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_842),
.B(n_626),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_781),
.B(n_820),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_708),
.B(n_671),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_847),
.A2(n_643),
.B(n_691),
.C(n_671),
.Y(n_927)
);

BUFx8_ASAP7_75t_L g928 ( 
.A(n_726),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_779),
.B(n_759),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_819),
.A2(n_333),
.B(n_332),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_826),
.A2(n_327),
.B1(n_30),
.B2(n_32),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_824),
.A2(n_198),
.B(n_210),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_821),
.B(n_855),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_733),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_827),
.A2(n_834),
.B(n_829),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_832),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_844),
.B(n_845),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_730),
.A2(n_198),
.B(n_210),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_847),
.A2(n_210),
.B(n_34),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_708),
.B(n_635),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_850),
.A2(n_210),
.B(n_38),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_855),
.B(n_210),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_708),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_856),
.B(n_210),
.Y(n_944)
);

BUFx8_ASAP7_75t_L g945 ( 
.A(n_725),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_764),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_812),
.Y(n_947)
);

NOR3xp33_ASAP7_75t_L g948 ( 
.A(n_853),
.B(n_33),
.C(n_39),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_713),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_858),
.B(n_42),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_850),
.A2(n_42),
.B(n_46),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_712),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_830),
.A2(n_112),
.B(n_189),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_857),
.A2(n_46),
.B(n_48),
.C(n_53),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_830),
.A2(n_852),
.B(n_798),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_712),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_863),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_852),
.A2(n_131),
.B(n_187),
.Y(n_958)
);

AO32x2_ASAP7_75t_L g959 ( 
.A1(n_744),
.A2(n_53),
.A3(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_851),
.A2(n_61),
.B(n_63),
.Y(n_960)
);

NAND3xp33_ASAP7_75t_L g961 ( 
.A(n_857),
.B(n_68),
.C(n_82),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_805),
.A2(n_91),
.B(n_96),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_713),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_806),
.A2(n_99),
.B(n_104),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_747),
.B(n_109),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_800),
.B(n_111),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_851),
.A2(n_135),
.B(n_141),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_810),
.A2(n_146),
.B(n_153),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_748),
.B(n_154),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_825),
.A2(n_160),
.B(n_164),
.Y(n_970)
);

NOR3xp33_ASAP7_75t_L g971 ( 
.A(n_803),
.B(n_171),
.C(n_174),
.Y(n_971)
);

BUFx4f_ASAP7_75t_L g972 ( 
.A(n_713),
.Y(n_972)
);

BUFx8_ASAP7_75t_SL g973 ( 
.A(n_816),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_734),
.B(n_183),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_774),
.B(n_193),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_816),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_774),
.B(n_710),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_793),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_771),
.Y(n_979)
);

O2A1O1Ixp5_ASAP7_75t_L g980 ( 
.A1(n_728),
.A2(n_750),
.B(n_862),
.C(n_714),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_799),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_710),
.B(n_727),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_837),
.A2(n_840),
.B(n_797),
.Y(n_983)
);

BUFx4f_ASAP7_75t_L g984 ( 
.A(n_816),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_808),
.B(n_811),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_813),
.B(n_831),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_817),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_835),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_723),
.B(n_828),
.Y(n_989)
);

NAND3xp33_ASAP7_75t_L g990 ( 
.A(n_864),
.B(n_841),
.C(n_839),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_773),
.A2(n_861),
.B(n_775),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_818),
.A2(n_790),
.B(n_788),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_717),
.B(n_796),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_791),
.B(n_795),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_746),
.B(n_832),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_784),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_839),
.A2(n_841),
.B1(n_757),
.B2(n_746),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_854),
.B(n_769),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_861),
.A2(n_802),
.B(n_758),
.Y(n_999)
);

BUFx8_ASAP7_75t_L g1000 ( 
.A(n_771),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_709),
.B(n_711),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_771),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_736),
.A2(n_740),
.B(n_739),
.C(n_787),
.Y(n_1003)
);

AND2x2_ASAP7_75t_SL g1004 ( 
.A(n_738),
.B(n_718),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_792),
.B(n_771),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_786),
.B(n_720),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_860),
.A2(n_849),
.B(n_721),
.C(n_823),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_833),
.A2(n_859),
.B(n_848),
.Y(n_1008)
);

AND2x2_ASAP7_75t_SL g1009 ( 
.A(n_794),
.B(n_682),
.Y(n_1009)
);

OAI21xp33_ASAP7_75t_L g1010 ( 
.A1(n_735),
.A2(n_804),
.B(n_741),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_822),
.A2(n_852),
.B(n_830),
.Y(n_1011)
);

BUFx12f_ASAP7_75t_L g1012 ( 
.A(n_812),
.Y(n_1012)
);

AO21x1_ASAP7_75t_L g1013 ( 
.A1(n_716),
.A2(n_760),
.B(n_853),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_735),
.A2(n_847),
.B(n_850),
.C(n_843),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_SL g1015 ( 
.A1(n_836),
.A2(n_745),
.B(n_862),
.C(n_772),
.Y(n_1015)
);

NAND3xp33_ASAP7_75t_L g1016 ( 
.A(n_735),
.B(n_537),
.C(n_529),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_742),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_742),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_776),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_776),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_776),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_742),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_737),
.B(n_708),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_735),
.A2(n_847),
.B(n_850),
.C(n_843),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_737),
.B(n_584),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_742),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_735),
.B(n_391),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_846),
.B(n_807),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_776),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_712),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_L g1031 ( 
.A(n_745),
.B(n_491),
.Y(n_1031)
);

OAI21xp33_ASAP7_75t_L g1032 ( 
.A1(n_735),
.A2(n_804),
.B(n_741),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_761),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_895),
.A2(n_896),
.B(n_922),
.Y(n_1034)
);

NAND2x1_ASAP7_75t_L g1035 ( 
.A(n_916),
.B(n_979),
.Y(n_1035)
);

NOR2xp67_ASAP7_75t_SL g1036 ( 
.A(n_1016),
.B(n_1012),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_868),
.A2(n_915),
.B(n_913),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_883),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_917),
.A2(n_919),
.B(n_906),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_907),
.A2(n_977),
.B1(n_1027),
.B2(n_990),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_1033),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1028),
.B(n_870),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1028),
.B(n_933),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_929),
.B(n_880),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1031),
.A2(n_900),
.B(n_992),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_902),
.A2(n_908),
.B(n_872),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_1023),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_1023),
.B(n_1005),
.Y(n_1048)
);

OAI211xp5_ASAP7_75t_L g1049 ( 
.A1(n_1032),
.A2(n_1010),
.B(n_871),
.C(n_960),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_SL g1050 ( 
.A1(n_884),
.A2(n_931),
.B(n_951),
.Y(n_1050)
);

OA21x2_ASAP7_75t_L g1051 ( 
.A1(n_938),
.A2(n_932),
.B(n_980),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_974),
.A2(n_941),
.B(n_939),
.C(n_994),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_1011),
.A2(n_944),
.B(n_885),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_SL g1054 ( 
.A1(n_927),
.A2(n_975),
.B(n_967),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_944),
.A2(n_886),
.B(n_882),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1015),
.A2(n_982),
.B(n_866),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_933),
.B(n_995),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_972),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_866),
.A2(n_889),
.B(n_898),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_SL g1060 ( 
.A(n_904),
.B(n_972),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_SL g1061 ( 
.A1(n_939),
.A2(n_941),
.B(n_951),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_955),
.A2(n_1003),
.B(n_1007),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_890),
.A2(n_891),
.B(n_899),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_995),
.B(n_867),
.Y(n_1064)
);

INVxp67_ASAP7_75t_SL g1065 ( 
.A(n_1000),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_925),
.B(n_996),
.Y(n_1066)
);

NOR2x1_ASAP7_75t_SL g1067 ( 
.A(n_910),
.B(n_952),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_1000),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_925),
.B(n_997),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_873),
.A2(n_911),
.B(n_999),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_999),
.A2(n_993),
.B(n_997),
.C(n_960),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_947),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_879),
.A2(n_967),
.B(n_875),
.C(n_991),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_1005),
.B(n_926),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_893),
.A2(n_912),
.B(n_911),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_910),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1006),
.B(n_876),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_874),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_952),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_983),
.A2(n_912),
.B(n_937),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_878),
.B(n_903),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_923),
.A2(n_991),
.B(n_1008),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_921),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1017),
.B(n_1018),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_952),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_924),
.A2(n_950),
.B(n_964),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_984),
.B(n_905),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_962),
.A2(n_968),
.B(n_950),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1001),
.A2(n_965),
.B(n_969),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_884),
.B(n_894),
.Y(n_1090)
);

AOI31xp33_ASAP7_75t_L g1091 ( 
.A1(n_931),
.A2(n_936),
.A3(n_865),
.B(n_940),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_930),
.A2(n_1026),
.B(n_1022),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_973),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_985),
.A2(n_986),
.B(n_970),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_934),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_957),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_985),
.A2(n_986),
.B(n_1002),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_877),
.B(n_1029),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_942),
.A2(n_966),
.B(n_914),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_943),
.B(n_963),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_914),
.A2(n_953),
.B(n_958),
.Y(n_1101)
);

INVx3_ASAP7_75t_SL g1102 ( 
.A(n_887),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1019),
.B(n_1021),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1020),
.B(n_1004),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_910),
.A2(n_961),
.B(n_1030),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_910),
.A2(n_1030),
.B(n_956),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_920),
.B(n_949),
.Y(n_1107)
);

INVx5_ASAP7_75t_L g1108 ( 
.A(n_956),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_887),
.Y(n_1109)
);

AO31x2_ASAP7_75t_L g1110 ( 
.A1(n_942),
.A2(n_881),
.A3(n_978),
.B(n_981),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_926),
.B(n_888),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_936),
.A2(n_948),
.B1(n_897),
.B2(n_989),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_954),
.A2(n_971),
.B(n_998),
.C(n_1025),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_956),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_987),
.A2(n_909),
.B(n_901),
.C(n_946),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_918),
.A2(n_988),
.B(n_976),
.Y(n_1116)
);

OAI22x1_ASAP7_75t_L g1117 ( 
.A1(n_888),
.A2(n_1009),
.B1(n_945),
.B2(n_928),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1030),
.A2(n_959),
.B(n_928),
.Y(n_1118)
);

OA22x2_ASAP7_75t_L g1119 ( 
.A1(n_945),
.A2(n_884),
.B1(n_871),
.B2(n_870),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_959),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_959),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1014),
.A2(n_1024),
.B(n_907),
.C(n_1010),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1028),
.B(n_907),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_869),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_869),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1014),
.A2(n_1024),
.B(n_935),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1014),
.A2(n_1024),
.B(n_907),
.C(n_1010),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_868),
.A2(n_892),
.B(n_760),
.Y(n_1128)
);

NAND2xp33_ASAP7_75t_SL g1129 ( 
.A(n_907),
.B(n_977),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1014),
.A2(n_1024),
.B(n_907),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_984),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_929),
.B(n_783),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_896),
.A2(n_1013),
.A3(n_922),
.B(n_836),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_868),
.A2(n_892),
.B(n_760),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1028),
.B(n_907),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_868),
.A2(n_892),
.B(n_760),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1028),
.B(n_907),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_952),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_870),
.B(n_648),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_868),
.A2(n_892),
.B(n_760),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1014),
.A2(n_1024),
.B(n_935),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1014),
.A2(n_1024),
.B(n_935),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_929),
.B(n_783),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_984),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1014),
.A2(n_1024),
.B(n_907),
.Y(n_1145)
);

NAND2x1p5_ASAP7_75t_L g1146 ( 
.A(n_1023),
.B(n_737),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_868),
.A2(n_892),
.B(n_760),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_952),
.Y(n_1148)
);

INVx3_ASAP7_75t_SL g1149 ( 
.A(n_904),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_869),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_952),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1014),
.A2(n_1024),
.B(n_907),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_870),
.B(n_648),
.Y(n_1153)
);

OAI21xp33_ASAP7_75t_L g1154 ( 
.A1(n_907),
.A2(n_735),
.B(n_1027),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1028),
.B(n_907),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1028),
.B(n_907),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1028),
.B(n_907),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_868),
.A2(n_892),
.B(n_760),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_869),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1028),
.B(n_907),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1014),
.A2(n_1024),
.B(n_907),
.C(n_1010),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1027),
.B(n_391),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1028),
.B(n_907),
.Y(n_1163)
);

AOI21xp33_ASAP7_75t_L g1164 ( 
.A1(n_1014),
.A2(n_1024),
.B(n_977),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_883),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_868),
.A2(n_892),
.B(n_760),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1027),
.B(n_596),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_868),
.A2(n_892),
.B(n_760),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_868),
.A2(n_892),
.B(n_760),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1023),
.B(n_1005),
.Y(n_1170)
);

INVx3_ASAP7_75t_SL g1171 ( 
.A(n_1149),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1081),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1093),
.Y(n_1173)
);

BUFx10_ASAP7_75t_L g1174 ( 
.A(n_1162),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1123),
.B(n_1135),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_1038),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1078),
.Y(n_1177)
);

NOR2xp67_ASAP7_75t_L g1178 ( 
.A(n_1131),
.B(n_1144),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1123),
.B(n_1135),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1052),
.A2(n_1054),
.B(n_1071),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1050),
.A2(n_1069),
.B1(n_1154),
.B2(n_1040),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1132),
.B(n_1143),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1108),
.Y(n_1183)
);

BUFx2_ASAP7_75t_R g1184 ( 
.A(n_1072),
.Y(n_1184)
);

INVx5_ASAP7_75t_L g1185 ( 
.A(n_1047),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1042),
.B(n_1137),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1137),
.B(n_1155),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1044),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1130),
.A2(n_1152),
.B(n_1145),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1041),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1042),
.B(n_1155),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1090),
.A2(n_1069),
.B(n_1129),
.C(n_1049),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1165),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1108),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1156),
.B(n_1157),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1117),
.Y(n_1196)
);

AO21x2_ASAP7_75t_L g1197 ( 
.A1(n_1061),
.A2(n_1088),
.B(n_1034),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1058),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1156),
.B(n_1157),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1160),
.B(n_1163),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1119),
.A2(n_1139),
.B1(n_1153),
.B2(n_1109),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1160),
.B(n_1163),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1083),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1066),
.B(n_1077),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1043),
.B(n_1064),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1108),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_1079),
.Y(n_1207)
);

INVx5_ASAP7_75t_L g1208 ( 
.A(n_1108),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1122),
.A2(n_1161),
.B(n_1127),
.C(n_1164),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1074),
.B(n_1048),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1074),
.B(n_1048),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1084),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1146),
.Y(n_1213)
);

INVx8_ASAP7_75t_L g1214 ( 
.A(n_1111),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1164),
.A2(n_1073),
.B(n_1113),
.C(n_1126),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1076),
.Y(n_1216)
);

OR2x6_ASAP7_75t_L g1217 ( 
.A(n_1111),
.B(n_1170),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1091),
.A2(n_1043),
.B1(n_1066),
.B2(n_1119),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1065),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1126),
.A2(n_1141),
.B(n_1142),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1142),
.A2(n_1056),
.B(n_1088),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1167),
.B(n_1112),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1096),
.Y(n_1223)
);

NOR2xp67_ASAP7_75t_L g1224 ( 
.A(n_1068),
.B(n_1114),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1084),
.A2(n_1077),
.B(n_1070),
.C(n_1104),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1102),
.Y(n_1226)
);

INVx4_ASAP7_75t_L g1227 ( 
.A(n_1068),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1100),
.B(n_1060),
.Y(n_1228)
);

INVx3_ASAP7_75t_SL g1229 ( 
.A(n_1079),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1095),
.B(n_1107),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1124),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1076),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1089),
.A2(n_1099),
.B(n_1092),
.C(n_1118),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1064),
.B(n_1057),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1104),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1079),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_1125),
.Y(n_1237)
);

O2A1O1Ixp5_ASAP7_75t_L g1238 ( 
.A1(n_1062),
.A2(n_1045),
.B(n_1070),
.C(n_1082),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1120),
.A2(n_1150),
.B1(n_1159),
.B2(n_1121),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1059),
.B(n_1087),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1146),
.B(n_1116),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1138),
.Y(n_1242)
);

BUFx12f_ASAP7_75t_L g1243 ( 
.A(n_1138),
.Y(n_1243)
);

INVx5_ASAP7_75t_L g1244 ( 
.A(n_1148),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1098),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1098),
.B(n_1103),
.Y(n_1246)
);

BUFx4f_ASAP7_75t_L g1247 ( 
.A(n_1148),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1110),
.Y(n_1248)
);

AND2x2_ASAP7_75t_SL g1249 ( 
.A(n_1148),
.B(n_1151),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1115),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1151),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1092),
.A2(n_1036),
.B1(n_1089),
.B2(n_1080),
.Y(n_1252)
);

OR2x6_ASAP7_75t_L g1253 ( 
.A(n_1106),
.B(n_1035),
.Y(n_1253)
);

BUFx12f_ASAP7_75t_L g1254 ( 
.A(n_1151),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1085),
.B(n_1067),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1105),
.A2(n_1051),
.B(n_1086),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_SL g1257 ( 
.A(n_1133),
.B(n_1075),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1133),
.A2(n_1101),
.B1(n_1169),
.B2(n_1128),
.Y(n_1258)
);

INVx5_ASAP7_75t_L g1259 ( 
.A(n_1134),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1136),
.A2(n_1168),
.B(n_1140),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1097),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1094),
.B(n_1166),
.Y(n_1262)
);

OR2x6_ASAP7_75t_SL g1263 ( 
.A(n_1037),
.B(n_1053),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1147),
.B(n_1158),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1046),
.A2(n_1063),
.B(n_1039),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1055),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1132),
.B(n_1143),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1123),
.B(n_1135),
.Y(n_1268)
);

CKINVDCx6p67_ASAP7_75t_R g1269 ( 
.A(n_1149),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1081),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1123),
.B(n_1135),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_SL g1272 ( 
.A1(n_1052),
.A2(n_1024),
.B(n_1014),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1132),
.B(n_1143),
.Y(n_1273)
);

NOR2x1_ASAP7_75t_SL g1274 ( 
.A(n_1108),
.B(n_1087),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1123),
.B(n_1135),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1081),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1081),
.Y(n_1277)
);

BUFx4_ASAP7_75t_R g1278 ( 
.A(n_1093),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1162),
.B(n_1027),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1132),
.B(n_1143),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1123),
.B(n_1135),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1041),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1090),
.A2(n_1027),
.B1(n_1162),
.B2(n_1119),
.Y(n_1283)
);

BUFx8_ASAP7_75t_SL g1284 ( 
.A(n_1093),
.Y(n_1284)
);

BUFx4_ASAP7_75t_SL g1285 ( 
.A(n_1093),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1047),
.B(n_1074),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1149),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1123),
.B(n_1135),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1047),
.B(n_1074),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1052),
.A2(n_1024),
.B(n_1014),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1149),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1041),
.Y(n_1292)
);

INVx4_ASAP7_75t_L g1293 ( 
.A(n_1108),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1052),
.A2(n_1054),
.B(n_1071),
.Y(n_1294)
);

BUFx12f_ASAP7_75t_L g1295 ( 
.A(n_1093),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1108),
.Y(n_1296)
);

AO22x1_ASAP7_75t_L g1297 ( 
.A1(n_1162),
.A2(n_1027),
.B1(n_1090),
.B2(n_630),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1041),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1047),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1081),
.Y(n_1300)
);

AND2x6_ASAP7_75t_L g1301 ( 
.A(n_1090),
.B(n_926),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1052),
.A2(n_1054),
.B(n_1071),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1162),
.B(n_1027),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1047),
.B(n_1074),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1050),
.A2(n_1069),
.B1(n_1071),
.B2(n_1052),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1047),
.Y(n_1306)
);

BUFx8_ASAP7_75t_L g1307 ( 
.A(n_1093),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1231),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1208),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1279),
.A2(n_1303),
.B1(n_1283),
.B2(n_1218),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1218),
.A2(n_1201),
.B1(n_1222),
.B2(n_1181),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1237),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1263),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1177),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1253),
.Y(n_1315)
);

AO21x1_ASAP7_75t_SL g1316 ( 
.A1(n_1220),
.A2(n_1240),
.B(n_1252),
.Y(n_1316)
);

CKINVDCx11_ASAP7_75t_R g1317 ( 
.A(n_1291),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1248),
.Y(n_1318)
);

AO21x2_ASAP7_75t_L g1319 ( 
.A1(n_1260),
.A2(n_1256),
.B(n_1262),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1208),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1245),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1301),
.A2(n_1305),
.B1(n_1182),
.B2(n_1267),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1221),
.A2(n_1238),
.B(n_1265),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1305),
.B(n_1172),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1273),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1193),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1207),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1212),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1301),
.A2(n_1280),
.B1(n_1235),
.B2(n_1250),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1270),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1203),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1239),
.B(n_1205),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1220),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1204),
.B(n_1297),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1276),
.B(n_1277),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1300),
.Y(n_1336)
);

BUFx8_ASAP7_75t_SL g1337 ( 
.A(n_1284),
.Y(n_1337)
);

OAI21xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1272),
.A2(n_1290),
.B(n_1302),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1230),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1301),
.A2(n_1174),
.B1(n_1196),
.B2(n_1294),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1240),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1244),
.Y(n_1342)
);

NAND2x1p5_ASAP7_75t_L g1343 ( 
.A(n_1185),
.B(n_1244),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1246),
.Y(n_1344)
);

NAND2x1p5_ASAP7_75t_L g1345 ( 
.A(n_1185),
.B(n_1244),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1239),
.B(n_1205),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1184),
.Y(n_1347)
);

BUFx8_ASAP7_75t_L g1348 ( 
.A(n_1295),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1301),
.A2(n_1174),
.B1(n_1180),
.B2(n_1189),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_SL g1350 ( 
.A(n_1286),
.Y(n_1350)
);

CKINVDCx11_ASAP7_75t_R g1351 ( 
.A(n_1171),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1188),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1234),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1278),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1225),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1261),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1198),
.B(n_1190),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1243),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1175),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1175),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1298),
.B(n_1292),
.Y(n_1361)
);

CKINVDCx6p67_ASAP7_75t_R g1362 ( 
.A(n_1269),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1192),
.B(n_1179),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1197),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1179),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1228),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1187),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_1307),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1187),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1195),
.A2(n_1268),
.B1(n_1271),
.B2(n_1275),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1249),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1195),
.A2(n_1275),
.B1(n_1288),
.B2(n_1281),
.Y(n_1372)
);

BUFx4f_ASAP7_75t_SL g1373 ( 
.A(n_1307),
.Y(n_1373)
);

AO21x2_ASAP7_75t_L g1374 ( 
.A1(n_1260),
.A2(n_1264),
.B(n_1258),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1200),
.B(n_1268),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1253),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1259),
.Y(n_1377)
);

AO21x1_ASAP7_75t_L g1378 ( 
.A1(n_1209),
.A2(n_1257),
.B(n_1191),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1259),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1226),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1200),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1197),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1214),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1266),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1176),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1271),
.B(n_1288),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1281),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1217),
.B(n_1241),
.Y(n_1388)
);

BUFx12f_ASAP7_75t_L g1389 ( 
.A(n_1287),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1186),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1215),
.B(n_1199),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1219),
.B(n_1282),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1216),
.A2(n_1232),
.B(n_1296),
.Y(n_1393)
);

INVx5_ASAP7_75t_L g1394 ( 
.A(n_1214),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1244),
.Y(n_1395)
);

NAND2x1p5_ASAP7_75t_L g1396 ( 
.A(n_1185),
.B(n_1213),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1202),
.B(n_1233),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_SL g1398 ( 
.A1(n_1173),
.A2(n_1304),
.B1(n_1289),
.B2(n_1286),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1236),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1254),
.Y(n_1400)
);

INVx4_ASAP7_75t_L g1401 ( 
.A(n_1293),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1251),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1229),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1183),
.A2(n_1206),
.B(n_1296),
.Y(n_1404)
);

AOI222xp33_ASAP7_75t_L g1405 ( 
.A1(n_1178),
.A2(n_1210),
.B1(n_1211),
.B2(n_1304),
.C1(n_1289),
.C2(n_1224),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1293),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1242),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1242),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1242),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1183),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1274),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1255),
.Y(n_1412)
);

OAI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1299),
.A2(n_1306),
.B1(n_1227),
.B2(n_1213),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1213),
.Y(n_1414)
);

AOI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1257),
.A2(n_1210),
.B(n_1211),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1194),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1299),
.A2(n_1306),
.B1(n_1247),
.B2(n_1285),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1279),
.A2(n_1090),
.B1(n_1119),
.B2(n_1303),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1182),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1253),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1223),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1223),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1291),
.Y(n_1423)
);

AO21x1_ASAP7_75t_SL g1424 ( 
.A1(n_1220),
.A2(n_1240),
.B(n_1164),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1223),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1203),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1279),
.A2(n_1303),
.B1(n_1027),
.B2(n_1162),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1279),
.A2(n_1090),
.B1(n_1119),
.B2(n_1303),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1223),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1279),
.A2(n_1090),
.B1(n_1119),
.B2(n_1303),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1279),
.B(n_1303),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1279),
.A2(n_1090),
.B1(n_1119),
.B2(n_1303),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1223),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1253),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1341),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1317),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1333),
.B(n_1332),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1318),
.Y(n_1438)
);

AO21x2_ASAP7_75t_L g1439 ( 
.A1(n_1378),
.A2(n_1382),
.B(n_1355),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1321),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1378),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1375),
.B(n_1386),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1363),
.B(n_1370),
.Y(n_1443)
);

NOR2x1_ASAP7_75t_R g1444 ( 
.A(n_1354),
.B(n_1351),
.Y(n_1444)
);

INVxp33_ASAP7_75t_L g1445 ( 
.A(n_1357),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1333),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1313),
.Y(n_1447)
);

AO21x2_ASAP7_75t_L g1448 ( 
.A1(n_1384),
.A2(n_1334),
.B(n_1319),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1324),
.B(n_1424),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1324),
.B(n_1424),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1316),
.B(n_1363),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1359),
.B(n_1360),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1332),
.B(n_1346),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1331),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1365),
.B(n_1367),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1426),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1323),
.A2(n_1393),
.B(n_1376),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1369),
.B(n_1381),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1335),
.B(n_1391),
.Y(n_1459)
);

AOI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1364),
.A2(n_1323),
.B(n_1313),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1385),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1346),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1427),
.B(n_1431),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1328),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1374),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1352),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1330),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1336),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1397),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1374),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1356),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1317),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1315),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1315),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1323),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_SL g1476 ( 
.A1(n_1338),
.A2(n_1428),
.B1(n_1391),
.B2(n_1398),
.Y(n_1476)
);

CKINVDCx12_ASAP7_75t_R g1477 ( 
.A(n_1373),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1387),
.B(n_1372),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1311),
.A2(n_1377),
.B(n_1379),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1412),
.B(n_1339),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1434),
.B(n_1315),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1376),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1420),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1344),
.B(n_1353),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1312),
.B(n_1322),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1337),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1308),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1390),
.B(n_1418),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1415),
.A2(n_1433),
.B(n_1425),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1325),
.B(n_1419),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1421),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1422),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1429),
.Y(n_1493)
);

INVx8_ASAP7_75t_L g1494 ( 
.A(n_1350),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1399),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1402),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1388),
.B(n_1349),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1329),
.A2(n_1404),
.B(n_1432),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1401),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1430),
.B(n_1310),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1314),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1416),
.B(n_1309),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1416),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1410),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1410),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1366),
.B(n_1410),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1414),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1408),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1409),
.Y(n_1509)
);

BUFx4f_ASAP7_75t_L g1510 ( 
.A(n_1309),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1411),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1407),
.B(n_1392),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1380),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1407),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1407),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1340),
.A2(n_1371),
.B1(n_1405),
.B2(n_1347),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1342),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1459),
.B(n_1361),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1441),
.A2(n_1463),
.B(n_1443),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1449),
.B(n_1326),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1459),
.B(n_1413),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1454),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1450),
.B(n_1354),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1464),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1436),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1464),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1503),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1476),
.A2(n_1417),
.B1(n_1403),
.B2(n_1423),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1467),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1467),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1450),
.B(n_1395),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1442),
.B(n_1403),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1468),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1468),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1440),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1451),
.B(n_1320),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1437),
.B(n_1362),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1440),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1503),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1503),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1462),
.B(n_1406),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1456),
.Y(n_1542)
);

NOR2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1453),
.B(n_1406),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1462),
.B(n_1401),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1506),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1438),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1453),
.B(n_1446),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1469),
.B(n_1446),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1469),
.B(n_1406),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1447),
.Y(n_1550)
);

AOI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1500),
.A2(n_1488),
.B1(n_1478),
.B2(n_1485),
.C(n_1484),
.Y(n_1551)
);

NAND4xp25_ASAP7_75t_L g1552 ( 
.A(n_1461),
.B(n_1327),
.C(n_1358),
.D(n_1400),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1502),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1447),
.B(n_1358),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1485),
.A2(n_1350),
.B1(n_1383),
.B2(n_1394),
.Y(n_1555)
);

BUFx12f_ASAP7_75t_L g1556 ( 
.A(n_1472),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1481),
.B(n_1394),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1457),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1466),
.B(n_1327),
.Y(n_1559)
);

OAI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1501),
.A2(n_1394),
.B1(n_1396),
.B2(n_1400),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1452),
.B(n_1351),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1457),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1477),
.Y(n_1563)
);

OAI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1445),
.A2(n_1345),
.B(n_1343),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1471),
.B(n_1383),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1506),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1435),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1545),
.B(n_1460),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1545),
.B(n_1460),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1552),
.B(n_1444),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1519),
.B(n_1495),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1522),
.B(n_1496),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1542),
.B(n_1513),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1547),
.B(n_1455),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1528),
.A2(n_1516),
.B1(n_1497),
.B2(n_1510),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1547),
.B(n_1458),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_L g1577 ( 
.A(n_1551),
.B(n_1509),
.C(n_1507),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1521),
.A2(n_1498),
.B1(n_1479),
.B2(n_1489),
.Y(n_1578)
);

NAND3xp33_ASAP7_75t_L g1579 ( 
.A(n_1559),
.B(n_1509),
.C(n_1507),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1566),
.B(n_1512),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_SL g1581 ( 
.A1(n_1523),
.A2(n_1490),
.B(n_1499),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1550),
.B(n_1512),
.Y(n_1582)
);

OAI221xp5_ASAP7_75t_SL g1583 ( 
.A1(n_1537),
.A2(n_1511),
.B1(n_1470),
.B2(n_1465),
.C(n_1490),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_L g1584 ( 
.A(n_1559),
.B(n_1511),
.C(n_1508),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1518),
.B(n_1480),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1555),
.A2(n_1498),
.B1(n_1479),
.B2(n_1489),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1566),
.B(n_1517),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1548),
.B(n_1524),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1560),
.A2(n_1498),
.B1(n_1494),
.B2(n_1439),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1546),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1548),
.B(n_1448),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1553),
.B(n_1482),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1524),
.B(n_1448),
.Y(n_1593)
);

AOI221xp5_ASAP7_75t_L g1594 ( 
.A1(n_1567),
.A2(n_1491),
.B1(n_1487),
.B2(n_1492),
.C(n_1493),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1553),
.B(n_1482),
.Y(n_1595)
);

AND4x1_ASAP7_75t_L g1596 ( 
.A(n_1564),
.B(n_1444),
.C(n_1477),
.D(n_1337),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1526),
.B(n_1529),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1553),
.B(n_1482),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1529),
.B(n_1504),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1556),
.B(n_1389),
.Y(n_1600)
);

OAI211xp5_ASAP7_75t_SL g1601 ( 
.A1(n_1561),
.A2(n_1532),
.B(n_1554),
.C(n_1562),
.Y(n_1601)
);

NAND4xp25_ASAP7_75t_L g1602 ( 
.A(n_1554),
.B(n_1505),
.C(n_1504),
.D(n_1475),
.Y(n_1602)
);

OAI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1565),
.A2(n_1498),
.B1(n_1487),
.B2(n_1492),
.C(n_1491),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1530),
.B(n_1505),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1531),
.B(n_1520),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1530),
.B(n_1473),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1533),
.B(n_1473),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1556),
.B(n_1389),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1533),
.B(n_1474),
.Y(n_1609)
);

NOR3xp33_ASAP7_75t_SL g1610 ( 
.A(n_1563),
.B(n_1515),
.C(n_1514),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1534),
.B(n_1515),
.C(n_1514),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1534),
.B(n_1541),
.Y(n_1612)
);

NOR3xp33_ASAP7_75t_L g1613 ( 
.A(n_1558),
.B(n_1465),
.C(n_1470),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1544),
.B(n_1474),
.Y(n_1614)
);

NAND3xp33_ASAP7_75t_L g1615 ( 
.A(n_1549),
.B(n_1470),
.C(n_1483),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1600),
.Y(n_1616)
);

NOR2x1_ASAP7_75t_L g1617 ( 
.A(n_1571),
.B(n_1543),
.Y(n_1617)
);

NOR2xp67_ASAP7_75t_L g1618 ( 
.A(n_1602),
.B(n_1558),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1605),
.B(n_1527),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1572),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1590),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1573),
.Y(n_1622)
);

AND2x4_ASAP7_75t_SL g1623 ( 
.A(n_1610),
.B(n_1557),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1605),
.B(n_1539),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1568),
.B(n_1539),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1593),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1568),
.B(n_1540),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1597),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1569),
.B(n_1536),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1591),
.B(n_1535),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1580),
.B(n_1536),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1615),
.B(n_1557),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1608),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1599),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1604),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1611),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1606),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1584),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1611),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1579),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1607),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1609),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1588),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1574),
.B(n_1535),
.Y(n_1644)
);

NAND4xp25_ASAP7_75t_L g1645 ( 
.A(n_1570),
.B(n_1523),
.C(n_1475),
.D(n_1562),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1603),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1576),
.B(n_1538),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1615),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_R g1649 ( 
.A(n_1596),
.B(n_1486),
.Y(n_1649)
);

NOR2xp67_ASAP7_75t_L g1650 ( 
.A(n_1602),
.B(n_1558),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1596),
.B(n_1525),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1629),
.B(n_1581),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1632),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1636),
.B(n_1612),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1629),
.B(n_1581),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1634),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1634),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1618),
.B(n_1613),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1635),
.Y(n_1659)
);

INVxp67_ASAP7_75t_SL g1660 ( 
.A(n_1638),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1636),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1635),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1637),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1629),
.B(n_1592),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1617),
.B(n_1595),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1638),
.B(n_1579),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1637),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1617),
.B(n_1595),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1641),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1619),
.B(n_1598),
.Y(n_1670)
);

INVxp67_ASAP7_75t_SL g1671 ( 
.A(n_1640),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1636),
.B(n_1594),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_1616),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1639),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1639),
.B(n_1584),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1641),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1642),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1639),
.B(n_1585),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1628),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1628),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1640),
.B(n_1614),
.Y(n_1681)
);

NAND2x1_ASAP7_75t_L g1682 ( 
.A(n_1632),
.B(n_1618),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1643),
.B(n_1582),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1621),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1621),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1646),
.B(n_1587),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1643),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1619),
.B(n_1624),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1646),
.B(n_1583),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1630),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1660),
.B(n_1646),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1679),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1679),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1672),
.B(n_1648),
.Y(n_1694)
);

A2O1A1Ixp33_ASAP7_75t_L g1695 ( 
.A1(n_1689),
.A2(n_1650),
.B(n_1648),
.C(n_1645),
.Y(n_1695)
);

NOR2x1p5_ASAP7_75t_SL g1696 ( 
.A(n_1661),
.B(n_1648),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1672),
.A2(n_1577),
.B1(n_1589),
.B2(n_1575),
.C(n_1650),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1680),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1684),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1652),
.B(n_1632),
.Y(n_1700)
);

NAND2x2_ASAP7_75t_L g1701 ( 
.A(n_1673),
.B(n_1649),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1675),
.B(n_1644),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1682),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1671),
.Y(n_1704)
);

INVxp67_ASAP7_75t_SL g1705 ( 
.A(n_1666),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_L g1706 ( 
.A(n_1661),
.B(n_1577),
.C(n_1645),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1652),
.B(n_1632),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1655),
.B(n_1625),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1655),
.B(n_1625),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1661),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1680),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1674),
.B(n_1630),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1684),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1688),
.B(n_1625),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1688),
.B(n_1625),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1658),
.B(n_1623),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1656),
.Y(n_1717)
);

INVxp67_ASAP7_75t_SL g1718 ( 
.A(n_1675),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1674),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1656),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1674),
.B(n_1626),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1653),
.B(n_1627),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1684),
.Y(n_1723)
);

AOI21xp33_ASAP7_75t_L g1724 ( 
.A1(n_1689),
.A2(n_1626),
.B(n_1601),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1685),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1654),
.B(n_1644),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1673),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1653),
.B(n_1665),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1685),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1665),
.B(n_1631),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1673),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1657),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1685),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1668),
.B(n_1631),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1654),
.B(n_1647),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1687),
.B(n_1647),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1668),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1700),
.B(n_1653),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1694),
.B(n_1678),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1703),
.B(n_1653),
.Y(n_1740)
);

INVx1_ASAP7_75t_SL g1741 ( 
.A(n_1731),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1694),
.B(n_1702),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1722),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1697),
.A2(n_1706),
.B1(n_1691),
.B2(n_1724),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1692),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1731),
.B(n_1651),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1692),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1722),
.Y(n_1748)
);

INVx11_ASAP7_75t_L g1749 ( 
.A(n_1727),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1693),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1693),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1691),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1707),
.B(n_1658),
.Y(n_1753)
);

CKINVDCx16_ASAP7_75t_R g1754 ( 
.A(n_1701),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1698),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1697),
.A2(n_1686),
.B1(n_1658),
.B2(n_1681),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1698),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1711),
.Y(n_1758)
);

BUFx2_ASAP7_75t_L g1759 ( 
.A(n_1704),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1711),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1703),
.Y(n_1761)
);

BUFx12f_ASAP7_75t_L g1762 ( 
.A(n_1704),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1707),
.B(n_1658),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1727),
.B(n_1368),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1706),
.A2(n_1686),
.B1(n_1578),
.B2(n_1586),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1730),
.B(n_1734),
.Y(n_1766)
);

NAND3x1_ASAP7_75t_L g1767 ( 
.A(n_1703),
.B(n_1664),
.C(n_1368),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1717),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1717),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1728),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1720),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1703),
.B(n_1682),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1695),
.A2(n_1623),
.B1(n_1683),
.B2(n_1670),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1754),
.B(n_1705),
.Y(n_1774)
);

O2A1O1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1744),
.A2(n_1705),
.B(n_1718),
.C(n_1724),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1741),
.B(n_1718),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1761),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1742),
.B(n_1752),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1756),
.A2(n_1701),
.B1(n_1716),
.B2(n_1702),
.Y(n_1779)
);

XOR2x2_ASAP7_75t_L g1780 ( 
.A(n_1767),
.B(n_1701),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1737),
.B(n_1730),
.Y(n_1781)
);

AOI322xp5_ASAP7_75t_L g1782 ( 
.A1(n_1765),
.A2(n_1719),
.A3(n_1710),
.B1(n_1696),
.B2(n_1712),
.C1(n_1721),
.C2(n_1734),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_SL g1783 ( 
.A(n_1759),
.B(n_1728),
.C(n_1696),
.Y(n_1783)
);

INVxp67_ASAP7_75t_L g1784 ( 
.A(n_1764),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1742),
.B(n_1726),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1759),
.B(n_1726),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1746),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1770),
.B(n_1735),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1767),
.A2(n_1719),
.B1(n_1710),
.B2(n_1728),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1749),
.B(n_1633),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1747),
.Y(n_1791)
);

AOI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1739),
.A2(n_1712),
.B1(n_1721),
.B2(n_1720),
.C(n_1732),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1739),
.B(n_1735),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1773),
.A2(n_1722),
.B(n_1709),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1747),
.Y(n_1795)
);

OAI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1753),
.A2(n_1723),
.B1(n_1733),
.B2(n_1713),
.C(n_1729),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1761),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1762),
.A2(n_1708),
.B1(n_1709),
.B2(n_1714),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1762),
.A2(n_1713),
.B1(n_1733),
.B2(n_1699),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1766),
.B(n_1687),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1787),
.B(n_1766),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1781),
.B(n_1737),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1785),
.B(n_1776),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1775),
.B(n_1793),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1783),
.A2(n_1753),
.B1(n_1763),
.B2(n_1738),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1791),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1775),
.B(n_1743),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1795),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1788),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1777),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1797),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1780),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1786),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1778),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1784),
.B(n_1743),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1800),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1790),
.B(n_1763),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1774),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1799),
.B(n_1782),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1783),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1789),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1818),
.B(n_1749),
.Y(n_1822)
);

NOR3x1_ASAP7_75t_L g1823 ( 
.A(n_1819),
.B(n_1801),
.C(n_1804),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1802),
.Y(n_1824)
);

NOR3xp33_ASAP7_75t_L g1825 ( 
.A(n_1812),
.B(n_1779),
.C(n_1796),
.Y(n_1825)
);

AOI221x1_ASAP7_75t_L g1826 ( 
.A1(n_1820),
.A2(n_1798),
.B1(n_1761),
.B2(n_1760),
.C(n_1745),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1820),
.A2(n_1792),
.B1(n_1755),
.B2(n_1750),
.C(n_1771),
.Y(n_1827)
);

OAI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1807),
.A2(n_1794),
.B(n_1792),
.C(n_1748),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1805),
.A2(n_1748),
.B1(n_1772),
.B2(n_1738),
.Y(n_1829)
);

AOI222xp33_ASAP7_75t_L g1830 ( 
.A1(n_1821),
.A2(n_1750),
.B1(n_1755),
.B2(n_1768),
.C1(n_1751),
.C2(n_1758),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1817),
.B(n_1772),
.Y(n_1831)
);

AOI211xp5_ASAP7_75t_SL g1832 ( 
.A1(n_1814),
.A2(n_1772),
.B(n_1740),
.C(n_1757),
.Y(n_1832)
);

OAI21xp5_ASAP7_75t_SL g1833 ( 
.A1(n_1813),
.A2(n_1740),
.B(n_1769),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1802),
.B(n_1736),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1824),
.B(n_1817),
.Y(n_1835)
);

NOR2x1_ASAP7_75t_L g1836 ( 
.A(n_1822),
.B(n_1810),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1823),
.B(n_1814),
.Y(n_1837)
);

NOR2x1_ASAP7_75t_L g1838 ( 
.A(n_1833),
.B(n_1810),
.Y(n_1838)
);

NOR3xp33_ASAP7_75t_L g1839 ( 
.A(n_1825),
.B(n_1828),
.C(n_1827),
.Y(n_1839)
);

NOR3xp33_ASAP7_75t_L g1840 ( 
.A(n_1831),
.B(n_1821),
.C(n_1809),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1832),
.B(n_1816),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1826),
.B(n_1811),
.C(n_1815),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1834),
.Y(n_1843)
);

NOR4xp25_ASAP7_75t_L g1844 ( 
.A(n_1829),
.B(n_1808),
.C(n_1806),
.D(n_1811),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1830),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1835),
.B(n_1838),
.Y(n_1846)
);

NAND4xp25_ASAP7_75t_L g1847 ( 
.A(n_1839),
.B(n_1803),
.C(n_1817),
.D(n_1816),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1836),
.Y(n_1848)
);

OAI221xp5_ASAP7_75t_L g1849 ( 
.A1(n_1842),
.A2(n_1803),
.B1(n_1699),
.B2(n_1733),
.C(n_1713),
.Y(n_1849)
);

NAND3xp33_ASAP7_75t_SL g1850 ( 
.A(n_1844),
.B(n_1708),
.C(n_1348),
.Y(n_1850)
);

NAND4xp25_ASAP7_75t_L g1851 ( 
.A(n_1840),
.B(n_1740),
.C(n_1714),
.D(n_1715),
.Y(n_1851)
);

NOR3xp33_ASAP7_75t_SL g1852 ( 
.A(n_1837),
.B(n_1348),
.C(n_1732),
.Y(n_1852)
);

NOR2xp67_ASAP7_75t_SL g1853 ( 
.A(n_1843),
.B(n_1841),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1846),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1849),
.A2(n_1845),
.B1(n_1699),
.B2(n_1729),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1848),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1853),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1851),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1850),
.A2(n_1723),
.B1(n_1725),
.B2(n_1729),
.Y(n_1859)
);

OAI22x1_ASAP7_75t_L g1860 ( 
.A1(n_1847),
.A2(n_1725),
.B1(n_1723),
.B2(n_1715),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_R g1861 ( 
.A(n_1857),
.B(n_1852),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1854),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1860),
.Y(n_1863)
);

NOR2x1_ASAP7_75t_L g1864 ( 
.A(n_1856),
.B(n_1736),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1858),
.Y(n_1865)
);

OAI211xp5_ASAP7_75t_L g1866 ( 
.A1(n_1855),
.A2(n_1620),
.B(n_1725),
.C(n_1622),
.Y(n_1866)
);

INVx3_ASAP7_75t_L g1867 ( 
.A(n_1862),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1864),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1865),
.B(n_1859),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1869),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1870),
.B(n_1869),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1871),
.A2(n_1863),
.B(n_1868),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1871),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1873),
.B(n_1869),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1872),
.B(n_1867),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1875),
.A2(n_1867),
.B1(n_1866),
.B2(n_1859),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1874),
.A2(n_1867),
.B1(n_1861),
.B2(n_1663),
.Y(n_1877)
);

OAI21x1_ASAP7_75t_L g1878 ( 
.A1(n_1877),
.A2(n_1876),
.B(n_1659),
.Y(n_1878)
);

AOI322xp5_ASAP7_75t_L g1879 ( 
.A1(n_1878),
.A2(n_1690),
.A3(n_1663),
.B1(n_1667),
.B2(n_1677),
.C1(n_1657),
.C2(n_1659),
.Y(n_1879)
);

OAI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1879),
.A2(n_1676),
.B1(n_1662),
.B2(n_1667),
.C(n_1669),
.Y(n_1880)
);

AOI211xp5_ASAP7_75t_L g1881 ( 
.A1(n_1880),
.A2(n_1677),
.B(n_1662),
.C(n_1669),
.Y(n_1881)
);


endmodule