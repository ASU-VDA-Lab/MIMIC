module fake_netlist_1_12435_n_727 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_727);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_727;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_420;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_78), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_59), .Y(n_102) );
HB1xp67_ASAP7_75t_SL g103 ( .A(n_82), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_9), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_61), .Y(n_105) );
INVx2_ASAP7_75t_SL g106 ( .A(n_87), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_80), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_4), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_39), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_71), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_55), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_54), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_10), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_41), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_50), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_33), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_56), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_70), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_67), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_81), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_25), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_43), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_47), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_31), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_86), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_89), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_66), .Y(n_128) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_2), .Y(n_129) );
INVxp67_ASAP7_75t_SL g130 ( .A(n_57), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_53), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_72), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_16), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_14), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_13), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_35), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_63), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_97), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_14), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_58), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_91), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_69), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_48), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_104), .B(n_0), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_104), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_124), .B(n_1), .Y(n_146) );
INVx6_ASAP7_75t_L g147 ( .A(n_119), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_114), .Y(n_149) );
INVxp67_ASAP7_75t_L g150 ( .A(n_103), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_133), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_151) );
INVx5_ASAP7_75t_L g152 ( .A(n_123), .Y(n_152) );
XNOR2x2_ASAP7_75t_L g153 ( .A(n_111), .B(n_3), .Y(n_153) );
INVx6_ASAP7_75t_L g154 ( .A(n_119), .Y(n_154) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_136), .A2(n_45), .B(n_99), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_136), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_136), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_106), .B(n_4), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_102), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_102), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_119), .B(n_5), .Y(n_161) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_105), .A2(n_46), .B(n_98), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_105), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_150), .B(n_112), .Y(n_164) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_144), .B(n_112), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_150), .B(n_126), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_152), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_159), .B(n_131), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_159), .B(n_106), .Y(n_169) );
NAND2xp33_ASAP7_75t_L g170 ( .A(n_160), .B(n_101), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_160), .B(n_163), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
OAI21xp33_ASAP7_75t_SL g173 ( .A1(n_163), .A2(n_111), .B(n_129), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_152), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
AND2x6_ASAP7_75t_L g176 ( .A(n_161), .B(n_138), .Y(n_176) );
INVxp67_ASAP7_75t_SL g177 ( .A(n_144), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_161), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_151), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_161), .B(n_114), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_151), .Y(n_185) );
OAI22xp33_ASAP7_75t_L g186 ( .A1(n_158), .A2(n_126), .B1(n_108), .B2(n_134), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_149), .B(n_138), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_161), .B(n_109), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_161), .B(n_139), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_144), .B(n_115), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_145), .B(n_113), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_149), .B(n_138), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_164), .B(n_146), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_165), .B(n_144), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_165), .A2(n_144), .B1(n_146), .B2(n_158), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_165), .B(n_154), .Y(n_196) );
NOR2xp33_ASAP7_75t_SL g197 ( .A(n_178), .B(n_107), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_178), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_166), .B(n_149), .Y(n_199) );
AND2x6_ASAP7_75t_SL g200 ( .A(n_166), .B(n_153), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_176), .A2(n_153), .B1(n_148), .B2(n_145), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_168), .B(n_171), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_188), .B(n_149), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_178), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_178), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_176), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_176), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_183), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_189), .B(n_154), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_189), .B(n_154), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_177), .A2(n_148), .B(n_155), .C(n_157), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_175), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_183), .B(n_157), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_186), .B(n_118), .Y(n_214) );
AOI21x1_ASAP7_75t_L g215 ( .A1(n_190), .A2(n_155), .B(n_162), .Y(n_215) );
NOR2xp67_ASAP7_75t_L g216 ( .A(n_173), .B(n_157), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_175), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_180), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_176), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_179), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_176), .B(n_154), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_173), .A2(n_132), .B1(n_121), .B2(n_139), .Y(n_222) );
OAI221xp5_ASAP7_75t_L g223 ( .A1(n_169), .A2(n_135), .B1(n_110), .B2(n_130), .C(n_137), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_185), .A2(n_147), .B1(n_154), .B2(n_117), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_176), .B(n_154), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_176), .Y(n_226) );
INVx8_ASAP7_75t_L g227 ( .A(n_176), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_183), .B(n_147), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_183), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_170), .B(n_147), .Y(n_230) );
INVx2_ASAP7_75t_SL g231 ( .A(n_179), .Y(n_231) );
OAI22xp33_ASAP7_75t_L g232 ( .A1(n_197), .A2(n_191), .B1(n_184), .B2(n_153), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_195), .B(n_184), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_211), .A2(n_191), .B(n_155), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_194), .A2(n_162), .B(n_172), .Y(n_235) );
NOR2xp67_ASAP7_75t_L g236 ( .A(n_222), .B(n_187), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_195), .A2(n_192), .B1(n_147), .B2(n_141), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_196), .A2(n_162), .B(n_172), .Y(n_238) );
OAI21xp33_ASAP7_75t_L g239 ( .A1(n_197), .A2(n_172), .B(n_140), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_224), .A2(n_128), .B(n_116), .C(n_117), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_216), .A2(n_137), .B(n_116), .C(n_120), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_193), .B(n_142), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_208), .A2(n_141), .B1(n_120), .B2(n_122), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_229), .A2(n_122), .B1(n_127), .B2(n_128), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_222), .B(n_5), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_218), .Y(n_246) );
OAI22x1_ASAP7_75t_L g247 ( .A1(n_200), .A2(n_162), .B1(n_127), .B2(n_143), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_227), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_231), .A2(n_113), .B(n_181), .C(n_174), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_206), .B(n_167), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_199), .B(n_162), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_202), .B(n_6), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_216), .A2(n_182), .B(n_181), .C(n_174), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_231), .B(n_167), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_198), .A2(n_182), .B(n_181), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_220), .A2(n_182), .B(n_174), .C(n_167), .Y(n_256) );
O2A1O1Ixp5_ASAP7_75t_L g257 ( .A1(n_215), .A2(n_214), .B(n_224), .C(n_203), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_223), .B(n_6), .Y(n_258) );
OR2x6_ASAP7_75t_L g259 ( .A(n_227), .B(n_123), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_229), .B(n_7), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_227), .A2(n_201), .B1(n_208), .B2(n_212), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_227), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_206), .B(n_125), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_212), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_208), .A2(n_7), .B(n_8), .C(n_9), .Y(n_265) );
OAI21x1_ASAP7_75t_SL g266 ( .A1(n_233), .A2(n_219), .B(n_207), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_251), .A2(n_230), .B(n_221), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_235), .A2(n_215), .B(n_198), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_234), .A2(n_220), .B(n_212), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_264), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_246), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_252), .A2(n_217), .B(n_208), .C(n_210), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_264), .B(n_200), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_260), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_245), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_238), .A2(n_225), .B(n_209), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_258), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_232), .A2(n_228), .B(n_213), .C(n_198), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_248), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_265), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_254), .A2(n_204), .B(n_205), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_236), .B(n_217), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_240), .A2(n_217), .B(n_213), .C(n_204), .Y(n_283) );
BUFx4f_ASAP7_75t_L g284 ( .A(n_259), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_249), .A2(n_205), .B(n_204), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_241), .Y(n_286) );
A2O1A1Ixp33_ASAP7_75t_L g287 ( .A1(n_257), .A2(n_205), .B(n_226), .C(n_219), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_253), .A2(n_227), .B(n_226), .Y(n_288) );
OA21x2_ASAP7_75t_L g289 ( .A1(n_256), .A2(n_207), .B(n_125), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_277), .B(n_232), .Y(n_290) );
OA21x2_ASAP7_75t_L g291 ( .A1(n_287), .A2(n_243), .B(n_239), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_276), .A2(n_247), .B(n_261), .Y(n_292) );
AO31x2_ASAP7_75t_L g293 ( .A1(n_287), .A2(n_237), .A3(n_255), .B(n_242), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_275), .A2(n_243), .B1(n_244), .B2(n_259), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_279), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_286), .B(n_250), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_280), .B(n_270), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_279), .B(n_248), .Y(n_298) );
OA21x2_ASAP7_75t_L g299 ( .A1(n_268), .A2(n_269), .B(n_272), .Y(n_299) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_272), .A2(n_267), .B(n_285), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_282), .Y(n_301) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_289), .A2(n_263), .B(n_259), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_279), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_289), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_278), .A2(n_262), .B(n_248), .C(n_125), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_283), .B(n_248), .Y(n_306) );
OA21x2_ASAP7_75t_L g307 ( .A1(n_288), .A2(n_125), .B(n_123), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_289), .A2(n_123), .B(n_125), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_283), .B(n_8), .Y(n_309) );
OA21x2_ASAP7_75t_L g310 ( .A1(n_266), .A2(n_125), .B(n_123), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_271), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_304), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_290), .B(n_273), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_290), .B(n_274), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_297), .B(n_281), .Y(n_315) );
AOI22xp5_ASAP7_75t_SL g316 ( .A1(n_311), .A2(n_284), .B1(n_279), .B2(n_123), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_298), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_304), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_301), .B(n_284), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_304), .Y(n_320) );
OAI21x1_ASAP7_75t_L g321 ( .A1(n_308), .A2(n_52), .B(n_100), .Y(n_321) );
OA21x2_ASAP7_75t_L g322 ( .A1(n_308), .A2(n_152), .B(n_51), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_297), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_301), .B(n_10), .Y(n_324) );
INVxp67_ASAP7_75t_L g325 ( .A(n_309), .Y(n_325) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_292), .A2(n_306), .B(n_308), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_295), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_309), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_299), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_293), .B(n_11), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_310), .Y(n_331) );
INVxp67_ASAP7_75t_L g332 ( .A(n_295), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_310), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_292), .B(n_60), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_293), .B(n_11), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_310), .Y(n_336) );
OAI21x1_ASAP7_75t_L g337 ( .A1(n_302), .A2(n_62), .B(n_96), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_295), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_310), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_294), .A2(n_306), .B1(n_291), .B2(n_296), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_317), .Y(n_341) );
INVx4_ASAP7_75t_R g342 ( .A(n_333), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_320), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_312), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_320), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_335), .B(n_299), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_312), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_330), .B(n_293), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_333), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_339), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_329), .B(n_293), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_312), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_323), .B(n_293), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_339), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_331), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_335), .B(n_299), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_335), .B(n_299), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_318), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_318), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_318), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_315), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_315), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_329), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_313), .B(n_293), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_329), .B(n_299), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_331), .Y(n_367) );
NOR2x1_ASAP7_75t_SL g368 ( .A(n_334), .B(n_303), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_336), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_316), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_336), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_317), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_336), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_323), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_340), .B(n_293), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_340), .B(n_300), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_330), .B(n_300), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_328), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_326), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_326), .Y(n_380) );
INVx2_ASAP7_75t_SL g381 ( .A(n_316), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_327), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_328), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_325), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_317), .B(n_303), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_326), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_325), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_319), .A2(n_294), .B1(n_291), .B2(n_296), .Y(n_388) );
BUFx2_ASAP7_75t_SL g389 ( .A(n_370), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_364), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_344), .Y(n_391) );
NAND3xp33_ASAP7_75t_L g392 ( .A(n_370), .B(n_324), .C(n_313), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_374), .B(n_324), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_349), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_374), .B(n_324), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_344), .Y(n_396) );
CKINVDCx16_ASAP7_75t_R g397 ( .A(n_370), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_349), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_384), .B(n_314), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_350), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_384), .B(n_314), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_343), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_368), .B(n_317), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_346), .B(n_326), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_343), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_382), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_346), .B(n_326), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_379), .Y(n_408) );
BUFx3_ASAP7_75t_L g409 ( .A(n_381), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_344), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_346), .B(n_317), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_356), .B(n_334), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_356), .B(n_334), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_387), .B(n_319), .Y(n_414) );
INVxp67_ASAP7_75t_L g415 ( .A(n_381), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_350), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_356), .B(n_334), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_364), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_381), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_382), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_357), .B(n_334), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_357), .B(n_334), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_357), .B(n_327), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_375), .B(n_338), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_364), .Y(n_425) );
AOI211xp5_ASAP7_75t_SL g426 ( .A1(n_355), .A2(n_332), .B(n_319), .C(n_338), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_375), .B(n_332), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_378), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_387), .B(n_300), .Y(n_429) );
AND2x4_ASAP7_75t_SL g430 ( .A(n_385), .B(n_298), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_361), .B(n_300), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_375), .B(n_300), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_378), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_376), .B(n_337), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_345), .B(n_310), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_376), .B(n_337), .Y(n_436) );
NAND2xp67_ASAP7_75t_L g437 ( .A(n_376), .B(n_12), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_351), .B(n_337), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_383), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_368), .B(n_303), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_345), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_361), .B(n_305), .C(n_322), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_365), .B(n_12), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_363), .B(n_291), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_383), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_363), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_354), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_365), .B(n_291), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_354), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_347), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_358), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_388), .A2(n_322), .B1(n_298), .B2(n_291), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_358), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_351), .B(n_307), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_360), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_385), .B(n_13), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_360), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_347), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_351), .B(n_307), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_351), .B(n_307), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_404), .B(n_351), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_441), .B(n_353), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_394), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_402), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_423), .B(n_341), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_394), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_398), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_423), .B(n_341), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_397), .B(n_355), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_398), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_409), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_446), .B(n_353), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_427), .B(n_341), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_400), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_427), .B(n_372), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_446), .B(n_367), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_424), .B(n_397), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_404), .B(n_367), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_390), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_400), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_416), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_443), .A2(n_371), .B1(n_385), .B2(n_362), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_407), .B(n_371), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_399), .B(n_362), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_416), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_428), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_401), .B(n_369), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_424), .B(n_372), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_406), .B(n_369), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_415), .B(n_386), .C(n_379), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_428), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_390), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_433), .B(n_373), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_433), .B(n_373), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_411), .B(n_372), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_402), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_439), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_420), .B(n_347), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_405), .B(n_352), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_439), .B(n_366), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_445), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_445), .B(n_366), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_447), .Y(n_503) );
OAI21xp33_ASAP7_75t_SL g504 ( .A1(n_419), .A2(n_342), .B(n_348), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_447), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_412), .B(n_385), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_393), .B(n_366), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_412), .B(n_359), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_395), .B(n_348), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_449), .B(n_348), .Y(n_510) );
INVx2_ASAP7_75t_SL g511 ( .A(n_409), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_409), .B(n_386), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_405), .B(n_359), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_413), .B(n_359), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_403), .B(n_386), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_417), .B(n_352), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_403), .B(n_380), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_449), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_414), .B(n_377), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_403), .B(n_380), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_389), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_451), .Y(n_522) );
AOI21xp5_ASAP7_75t_SL g523 ( .A1(n_392), .A2(n_342), .B(n_322), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_390), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_403), .B(n_380), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_392), .B(n_377), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_440), .B(n_379), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_407), .B(n_377), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_408), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_451), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_432), .B(n_15), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_453), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_440), .B(n_321), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_437), .B(n_15), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_453), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_418), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_408), .Y(n_537) );
AND2x2_ASAP7_75t_SL g538 ( .A(n_417), .B(n_322), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_389), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_408), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_421), .B(n_16), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_435), .B(n_17), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_421), .B(n_17), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_455), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_435), .B(n_18), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_503), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_528), .B(n_429), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_505), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_471), .B(n_440), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_478), .B(n_432), .Y(n_550) );
NOR2x1_ASAP7_75t_L g551 ( .A(n_523), .B(n_440), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_518), .Y(n_552) );
NAND2xp33_ASAP7_75t_SL g553 ( .A(n_477), .B(n_422), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_461), .B(n_422), .Y(n_554) );
OAI21xp33_ASAP7_75t_L g555 ( .A1(n_504), .A2(n_437), .B(n_456), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_478), .B(n_454), .Y(n_556) );
NAND2xp33_ASAP7_75t_SL g557 ( .A(n_511), .B(n_454), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_483), .B(n_455), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_483), .B(n_507), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_531), .B(n_430), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_463), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_461), .B(n_438), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_499), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_466), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_467), .Y(n_565) );
NOR2xp67_ASAP7_75t_SL g566 ( .A(n_542), .B(n_442), .Y(n_566) );
NOR2xp67_ASAP7_75t_SL g567 ( .A(n_545), .B(n_442), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_534), .B(n_457), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_513), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_470), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_474), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_498), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_480), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_534), .A2(n_434), .B1(n_436), .B2(n_460), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_482), .A2(n_434), .B1(n_436), .B2(n_460), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_469), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_510), .B(n_457), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_465), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_481), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_479), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_485), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_500), .B(n_408), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_521), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_486), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_464), .Y(n_585) );
INVxp67_ASAP7_75t_SL g586 ( .A(n_529), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_506), .B(n_426), .Y(n_587) );
CKINVDCx14_ASAP7_75t_R g588 ( .A(n_468), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_539), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_479), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_491), .Y(n_591) );
NAND2x1p5_ASAP7_75t_L g592 ( .A(n_471), .B(n_459), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_495), .B(n_459), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_502), .B(n_448), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_508), .B(n_430), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_497), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_464), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_489), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_501), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_492), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_514), .B(n_430), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_516), .B(n_418), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_496), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_462), .B(n_431), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_511), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_484), .B(n_425), .Y(n_606) );
NAND4xp25_ASAP7_75t_L g607 ( .A(n_541), .B(n_452), .C(n_444), .D(n_458), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_522), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_488), .B(n_425), .Y(n_609) );
INVxp67_ASAP7_75t_L g610 ( .A(n_496), .Y(n_610) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_529), .Y(n_611) );
INVxp67_ASAP7_75t_SL g612 ( .A(n_537), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_537), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_526), .A2(n_458), .B1(n_425), .B2(n_450), .Y(n_614) );
NOR2xp67_ASAP7_75t_L g615 ( .A(n_471), .B(n_450), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_530), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_487), .B(n_410), .Y(n_617) );
OR2x6_ASAP7_75t_L g618 ( .A(n_523), .B(n_533), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_473), .B(n_396), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_538), .B(n_396), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_583), .Y(n_621) );
OAI222xp33_ASAP7_75t_L g622 ( .A1(n_618), .A2(n_543), .B1(n_527), .B2(n_533), .C1(n_509), .C2(n_475), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_551), .B(n_515), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_557), .A2(n_527), .B(n_490), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_607), .A2(n_472), .B1(n_519), .B2(n_532), .C(n_535), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_568), .A2(n_544), .B1(n_493), .B2(n_494), .C(n_540), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_558), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_604), .B(n_476), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g629 ( .A1(n_555), .A2(n_533), .B(n_538), .C(n_515), .Y(n_629) );
OAI321xp33_ASAP7_75t_L g630 ( .A1(n_618), .A2(n_536), .A3(n_524), .B1(n_492), .B2(n_391), .C(n_410), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_589), .B(n_520), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_604), .B(n_540), .Y(n_632) );
OAI221xp5_ASAP7_75t_L g633 ( .A1(n_618), .A2(n_536), .B1(n_524), .B2(n_391), .C(n_307), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_585), .A2(n_525), .B(n_520), .Y(n_634) );
OAI32xp33_ASAP7_75t_L g635 ( .A1(n_553), .A2(n_520), .A3(n_517), .B1(n_515), .B2(n_525), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_588), .B(n_525), .Y(n_636) );
AOI21xp33_ASAP7_75t_SL g637 ( .A1(n_592), .A2(n_517), .B(n_512), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_562), .B(n_517), .Y(n_638) );
AOI22xp33_ASAP7_75t_SL g639 ( .A1(n_587), .A2(n_512), .B1(n_322), .B2(n_321), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_592), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_576), .B(n_18), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_580), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_546), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_594), .B(n_307), .Y(n_644) );
CKINVDCx16_ASAP7_75t_R g645 ( .A(n_578), .Y(n_645) );
AO21x1_ASAP7_75t_L g646 ( .A1(n_586), .A2(n_321), .B(n_302), .Y(n_646) );
AOI322xp5_ASAP7_75t_L g647 ( .A1(n_550), .A2(n_19), .A3(n_20), .B1(n_21), .B2(n_22), .C1(n_23), .C2(n_298), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_597), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_548), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_552), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_594), .B(n_19), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_590), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_605), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g654 ( .A1(n_549), .A2(n_298), .B(n_22), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_617), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_574), .B(n_21), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g657 ( .A1(n_550), .A2(n_23), .A3(n_152), .B1(n_302), .B2(n_27), .C1(n_28), .C2(n_29), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_620), .A2(n_152), .B(n_26), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_561), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_566), .A2(n_152), .B1(n_30), .B2(n_32), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_564), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_597), .Y(n_662) );
NAND2x1_ASAP7_75t_SL g663 ( .A(n_549), .B(n_24), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_577), .B(n_95), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_565), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_577), .B(n_34), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g667 ( .A1(n_629), .A2(n_575), .B1(n_610), .B2(n_585), .C(n_567), .Y(n_667) );
INVx3_ASAP7_75t_L g668 ( .A(n_623), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_654), .A2(n_598), .B1(n_560), .B2(n_610), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_625), .B(n_603), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g671 ( .A1(n_641), .A2(n_614), .B1(n_603), .B2(n_586), .C1(n_612), .C2(n_573), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_645), .A2(n_614), .B1(n_582), .B2(n_615), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_626), .B(n_559), .Y(n_673) );
OAI322xp33_ASAP7_75t_L g674 ( .A1(n_641), .A2(n_556), .A3(n_606), .B1(n_582), .B2(n_547), .C1(n_612), .C2(n_591), .Y(n_674) );
OAI222xp33_ASAP7_75t_L g675 ( .A1(n_624), .A2(n_601), .B1(n_595), .B2(n_554), .C1(n_611), .C2(n_613), .Y(n_675) );
AOI32xp33_ASAP7_75t_L g676 ( .A1(n_623), .A2(n_593), .A3(n_609), .B1(n_619), .B2(n_572), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_621), .A2(n_563), .B1(n_569), .B2(n_616), .Y(n_677) );
NAND2xp33_ASAP7_75t_SL g678 ( .A(n_636), .B(n_613), .Y(n_678) );
AOI321xp33_ASAP7_75t_L g679 ( .A1(n_635), .A2(n_596), .A3(n_608), .B1(n_571), .B2(n_579), .C(n_599), .Y(n_679) );
AOI211xp5_ASAP7_75t_L g680 ( .A1(n_622), .A2(n_611), .B(n_584), .C(n_581), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_656), .A2(n_570), .B1(n_602), .B2(n_600), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_629), .B(n_36), .C(n_37), .Y(n_682) );
NAND3xp33_ASAP7_75t_SL g683 ( .A(n_637), .B(n_94), .C(n_40), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_627), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_648), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_653), .A2(n_38), .B1(n_42), .B2(n_44), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_632), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_643), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_622), .A2(n_49), .B(n_64), .C(n_65), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_631), .A2(n_68), .B1(n_73), .B2(n_74), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_649), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_631), .A2(n_75), .B1(n_76), .B2(n_77), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_634), .A2(n_79), .B1(n_83), .B2(n_84), .C(n_85), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_650), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_651), .A2(n_88), .B1(n_90), .B2(n_92), .C(n_93), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_655), .B(n_628), .Y(n_696) );
AOI211xp5_ASAP7_75t_SL g697 ( .A1(n_630), .A2(n_633), .B(n_658), .C(n_666), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_659), .A2(n_661), .B1(n_665), .B2(n_662), .C(n_639), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_639), .A2(n_640), .B1(n_642), .B2(n_652), .C(n_664), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g700 ( .A1(n_660), .A2(n_644), .B(n_646), .C(n_642), .Y(n_700) );
NAND4xp25_ASAP7_75t_L g701 ( .A(n_647), .B(n_660), .C(n_657), .D(n_638), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g702 ( .A1(n_652), .A2(n_645), .B1(n_397), .B2(n_637), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_663), .B(n_636), .Y(n_703) );
NAND4xp75_ASAP7_75t_L g704 ( .A(n_698), .B(n_669), .C(n_699), .D(n_672), .Y(n_704) );
AO22x2_ASAP7_75t_L g705 ( .A1(n_670), .A2(n_668), .B1(n_673), .B2(n_691), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_696), .Y(n_706) );
NAND4xp75_ASAP7_75t_L g707 ( .A(n_703), .B(n_695), .C(n_692), .D(n_681), .Y(n_707) );
NOR4xp25_ASAP7_75t_L g708 ( .A(n_700), .B(n_674), .C(n_675), .D(n_667), .Y(n_708) );
NOR2x1_ASAP7_75t_L g709 ( .A(n_682), .B(n_683), .Y(n_709) );
NOR4xp25_ASAP7_75t_L g710 ( .A(n_679), .B(n_701), .C(n_702), .D(n_688), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_704), .B(n_690), .C(n_693), .Y(n_711) );
NOR4xp25_ASAP7_75t_L g712 ( .A(n_710), .B(n_668), .C(n_694), .D(n_676), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_706), .B(n_678), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_709), .B(n_689), .C(n_697), .D(n_680), .Y(n_714) );
NOR2x2_ASAP7_75t_L g715 ( .A(n_712), .B(n_707), .Y(n_715) );
INVxp67_ASAP7_75t_L g716 ( .A(n_713), .Y(n_716) );
AND4x2_ASAP7_75t_L g717 ( .A(n_714), .B(n_705), .C(n_708), .D(n_671), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_715), .Y(n_718) );
INVxp33_ASAP7_75t_L g719 ( .A(n_717), .Y(n_719) );
INVx3_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_719), .Y(n_721) );
OAI21xp5_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_716), .B(n_711), .Y(n_722) );
OAI21xp5_ASAP7_75t_SL g723 ( .A1(n_721), .A2(n_671), .B(n_686), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_723), .B(n_720), .Y(n_724) );
NOR3xp33_ASAP7_75t_L g725 ( .A(n_724), .B(n_720), .C(n_722), .Y(n_725) );
OA22x2_ASAP7_75t_L g726 ( .A1(n_725), .A2(n_720), .B1(n_677), .B2(n_687), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_726), .A2(n_720), .B1(n_685), .B2(n_684), .Y(n_727) );
endmodule