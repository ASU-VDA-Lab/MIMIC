module fake_jpeg_19864_n_344 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_17),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_29),
.C(n_38),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_63),
.Y(n_83)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_29),
.C(n_38),
.Y(n_63)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_36),
.CON(n_67),
.SN(n_67)
);

OR2x4_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_33),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_76),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_79),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_41),
.Y(n_79)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx4f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_46),
.B1(n_48),
.B2(n_44),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_58),
.B1(n_54),
.B2(n_57),
.Y(n_119)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_53),
.A2(n_21),
.B1(n_46),
.B2(n_19),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_92),
.B1(n_53),
.B2(n_58),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_57),
.Y(n_117)
);

NOR2xp67_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_30),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_91),
.B(n_99),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_21),
.B1(n_33),
.B2(n_23),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_93),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_53),
.B1(n_58),
.B2(n_66),
.Y(n_116)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_36),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_97),
.Y(n_129)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_35),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_31),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_63),
.CI(n_30),
.CON(n_105),
.SN(n_105)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_108),
.Y(n_136)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_113),
.Y(n_138)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_123),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_117),
.B(n_100),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_121),
.B1(n_128),
.B2(n_134),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_69),
.B1(n_49),
.B2(n_42),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_29),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_127),
.Y(n_139)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_126),
.Y(n_148)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_69),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_77),
.A2(n_35),
.B1(n_1),
.B2(n_3),
.Y(n_128)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_85),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_90),
.B(n_94),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_152),
.B(n_116),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_32),
.Y(n_184)
);

AOI21x1_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_105),
.B(n_87),
.Y(n_173)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_109),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_147),
.B(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_120),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_135),
.B1(n_126),
.B2(n_106),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_100),
.B(n_93),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_155),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_156),
.Y(n_163)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_104),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_159),
.Y(n_164)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_160),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_161),
.B(n_165),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_107),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_139),
.B(n_130),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_180),
.C(n_27),
.Y(n_211)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_183),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_172),
.B(n_173),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_134),
.B1(n_118),
.B2(n_105),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_144),
.B1(n_159),
.B2(n_151),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_131),
.B(n_119),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_123),
.B1(n_114),
.B2(n_113),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_179),
.B1(n_182),
.B2(n_185),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_133),
.B1(n_108),
.B2(n_77),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_80),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_89),
.B1(n_81),
.B2(n_88),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_181),
.A2(n_151),
.B1(n_155),
.B2(n_157),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_89),
.B1(n_4),
.B2(n_5),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_32),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_147),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_136),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_190),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_136),
.B1(n_158),
.B2(n_143),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_202),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_161),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_175),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_0),
.Y(n_242)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_137),
.Y(n_192)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_140),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_201),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_169),
.A2(n_138),
.B(n_148),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_198),
.A2(n_203),
.B(n_206),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_159),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_200),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_138),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_148),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_22),
.B(n_20),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_168),
.B(n_182),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_162),
.A2(n_145),
.B1(n_150),
.B2(n_141),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_185),
.B1(n_163),
.B2(n_170),
.Y(n_218)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_211),
.B(n_24),
.Y(n_221)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_141),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_214),
.B(n_22),
.Y(n_225)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_26),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_217),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_25),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_218),
.A2(n_231),
.B1(n_205),
.B2(n_204),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_170),
.B1(n_167),
.B2(n_166),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_203),
.B1(n_207),
.B2(n_208),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_215),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_241),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_191),
.B(n_24),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_20),
.C(n_5),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_198),
.C(n_195),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_196),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_240),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_188),
.B(n_0),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_235),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_201),
.C(n_203),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_262),
.C(n_232),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_212),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_256),
.Y(n_270)
);

INVxp33_ASAP7_75t_SL g249 ( 
.A(n_228),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_255),
.B1(n_263),
.B2(n_250),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_233),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_259),
.B1(n_265),
.B2(n_216),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_199),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_237),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_217),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_238),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_194),
.C(n_195),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_219),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_234),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_238),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_268),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_274),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_230),
.B(n_229),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_273),
.B(n_281),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_245),
.B(n_192),
.Y(n_274)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_243),
.C(n_224),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_280),
.C(n_255),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_218),
.B1(n_233),
.B2(n_224),
.Y(n_279)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_229),
.C(n_223),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_219),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_246),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_234),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_253),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_300),
.C(n_283),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_251),
.C(n_202),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_287),
.B(n_296),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_270),
.B(n_248),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_291),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_260),
.Y(n_294)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_294),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_239),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_271),
.B(n_278),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_299),
.B1(n_277),
.B2(n_297),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_258),
.B1(n_239),
.B2(n_223),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_209),
.C(n_210),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_298),
.A2(n_267),
.B(n_276),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_301),
.A2(n_307),
.B(n_10),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_310),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_266),
.C(n_222),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_309),
.C(n_290),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_311),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_202),
.B(n_277),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_202),
.C(n_254),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_192),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g313 ( 
.A(n_292),
.B(n_193),
.CI(n_199),
.CON(n_313),
.SN(n_313)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_10),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_290),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_315),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_286),
.B1(n_293),
.B2(n_295),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_318),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_193),
.C(n_7),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_7),
.C(n_9),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_322),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_313),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_321),
.B(n_302),
.Y(n_324)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_324),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_325),
.B(n_326),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_317),
.B(n_312),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_318),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_316),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_334),
.B(n_335),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_320),
.C(n_310),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_311),
.C(n_12),
.Y(n_336)
);

OAI21x1_ASAP7_75t_L g338 ( 
.A1(n_336),
.A2(n_330),
.B(n_331),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_332),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_337),
.Y(n_340)
);

AOI322xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_333),
.A3(n_329),
.B1(n_14),
.B2(n_15),
.C1(n_11),
.C2(n_17),
.Y(n_341)
);

OAI21x1_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_11),
.B(n_12),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_16),
.B(n_247),
.Y(n_344)
);


endmodule