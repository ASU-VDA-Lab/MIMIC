module fake_aes_7187_n_896 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_896);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_896;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_241;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_235;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g109 ( .A(n_36), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_108), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_8), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_99), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_38), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_47), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_12), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_102), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_98), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_66), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_105), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_26), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_63), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_37), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_46), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_57), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_79), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_24), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_82), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_0), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_20), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_1), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_53), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_30), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_20), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_74), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_11), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_67), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_21), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_106), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_41), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_1), .Y(n_140) );
BUFx2_ASAP7_75t_SL g141 ( .A(n_60), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_71), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_100), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_6), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_51), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_87), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_85), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_10), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_43), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_59), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_88), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_64), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_123), .B(n_0), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_123), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_109), .Y(n_156) );
INVx2_ASAP7_75t_SL g157 ( .A(n_117), .Y(n_157) );
BUFx8_ASAP7_75t_SL g158 ( .A(n_113), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_117), .B(n_2), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_147), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_147), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_147), .Y(n_162) );
BUFx12f_ASAP7_75t_L g163 ( .A(n_110), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_147), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_111), .B(n_2), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_109), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_147), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_147), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_116), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_116), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_111), .B(n_3), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_126), .B(n_3), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_126), .B(n_4), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_115), .B(n_4), .Y(n_174) );
INVx5_ASAP7_75t_L g175 ( .A(n_115), .Y(n_175) );
INVx6_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_122), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_168), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_155), .B(n_120), .Y(n_179) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_159), .B(n_122), .Y(n_180) );
INVxp33_ASAP7_75t_L g181 ( .A(n_174), .Y(n_181) );
OAI22xp33_ASAP7_75t_SL g182 ( .A1(n_171), .A2(n_129), .B1(n_148), .B2(n_144), .Y(n_182) );
AO22x2_ASAP7_75t_L g183 ( .A1(n_174), .A2(n_155), .B1(n_159), .B2(n_154), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_155), .B(n_129), .Y(n_184) );
OAI22xp33_ASAP7_75t_SL g185 ( .A1(n_171), .A2(n_148), .B1(n_144), .B2(n_150), .Y(n_185) );
AO22x2_ASAP7_75t_L g186 ( .A1(n_174), .A2(n_134), .B1(n_145), .B2(n_150), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_169), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g188 ( .A1(n_155), .A2(n_135), .B1(n_128), .B2(n_130), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_155), .A2(n_171), .B1(n_165), .B2(n_173), .Y(n_189) );
CKINVDCx6p67_ASAP7_75t_R g190 ( .A(n_175), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_155), .B(n_132), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_168), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_169), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_165), .A2(n_133), .B1(n_137), .B2(n_140), .Y(n_194) );
INVxp67_ASAP7_75t_SL g195 ( .A(n_156), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_169), .Y(n_196) );
OAI22xp5_ASAP7_75t_SL g197 ( .A1(n_172), .A2(n_153), .B1(n_136), .B2(n_138), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_154), .B(n_141), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_168), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_168), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_174), .A2(n_134), .B1(n_151), .B2(n_145), .Y(n_201) );
AND2x2_ASAP7_75t_SL g202 ( .A(n_159), .B(n_151), .Y(n_202) );
AO22x2_ASAP7_75t_L g203 ( .A1(n_159), .A2(n_125), .B1(n_6), .B2(n_7), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_154), .B(n_112), .Y(n_204) );
AO22x2_ASAP7_75t_L g205 ( .A1(n_159), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_154), .B(n_114), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_175), .B(n_118), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_159), .A2(n_139), .B1(n_149), .B2(n_146), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_175), .B(n_119), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_168), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_175), .B(n_121), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_168), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_175), .B(n_124), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_160), .Y(n_214) );
AO22x2_ASAP7_75t_L g215 ( .A1(n_159), .A2(n_5), .B1(n_9), .B2(n_10), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_167), .Y(n_216) );
OAI22xp33_ASAP7_75t_L g217 ( .A1(n_172), .A2(n_152), .B1(n_143), .B2(n_142), .Y(n_217) );
OAI22xp5_ASAP7_75t_SL g218 ( .A1(n_173), .A2(n_131), .B1(n_127), .B2(n_12), .Y(n_218) );
OAI22xp33_ASAP7_75t_L g219 ( .A1(n_175), .A2(n_9), .B1(n_11), .B2(n_13), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_167), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_169), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_169), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_175), .A2(n_156), .B1(n_170), .B2(n_157), .Y(n_223) );
INVx8_ASAP7_75t_L g224 ( .A(n_175), .Y(n_224) );
AO22x2_ASAP7_75t_L g225 ( .A1(n_156), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_167), .Y(n_226) );
INVxp67_ASAP7_75t_SL g227 ( .A(n_195), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_183), .B(n_175), .Y(n_228) );
XNOR2xp5_ASAP7_75t_L g229 ( .A(n_197), .B(n_158), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_195), .Y(n_230) );
XOR2xp5_ASAP7_75t_L g231 ( .A(n_197), .B(n_158), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_187), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_183), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_179), .B(n_175), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_178), .A2(n_170), .B(n_157), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_183), .Y(n_236) );
AOI21x1_ASAP7_75t_L g237 ( .A1(n_187), .A2(n_170), .B(n_162), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_193), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_193), .Y(n_239) );
INVx8_ASAP7_75t_L g240 ( .A(n_224), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_196), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_179), .B(n_175), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_183), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_183), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_191), .B(n_163), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_223), .Y(n_246) );
INVxp33_ASAP7_75t_L g247 ( .A(n_206), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_223), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_180), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_180), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_196), .Y(n_251) );
INVx4_ASAP7_75t_SL g252 ( .A(n_184), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_180), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_198), .B(n_166), .Y(n_254) );
INVxp67_ASAP7_75t_SL g255 ( .A(n_198), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_202), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_202), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_202), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_186), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_186), .Y(n_260) );
XOR2xp5_ASAP7_75t_L g261 ( .A(n_186), .B(n_14), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_206), .B(n_166), .Y(n_262) );
INVx1_ASAP7_75t_SL g263 ( .A(n_204), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_186), .Y(n_264) );
XOR2xp5_ASAP7_75t_L g265 ( .A(n_186), .B(n_15), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_184), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_206), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_204), .Y(n_268) );
AOI21x1_ASAP7_75t_L g269 ( .A1(n_222), .A2(n_199), .B(n_178), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_205), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_181), .B(n_166), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_205), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_205), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_222), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_205), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_189), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_189), .Y(n_277) );
XNOR2x2_ASAP7_75t_L g278 ( .A(n_203), .B(n_205), .Y(n_278) );
XOR2xp5_ASAP7_75t_L g279 ( .A(n_188), .B(n_16), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_201), .B(n_166), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_215), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_215), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_215), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_215), .Y(n_284) );
XNOR2x2_ASAP7_75t_L g285 ( .A(n_203), .B(n_170), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_208), .B(n_163), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_215), .Y(n_287) );
XOR2xp5_ASAP7_75t_L g288 ( .A(n_188), .B(n_16), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_225), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_218), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_255), .B(n_201), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_258), .B(n_203), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_258), .B(n_203), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_280), .B(n_203), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_254), .B(n_194), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_269), .A2(n_185), .B(n_178), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_280), .B(n_225), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_240), .Y(n_298) );
CKINVDCx14_ASAP7_75t_R g299 ( .A(n_261), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_227), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_254), .B(n_194), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_249), .B(n_225), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_249), .B(n_225), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_262), .B(n_185), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_250), .B(n_225), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_240), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_267), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_262), .B(n_217), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_269), .A2(n_199), .B(n_212), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_250), .B(n_190), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_230), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_260), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_253), .B(n_190), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_253), .B(n_190), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_261), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_265), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_237), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_265), .Y(n_319) );
INVx4_ASAP7_75t_L g320 ( .A(n_240), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_240), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_252), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_252), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_237), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_228), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_276), .B(n_217), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_256), .B(n_207), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_228), .Y(n_328) );
AND2x4_ASAP7_75t_SL g329 ( .A(n_236), .B(n_207), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_260), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_247), .B(n_268), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_256), .B(n_207), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_277), .B(n_182), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_236), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_243), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_257), .B(n_182), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_286), .B(n_218), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_257), .B(n_209), .Y(n_338) );
INVx4_ASAP7_75t_L g339 ( .A(n_252), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_263), .B(n_176), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_232), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_243), .B(n_176), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_252), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_267), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_246), .B(n_209), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_320), .B(n_244), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_291), .B(n_266), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_291), .B(n_271), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_313), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_311), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_341), .B(n_270), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_318), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_313), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_320), .B(n_244), .Y(n_354) );
BUFx12f_ASAP7_75t_L g355 ( .A(n_339), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_291), .B(n_233), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_291), .B(n_259), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_291), .B(n_264), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_318), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_313), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_291), .B(n_271), .Y(n_361) );
NOR2x1_ASAP7_75t_SL g362 ( .A(n_320), .B(n_246), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_291), .B(n_248), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_320), .B(n_248), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_320), .B(n_289), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g366 ( .A(n_320), .B(n_270), .Y(n_366) );
CKINVDCx6p67_ASAP7_75t_R g367 ( .A(n_313), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_320), .B(n_272), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_318), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_311), .B(n_272), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_316), .B(n_279), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_311), .Y(n_372) );
INVx4_ASAP7_75t_L g373 ( .A(n_313), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_326), .B(n_273), .Y(n_374) );
INVx6_ASAP7_75t_L g375 ( .A(n_339), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_341), .B(n_273), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_312), .Y(n_377) );
CKINVDCx8_ASAP7_75t_R g378 ( .A(n_298), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_316), .B(n_279), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_373), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_373), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_350), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_367), .Y(n_383) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_359), .Y(n_384) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_355), .Y(n_385) );
CKINVDCx8_ASAP7_75t_R g386 ( .A(n_360), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_373), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_363), .B(n_333), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_360), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_350), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_363), .B(n_297), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_372), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_372), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_360), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_377), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_367), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_360), .Y(n_398) );
INVx1_ASAP7_75t_SL g399 ( .A(n_359), .Y(n_399) );
BUFx12f_ASAP7_75t_SL g400 ( .A(n_373), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_363), .B(n_333), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_353), .Y(n_402) );
INVx2_ASAP7_75t_SL g403 ( .A(n_360), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_377), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_360), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_378), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_360), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_353), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_359), .Y(n_409) );
OAI21xp5_ASAP7_75t_SL g410 ( .A1(n_402), .A2(n_229), .B(n_231), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_387), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_400), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_400), .A2(n_317), .B1(n_319), .B2(n_299), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_382), .B(n_348), .Y(n_414) );
NAND2x1p5_ASAP7_75t_L g415 ( .A(n_383), .B(n_373), .Y(n_415) );
CKINVDCx11_ASAP7_75t_R g416 ( .A(n_385), .Y(n_416) );
CKINVDCx11_ASAP7_75t_R g417 ( .A(n_385), .Y(n_417) );
BUFx4f_ASAP7_75t_L g418 ( .A(n_385), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_387), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_382), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_387), .Y(n_421) );
NAND2x1p5_ASAP7_75t_L g422 ( .A(n_383), .B(n_360), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_406), .A2(n_319), .B1(n_317), .B2(n_371), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_382), .B(n_348), .Y(n_424) );
OAI21xp5_ASAP7_75t_SL g425 ( .A1(n_402), .A2(n_229), .B(n_231), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_391), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_391), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_406), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_391), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g430 ( .A1(n_383), .A2(n_299), .B1(n_278), .B2(n_362), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_402), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_393), .B(n_337), .Y(n_432) );
BUFx10_ASAP7_75t_L g433 ( .A(n_403), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_393), .B(n_348), .Y(n_434) );
INVx6_ASAP7_75t_L g435 ( .A(n_383), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_408), .A2(n_378), .B1(n_367), .B2(n_347), .Y(n_436) );
INVx8_ASAP7_75t_L g437 ( .A(n_380), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_393), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_400), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_408), .Y(n_441) );
OAI22xp33_ASAP7_75t_L g442 ( .A1(n_397), .A2(n_379), .B1(n_371), .B2(n_378), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_394), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_400), .A2(n_290), .B1(n_379), .B2(n_371), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_397), .A2(n_278), .B1(n_362), .B2(n_285), .Y(n_445) );
BUFx8_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_380), .Y(n_447) );
BUFx2_ASAP7_75t_SL g448 ( .A(n_380), .Y(n_448) );
BUFx4f_ASAP7_75t_L g449 ( .A(n_380), .Y(n_449) );
BUFx8_ASAP7_75t_L g450 ( .A(n_394), .Y(n_450) );
BUFx10_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_380), .A2(n_285), .B1(n_294), .B2(n_307), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_394), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_442), .A2(n_379), .B1(n_297), .B2(n_288), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_411), .B(n_384), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_416), .Y(n_456) );
OAI21xp5_ASAP7_75t_SL g457 ( .A1(n_410), .A2(n_288), .B(n_297), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_450), .A2(n_380), .B1(n_381), .B2(n_388), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_430), .A2(n_297), .B1(n_294), .B2(n_361), .Y(n_459) );
BUFx12f_ASAP7_75t_L g460 ( .A(n_416), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_423), .A2(n_294), .B1(n_361), .B2(n_328), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_440), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_420), .Y(n_463) );
CKINVDCx6p67_ASAP7_75t_R g464 ( .A(n_417), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_452), .A2(n_294), .B1(n_361), .B2(n_328), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_450), .A2(n_328), .B1(n_364), .B2(n_389), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_426), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_450), .A2(n_328), .B1(n_364), .B2(n_389), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g469 ( .A1(n_418), .A2(n_388), .B1(n_381), .B2(n_328), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_448), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_412), .A2(n_388), .B1(n_381), .B2(n_384), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_417), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_427), .Y(n_473) );
BUFx12f_ASAP7_75t_L g474 ( .A(n_446), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_432), .B(n_396), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_445), .A2(n_328), .B1(n_364), .B2(n_401), .Y(n_476) );
OAI22xp33_ASAP7_75t_L g477 ( .A1(n_418), .A2(n_388), .B1(n_381), .B2(n_328), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_418), .A2(n_388), .B1(n_381), .B2(n_344), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_444), .A2(n_364), .B1(n_401), .B2(n_392), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_429), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_436), .A2(n_344), .B1(n_409), .B2(n_399), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_414), .A2(n_364), .B1(n_392), .B2(n_354), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_438), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_431), .Y(n_484) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_425), .A2(n_282), .B(n_275), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_441), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_414), .B(n_396), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_443), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_446), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_424), .A2(n_392), .B1(n_346), .B2(n_354), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_411), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_453), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_446), .A2(n_355), .B1(n_292), .B2(n_293), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_424), .B(n_396), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_419), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_434), .B(n_404), .Y(n_496) );
OAI22xp33_ASAP7_75t_L g497 ( .A1(n_439), .A2(n_355), .B1(n_349), .B2(n_358), .Y(n_497) );
INVx4_ASAP7_75t_L g498 ( .A(n_437), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_428), .B(n_331), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_437), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_439), .A2(n_409), .B1(n_399), .B2(n_358), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_419), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_434), .A2(n_354), .B1(n_346), .B2(n_349), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_421), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_413), .A2(n_354), .B1(n_346), .B2(n_349), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_441), .A2(n_354), .B1(n_346), .B2(n_349), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_449), .A2(n_282), .B(n_275), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_449), .A2(n_409), .B1(n_399), .B2(n_357), .Y(n_508) );
OAI21xp33_ASAP7_75t_L g509 ( .A1(n_415), .A2(n_219), .B(n_157), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_421), .Y(n_510) );
OAI21xp5_ASAP7_75t_SL g511 ( .A1(n_415), .A2(n_219), .B(n_292), .Y(n_511) );
OAI21xp5_ASAP7_75t_SL g512 ( .A1(n_422), .A2(n_293), .B(n_292), .Y(n_512) );
CKINVDCx11_ASAP7_75t_R g513 ( .A(n_433), .Y(n_513) );
INVx4_ASAP7_75t_L g514 ( .A(n_437), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_449), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_437), .A2(n_292), .B1(n_293), .B2(n_404), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_435), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_422), .Y(n_518) );
BUFx3_ASAP7_75t_L g519 ( .A(n_433), .Y(n_519) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_435), .A2(n_331), .B1(n_284), .B2(n_283), .C1(n_287), .C2(n_302), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_435), .B(n_356), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_447), .B(n_387), .Y(n_522) );
INVx3_ASAP7_75t_L g523 ( .A(n_433), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_435), .A2(n_346), .B1(n_368), .B2(n_293), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_487), .B(n_404), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_465), .A2(n_368), .B1(n_302), .B2(n_305), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_457), .A2(n_333), .B1(n_157), .B2(n_304), .C(n_326), .Y(n_527) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_498), .A2(n_447), .B1(n_451), .B2(n_422), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_454), .A2(n_357), .B1(n_287), .B2(n_284), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_466), .A2(n_447), .B1(n_386), .B2(n_283), .Y(n_530) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_512), .A2(n_369), .B(n_352), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_455), .B(n_405), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_499), .B(n_177), .C(n_169), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_459), .A2(n_368), .B1(n_302), .B2(n_305), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_494), .B(n_302), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_455), .Y(n_536) );
OAI21xp5_ASAP7_75t_SL g537 ( .A1(n_458), .A2(n_305), .B(n_303), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_468), .A2(n_386), .B1(n_407), .B2(n_403), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_496), .B(n_303), .Y(n_539) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_498), .A2(n_451), .B1(n_407), .B2(n_403), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_463), .B(n_405), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_463), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_476), .A2(n_368), .B1(n_305), .B2(n_303), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_509), .A2(n_368), .B1(n_365), .B2(n_325), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_467), .B(n_451), .Y(n_545) );
INVxp67_ASAP7_75t_L g546 ( .A(n_519), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_479), .A2(n_365), .B1(n_325), .B2(n_356), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_473), .Y(n_548) );
AO21x1_ASAP7_75t_SL g549 ( .A1(n_515), .A2(n_386), .B(n_323), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_498), .A2(n_386), .B1(n_407), .B2(n_281), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_493), .A2(n_325), .B1(n_375), .B2(n_374), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_485), .A2(n_325), .B1(n_375), .B2(n_374), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_485), .A2(n_325), .B1(n_375), .B2(n_407), .Y(n_553) );
AND2x2_ASAP7_75t_SL g554 ( .A(n_514), .B(n_390), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_480), .B(n_369), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_511), .B(n_177), .C(n_169), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_483), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_516), .A2(n_325), .B1(n_375), .B2(n_334), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_461), .A2(n_325), .B1(n_375), .B2(n_334), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_483), .B(n_369), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_474), .A2(n_304), .B1(n_326), .B2(n_308), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_488), .B(n_398), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_462), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_514), .A2(n_398), .B1(n_395), .B2(n_390), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_514), .A2(n_339), .B1(n_366), .B2(n_390), .Y(n_566) );
OAI222xp33_ASAP7_75t_L g567 ( .A1(n_471), .A2(n_352), .B1(n_339), .B2(n_366), .C1(n_304), .C2(n_308), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_488), .B(n_352), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_521), .A2(n_325), .B1(n_375), .B2(n_334), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_492), .B(n_390), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_464), .A2(n_366), .B1(n_395), .B2(n_390), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_513), .B(n_177), .C(n_169), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_474), .A2(n_325), .B1(n_334), .B2(n_335), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_505), .A2(n_334), .B1(n_335), .B2(n_366), .Y(n_574) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_470), .B(n_177), .C(n_169), .Y(n_575) );
OAI222xp33_ASAP7_75t_L g576 ( .A1(n_489), .A2(n_339), .B1(n_308), .B2(n_301), .C1(n_295), .C2(n_343), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_482), .A2(n_335), .B1(n_176), .B2(n_339), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_503), .A2(n_335), .B1(n_176), .B2(n_339), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_500), .A2(n_398), .B1(n_395), .B2(n_390), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_464), .A2(n_398), .B1(n_395), .B2(n_390), .Y(n_580) );
AOI222xp33_ASAP7_75t_L g581 ( .A1(n_460), .A2(n_336), .B1(n_301), .B2(n_295), .C1(n_176), .C2(n_177), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_520), .A2(n_335), .B1(n_176), .B2(n_390), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_492), .B(n_390), .Y(n_583) );
OAI222xp33_ASAP7_75t_L g584 ( .A1(n_489), .A2(n_322), .B1(n_323), .B2(n_343), .C1(n_370), .C2(n_336), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_490), .A2(n_176), .B1(n_395), .B2(n_398), .Y(n_585) );
INVx3_ASAP7_75t_L g586 ( .A(n_523), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_500), .A2(n_398), .B1(n_395), .B2(n_322), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_481), .A2(n_370), .B1(n_312), .B2(n_330), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_524), .A2(n_176), .B1(n_395), .B2(n_398), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_502), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_506), .A2(n_398), .B1(n_395), .B2(n_318), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_497), .A2(n_330), .B1(n_169), .B2(n_177), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_484), .A2(n_330), .B1(n_177), .B2(n_376), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_502), .B(n_177), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g595 ( .A1(n_519), .A2(n_321), .B1(n_298), .B2(n_340), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_478), .A2(n_321), .B1(n_298), .B2(n_318), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_501), .A2(n_340), .B1(n_300), .B2(n_376), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_523), .B(n_324), .Y(n_598) );
OAI222xp33_ASAP7_75t_L g599 ( .A1(n_517), .A2(n_351), .B1(n_324), .B2(n_340), .C1(n_300), .C2(n_306), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_484), .A2(n_177), .B1(n_351), .B2(n_342), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_523), .A2(n_324), .B1(n_300), .B2(n_321), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_469), .A2(n_177), .B1(n_342), .B2(n_345), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g603 ( .A1(n_456), .A2(n_324), .B1(n_306), .B2(n_245), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_477), .A2(n_342), .B1(n_345), .B2(n_329), .Y(n_604) );
BUFx2_ASAP7_75t_L g605 ( .A(n_518), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_456), .A2(n_296), .B1(n_345), .B2(n_341), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_486), .B(n_162), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_508), .A2(n_329), .B1(n_332), .B2(n_327), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_472), .A2(n_329), .B1(n_296), .B2(n_314), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_475), .A2(n_329), .B1(n_332), .B2(n_327), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_507), .A2(n_332), .B1(n_327), .B2(n_296), .Y(n_611) );
AOI222xp33_ASAP7_75t_L g612 ( .A1(n_472), .A2(n_235), .B1(n_327), .B2(n_162), .C1(n_242), .C2(n_338), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_522), .A2(n_338), .B1(n_162), .B2(n_341), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_522), .A2(n_338), .B1(n_341), .B2(n_315), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_510), .A2(n_315), .B1(n_314), .B2(n_310), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_491), .A2(n_315), .B1(n_314), .B2(n_310), .Y(n_616) );
BUFx2_ASAP7_75t_L g617 ( .A(n_491), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_495), .A2(n_310), .B1(n_160), .B2(n_161), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_564), .B(n_495), .Y(n_619) );
AND2x2_ASAP7_75t_SL g620 ( .A(n_554), .B(n_504), .Y(n_620) );
OAI221xp5_ASAP7_75t_SL g621 ( .A1(n_537), .A2(n_504), .B1(n_234), .B2(n_19), .C(n_21), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_536), .B(n_160), .Y(n_622) );
OAI221xp5_ASAP7_75t_SL g623 ( .A1(n_562), .A2(n_17), .B1(n_18), .B2(n_19), .C(n_22), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_536), .B(n_160), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_532), .B(n_18), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_532), .B(n_160), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_542), .B(n_22), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_554), .B(n_160), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_542), .B(n_23), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_563), .B(n_160), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_572), .B(n_164), .C(n_161), .Y(n_631) );
OAI221xp5_ASAP7_75t_SL g632 ( .A1(n_562), .A2(n_23), .B1(n_24), .B2(n_25), .C(n_26), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_548), .B(n_25), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_546), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_548), .B(n_27), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_556), .B(n_27), .Y(n_636) );
OA21x2_ASAP7_75t_L g637 ( .A1(n_598), .A2(n_309), .B(n_216), .Y(n_637) );
AOI21xp5_ASAP7_75t_SL g638 ( .A1(n_571), .A2(n_28), .B(n_29), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_556), .B(n_30), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_558), .B(n_31), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_558), .B(n_31), .Y(n_641) );
AOI211xp5_ASAP7_75t_L g642 ( .A1(n_606), .A2(n_164), .B(n_161), .C(n_160), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_605), .B(n_32), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_557), .B(n_164), .C(n_161), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_533), .B(n_164), .C(n_161), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_590), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_527), .A2(n_160), .B1(n_161), .B2(n_164), .C(n_167), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_525), .B(n_32), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_541), .B(n_33), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_531), .A2(n_167), .B1(n_309), .B2(n_35), .Y(n_650) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_595), .A2(n_164), .B1(n_161), .B2(n_160), .C(n_167), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_576), .A2(n_164), .B1(n_161), .B2(n_167), .C(n_35), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_605), .B(n_545), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_541), .B(n_33), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_545), .B(n_34), .Y(n_655) );
NOR2xp33_ASAP7_75t_R g656 ( .A(n_586), .B(n_34), .Y(n_656) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_575), .A2(n_167), .B(n_309), .Y(n_657) );
OAI21xp5_ASAP7_75t_SL g658 ( .A1(n_528), .A2(n_540), .B(n_609), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_565), .B(n_161), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_579), .B(n_164), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_590), .B(n_164), .Y(n_661) );
OAI21xp5_ASAP7_75t_SL g662 ( .A1(n_567), .A2(n_164), .B(n_213), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_617), .B(n_167), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_581), .B(n_214), .C(n_213), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_607), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_535), .B(n_39), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_612), .B(n_214), .C(n_211), .Y(n_667) );
NAND2xp33_ASAP7_75t_R g668 ( .A(n_531), .B(n_40), .Y(n_668) );
AND2x2_ASAP7_75t_SL g669 ( .A(n_531), .B(n_42), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_534), .A2(n_526), .B1(n_543), .B2(n_616), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_539), .B(n_44), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_580), .B(n_214), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_570), .B(n_45), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_588), .B(n_48), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_588), .B(n_49), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_607), .B(n_214), .C(n_221), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_547), .A2(n_214), .B1(n_221), .B2(n_216), .Y(n_677) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_584), .A2(n_50), .B(n_52), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_598), .B(n_226), .C(n_220), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_549), .B(n_54), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_583), .B(n_55), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_549), .B(n_56), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_594), .B(n_58), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_553), .A2(n_226), .B1(n_220), .B2(n_65), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_555), .B(n_61), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_529), .A2(n_274), .B1(n_251), .B2(n_241), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_594), .B(n_62), .Y(n_687) );
OA21x2_ASAP7_75t_L g688 ( .A1(n_568), .A2(n_274), .B(n_251), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_561), .B(n_68), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_591), .B(n_69), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_597), .B(n_538), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_552), .B(n_70), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_587), .B(n_72), .C(n_73), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_611), .B(n_75), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_592), .B(n_76), .C(n_77), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_608), .B(n_78), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_529), .B(n_80), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_544), .B(n_81), .C(n_83), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_550), .A2(n_84), .B1(n_86), .B2(n_90), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_585), .B(n_91), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_596), .B(n_92), .Y(n_701) );
OAI21xp5_ASAP7_75t_SL g702 ( .A1(n_599), .A2(n_93), .B(n_94), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_614), .B(n_95), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_582), .A2(n_241), .B1(n_239), .B2(n_238), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_603), .A2(n_239), .B1(n_238), .B2(n_232), .C(n_199), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_566), .A2(n_224), .B(n_212), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_589), .B(n_96), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_593), .B(n_97), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_551), .B(n_101), .C(n_103), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_610), .A2(n_192), .B1(n_200), .B2(n_210), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_613), .B(n_104), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_530), .B(n_107), .Y(n_712) );
OA21x2_ASAP7_75t_L g713 ( .A1(n_600), .A2(n_192), .B(n_200), .Y(n_713) );
AND2x2_ASAP7_75t_SL g714 ( .A(n_574), .B(n_192), .Y(n_714) );
AOI22xp33_ASAP7_75t_SL g715 ( .A1(n_601), .A2(n_224), .B1(n_210), .B2(n_212), .Y(n_715) );
INVx3_ASAP7_75t_L g716 ( .A(n_620), .Y(n_716) );
OA211x2_ASAP7_75t_L g717 ( .A1(n_628), .A2(n_559), .B(n_573), .C(n_604), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_653), .B(n_569), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_619), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_646), .B(n_618), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_634), .B(n_602), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_678), .B(n_577), .C(n_578), .Y(n_722) );
AOI211xp5_ASAP7_75t_L g723 ( .A1(n_658), .A2(n_560), .B(n_615), .C(n_210), .Y(n_723) );
AO21x1_ASAP7_75t_SL g724 ( .A1(n_663), .A2(n_661), .B(n_665), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g725 ( .A(n_638), .B(n_224), .C(n_702), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_625), .B(n_630), .Y(n_726) );
NOR3xp33_ASAP7_75t_L g727 ( .A(n_623), .B(n_632), .C(n_648), .Y(n_727) );
NAND2xp33_ASAP7_75t_SL g728 ( .A(n_656), .B(n_668), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_691), .A2(n_714), .B1(n_670), .B2(n_652), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_662), .A2(n_621), .B(n_669), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_688), .B(n_649), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_688), .B(n_654), .Y(n_732) );
AND2x4_ASAP7_75t_L g733 ( .A(n_672), .B(n_680), .Y(n_733) );
BUFx2_ASAP7_75t_L g734 ( .A(n_656), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_688), .B(n_622), .Y(n_735) );
INVx1_ASAP7_75t_SL g736 ( .A(n_643), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g737 ( .A(n_642), .B(n_668), .C(n_672), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_627), .B(n_629), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_633), .B(n_635), .Y(n_739) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_622), .Y(n_740) );
OA211x2_ASAP7_75t_L g741 ( .A1(n_659), .A2(n_660), .B(n_655), .C(n_693), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_624), .B(n_669), .Y(n_742) );
AOI211xp5_ASAP7_75t_L g743 ( .A1(n_659), .A2(n_667), .B(n_682), .C(n_660), .Y(n_743) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_631), .B(n_636), .C(n_641), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_639), .B(n_640), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_687), .B(n_637), .Y(n_746) );
NOR3xp33_ASAP7_75t_SL g747 ( .A(n_650), .B(n_664), .C(n_651), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_673), .B(n_681), .Y(n_748) );
NAND4xp25_ASAP7_75t_L g749 ( .A(n_670), .B(n_686), .C(n_710), .D(n_697), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_714), .A2(n_696), .B1(n_674), .B2(n_675), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_679), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_666), .B(n_671), .Y(n_752) );
NOR2x1_ASAP7_75t_L g753 ( .A(n_676), .B(n_645), .Y(n_753) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_713), .Y(n_754) );
BUFx2_ASAP7_75t_L g755 ( .A(n_713), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_644), .B(n_699), .C(n_698), .Y(n_756) );
AND2x4_ASAP7_75t_SL g757 ( .A(n_683), .B(n_696), .Y(n_757) );
AND2x4_ASAP7_75t_L g758 ( .A(n_690), .B(n_657), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_690), .B(n_700), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_685), .B(n_689), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_701), .B(n_686), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g762 ( .A(n_647), .B(n_709), .C(n_692), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_712), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_694), .B(n_706), .Y(n_764) );
OR2x2_ASAP7_75t_L g765 ( .A(n_703), .B(n_704), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_708), .B(n_700), .Y(n_766) );
AO21x2_ASAP7_75t_L g767 ( .A1(n_684), .A2(n_695), .B(n_707), .Y(n_767) );
NOR2x1_ASAP7_75t_L g768 ( .A(n_711), .B(n_715), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_704), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_705), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_677), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_653), .B(n_634), .Y(n_772) );
NOR3xp33_ASAP7_75t_L g773 ( .A(n_623), .B(n_632), .C(n_425), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g774 ( .A(n_658), .B(n_678), .C(n_564), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_691), .A2(n_658), .B1(n_457), .B2(n_678), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_653), .B(n_634), .Y(n_776) );
NOR3xp33_ASAP7_75t_L g777 ( .A(n_623), .B(n_632), .C(n_425), .Y(n_777) );
NAND3xp33_ASAP7_75t_L g778 ( .A(n_658), .B(n_678), .C(n_564), .Y(n_778) );
OR2x2_ASAP7_75t_L g779 ( .A(n_619), .B(n_564), .Y(n_779) );
AO21x2_ASAP7_75t_L g780 ( .A1(n_661), .A2(n_626), .B(n_630), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_653), .B(n_634), .Y(n_781) );
AO21x2_ASAP7_75t_L g782 ( .A1(n_661), .A2(n_626), .B(n_630), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_772), .B(n_776), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_780), .Y(n_784) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_779), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_775), .B(n_774), .Y(n_786) );
AND2x4_ASAP7_75t_SL g787 ( .A(n_733), .B(n_740), .Y(n_787) );
BUFx2_ASAP7_75t_L g788 ( .A(n_781), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_780), .B(n_782), .Y(n_789) );
OR2x2_ASAP7_75t_L g790 ( .A(n_719), .B(n_735), .Y(n_790) );
OR2x2_ASAP7_75t_L g791 ( .A(n_735), .B(n_782), .Y(n_791) );
NAND4xp75_ASAP7_75t_L g792 ( .A(n_717), .B(n_741), .C(n_730), .D(n_768), .Y(n_792) );
XOR2x2_ASAP7_75t_L g793 ( .A(n_778), .B(n_734), .Y(n_793) );
NAND4xp75_ASAP7_75t_L g794 ( .A(n_730), .B(n_747), .C(n_721), .D(n_750), .Y(n_794) );
INVx1_ASAP7_75t_SL g795 ( .A(n_726), .Y(n_795) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_731), .Y(n_796) );
XNOR2x2_ASAP7_75t_L g797 ( .A(n_737), .B(n_749), .Y(n_797) );
INVx2_ASAP7_75t_SL g798 ( .A(n_733), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_736), .B(n_738), .Y(n_799) );
NOR3xp33_ASAP7_75t_L g800 ( .A(n_762), .B(n_756), .C(n_744), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_739), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_732), .Y(n_802) );
NAND4xp75_ASAP7_75t_SL g803 ( .A(n_728), .B(n_742), .C(n_746), .D(n_759), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_720), .Y(n_804) );
XNOR2xp5_ASAP7_75t_L g805 ( .A(n_729), .B(n_718), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_720), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_716), .B(n_755), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_754), .B(n_724), .Y(n_808) );
INVx2_ASAP7_75t_SL g809 ( .A(n_757), .Y(n_809) );
INVx2_ASAP7_75t_SL g810 ( .A(n_753), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_771), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_763), .B(n_745), .Y(n_812) );
XOR2x2_ASAP7_75t_L g813 ( .A(n_773), .B(n_777), .Y(n_813) );
NAND4xp75_ASAP7_75t_L g814 ( .A(n_761), .B(n_752), .C(n_764), .D(n_760), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_769), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_761), .B(n_758), .Y(n_816) );
XNOR2xp5_ASAP7_75t_L g817 ( .A(n_723), .B(n_777), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_758), .B(n_751), .Y(n_818) );
CKINVDCx5p33_ASAP7_75t_R g819 ( .A(n_760), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_748), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_765), .Y(n_821) );
XOR2x2_ASAP7_75t_L g822 ( .A(n_773), .B(n_725), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_821), .B(n_748), .Y(n_823) );
INVx1_ASAP7_75t_SL g824 ( .A(n_787), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_790), .Y(n_825) );
INVxp67_ASAP7_75t_L g826 ( .A(n_786), .Y(n_826) );
XOR2x2_ASAP7_75t_L g827 ( .A(n_813), .B(n_727), .Y(n_827) );
XNOR2x1_ASAP7_75t_L g828 ( .A(n_813), .B(n_770), .Y(n_828) );
XNOR2xp5_ASAP7_75t_L g829 ( .A(n_822), .B(n_727), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_790), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_791), .Y(n_831) );
NOR2x1_ASAP7_75t_L g832 ( .A(n_792), .B(n_767), .Y(n_832) );
XOR2x2_ASAP7_75t_L g833 ( .A(n_794), .B(n_743), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_802), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_796), .Y(n_835) );
INVxp67_ASAP7_75t_L g836 ( .A(n_786), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_791), .Y(n_837) );
XNOR2xp5_ASAP7_75t_L g838 ( .A(n_822), .B(n_722), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_801), .Y(n_839) );
INVx1_ASAP7_75t_SL g840 ( .A(n_787), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_820), .Y(n_841) );
XOR2x2_ASAP7_75t_L g842 ( .A(n_797), .B(n_766), .Y(n_842) );
INVx2_ASAP7_75t_SL g843 ( .A(n_808), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_784), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_785), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_784), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_823), .Y(n_847) );
AOI22x1_ASAP7_75t_L g848 ( .A1(n_838), .A2(n_810), .B1(n_817), .B2(n_797), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_823), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_824), .A2(n_809), .B1(n_788), .B2(n_798), .Y(n_850) );
INVx1_ASAP7_75t_SL g851 ( .A(n_840), .Y(n_851) );
OA22x2_ASAP7_75t_L g852 ( .A1(n_829), .A2(n_805), .B1(n_810), .B2(n_809), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_845), .Y(n_853) );
AO22x1_ASAP7_75t_L g854 ( .A1(n_832), .A2(n_800), .B1(n_808), .B2(n_819), .Y(n_854) );
AO22x2_ASAP7_75t_L g855 ( .A1(n_843), .A2(n_803), .B1(n_814), .B2(n_811), .Y(n_855) );
OAI22x1_ASAP7_75t_L g856 ( .A1(n_838), .A2(n_819), .B1(n_798), .B2(n_821), .Y(n_856) );
OA22x2_ASAP7_75t_L g857 ( .A1(n_829), .A2(n_793), .B1(n_789), .B2(n_816), .Y(n_857) );
INVx1_ASAP7_75t_SL g858 ( .A(n_843), .Y(n_858) );
AOI22x1_ASAP7_75t_L g859 ( .A1(n_833), .A2(n_793), .B1(n_807), .B2(n_815), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_835), .Y(n_860) );
AOI22x1_ASAP7_75t_SL g861 ( .A1(n_827), .A2(n_806), .B1(n_804), .B2(n_795), .Y(n_861) );
INVx1_ASAP7_75t_SL g862 ( .A(n_827), .Y(n_862) );
INVx2_ASAP7_75t_L g863 ( .A(n_851), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_857), .A2(n_833), .B1(n_842), .B2(n_826), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_851), .Y(n_865) );
OAI322xp33_ASAP7_75t_L g866 ( .A1(n_862), .A2(n_836), .A3(n_828), .B1(n_837), .B2(n_831), .C1(n_835), .C2(n_812), .Y(n_866) );
BUFx2_ASAP7_75t_L g867 ( .A(n_858), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_853), .Y(n_868) );
INVxp67_ASAP7_75t_L g869 ( .A(n_848), .Y(n_869) );
NOR2x1_ASAP7_75t_SL g870 ( .A(n_850), .B(n_825), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_852), .A2(n_842), .B1(n_828), .B2(n_818), .Y(n_871) );
OAI22x1_ASAP7_75t_L g872 ( .A1(n_864), .A2(n_859), .B1(n_862), .B2(n_858), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_865), .Y(n_873) );
OA22x2_ASAP7_75t_L g874 ( .A1(n_871), .A2(n_856), .B1(n_861), .B2(n_854), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_863), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g876 ( .A1(n_869), .A2(n_855), .B1(n_860), .B2(n_849), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_875), .Y(n_877) );
A2O1A1Ixp33_ASAP7_75t_L g878 ( .A1(n_876), .A2(n_867), .B(n_868), .C(n_866), .Y(n_878) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_874), .A2(n_855), .B1(n_831), .B2(n_837), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_877), .Y(n_880) );
NAND2x1_ASAP7_75t_L g881 ( .A(n_879), .B(n_873), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_878), .B(n_872), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_882), .A2(n_812), .B1(n_866), .B2(n_799), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_881), .B(n_870), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_883), .Y(n_885) );
NOR2xp67_ASAP7_75t_L g886 ( .A(n_884), .B(n_880), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_885), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_886), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_887), .A2(n_846), .B1(n_844), .B2(n_847), .Y(n_889) );
INVx4_ASAP7_75t_L g890 ( .A(n_889), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_890), .A2(n_887), .B1(n_888), .B2(n_799), .Y(n_891) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_891), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_892), .A2(n_830), .B1(n_839), .B2(n_825), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_893), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g895 ( .A1(n_894), .A2(n_830), .B1(n_844), .B2(n_846), .C(n_834), .Y(n_895) );
AOI211xp5_ASAP7_75t_L g896 ( .A1(n_895), .A2(n_834), .B(n_783), .C(n_841), .Y(n_896) );
endmodule