module fake_netlist_5_2209_n_962 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_962);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_962;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_318;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_785;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_523;
wire n_268;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_372;
wire n_443;
wire n_677;
wire n_244;
wire n_293;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_247;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_946;
wire n_417;
wire n_932;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_624;
wire n_252;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_568;
wire n_509;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_448;
wire n_259;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_795;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_696;
wire n_255;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_580;
wire n_290;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_928;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_834;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_425;
wire n_237;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_832;
wire n_695;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_404;
wire n_233;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_565;
wire n_426;
wire n_566;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_960;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx2_ASAP7_75t_SL g198 ( 
.A(n_196),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_84),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_1),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_119),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_70),
.Y(n_205)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_110),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_136),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_38),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_180),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_160),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_64),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_197),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_51),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_65),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_57),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_13),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_14),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_171),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_68),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_105),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_120),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_135),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_151),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_111),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_10),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_155),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_97),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_83),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_96),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_159),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_162),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_45),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_185),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_116),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_17),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_126),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_112),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_161),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_21),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_147),
.Y(n_244)
);

CKINVDCx12_ASAP7_75t_R g245 ( 
.A(n_91),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_67),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_163),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_85),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_8),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_154),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_134),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_53),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_78),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_15),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_157),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_59),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_175),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_145),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_121),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_124),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_167),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_191),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_5),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_34),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_19),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_178),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_61),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_50),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_72),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_54),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_26),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_73),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_75),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_156),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_79),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_47),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_25),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_118),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_130),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_127),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_169),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_165),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_173),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_184),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_98),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_142),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_86),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_13),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_23),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_101),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_6),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_21),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_82),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_52),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_33),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_1),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_158),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_93),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_77),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_177),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_58),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_187),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_168),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_226),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_213),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_283),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_277),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_277),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_202),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_277),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_218),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_214),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_243),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_221),
.Y(n_315)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_238),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_256),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_199),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_241),
.Y(n_320)
);

INVxp33_ASAP7_75t_SL g321 ( 
.A(n_249),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_288),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_212),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_212),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_296),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_263),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_240),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_271),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_201),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_254),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_203),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_240),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_200),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_214),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_204),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_207),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_208),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_289),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_209),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_215),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_205),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_216),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_227),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_210),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_292),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_258),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_231),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_235),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_239),
.Y(n_350)
);

INVxp33_ASAP7_75t_SL g351 ( 
.A(n_217),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_246),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_250),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_264),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_278),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_270),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_272),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_274),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_211),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_282),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_287),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_254),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_285),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_291),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_294),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_284),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_299),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_234),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_219),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_220),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_234),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_291),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_222),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_275),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_223),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_347),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_307),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_305),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_308),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_327),
.Y(n_380)
);

OAI21x1_ASAP7_75t_L g381 ( 
.A1(n_320),
.A2(n_279),
.B(n_275),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_313),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_313),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_313),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_309),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_319),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_334),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_326),
.Y(n_389)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_0),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_336),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_330),
.Y(n_394)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_335),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_338),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_332),
.B(n_198),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_342),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_345),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_335),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

AND2x2_ASAP7_75t_SL g402 ( 
.A(n_304),
.B(n_279),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_335),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_340),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_335),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_343),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

NAND2x1p5_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_244),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_324),
.B(n_286),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_371),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_325),
.B(n_286),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_348),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_347),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_328),
.B(n_295),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_320),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_349),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_350),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_322),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_352),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_354),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_359),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_356),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_357),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_355),
.A2(n_273),
.B1(n_266),
.B2(n_300),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_333),
.B(n_273),
.Y(n_430)
);

AND2x6_ASAP7_75t_L g431 ( 
.A(n_322),
.B(n_214),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_329),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_362),
.Y(n_433)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_374),
.A2(n_295),
.B(n_206),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_418),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_406),
.B(n_369),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_418),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_388),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_421),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_421),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_421),
.Y(n_443)
);

INVx8_ASAP7_75t_L g444 ( 
.A(n_386),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_391),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_402),
.A2(n_306),
.B1(n_364),
.B2(n_363),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_397),
.B(n_316),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_389),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_402),
.A2(n_365),
.B1(n_367),
.B2(n_331),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_384),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_377),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_331),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_392),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_378),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_392),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_403),
.B(n_370),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_403),
.B(n_373),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_428),
.A2(n_321),
.B1(n_375),
.B2(n_339),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_400),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_378),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_400),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_362),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_409),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_409),
.Y(n_467)
);

NOR3xp33_ASAP7_75t_L g468 ( 
.A(n_416),
.B(n_323),
.C(n_310),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_412),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_376),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_412),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_410),
.B(n_312),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_383),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_403),
.B(n_224),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_383),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_393),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_379),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_431),
.B(n_241),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_435),
.B(n_396),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_434),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_410),
.B(n_351),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_434),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_383),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_387),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_386),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_404),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_381),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_411),
.B(n_314),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_L g492 ( 
.A(n_431),
.B(n_241),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_405),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_407),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_425),
.B(n_329),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_425),
.B(n_339),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_435),
.B(n_225),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_383),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_380),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_435),
.B(n_228),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_381),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_395),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_434),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_411),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_376),
.A2(n_366),
.B1(n_318),
.B2(n_315),
.Y(n_505)
);

INVxp33_ASAP7_75t_SL g506 ( 
.A(n_394),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_425),
.B(n_346),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_453),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_504),
.B(n_435),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_503),
.B(n_394),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_438),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_438),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_439),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_503),
.B(n_398),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_L g515 ( 
.A(n_504),
.B(n_398),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_454),
.B(n_435),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_454),
.B(n_399),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_480),
.B(n_399),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_447),
.B(n_414),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_439),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_491),
.B(n_415),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_465),
.B(n_419),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_486),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_465),
.A2(n_346),
.B1(n_366),
.B2(n_411),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_448),
.B(n_380),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_486),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_453),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_477),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_480),
.B(n_214),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_480),
.B(n_241),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_477),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_472),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_483),
.B(n_472),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_483),
.B(n_241),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_450),
.B(n_401),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_459),
.A2(n_422),
.B(n_420),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_444),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_466),
.Y(n_538)
);

NOR3xp33_ASAP7_75t_L g539 ( 
.A(n_482),
.B(n_432),
.C(n_401),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_483),
.B(n_423),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_441),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_507),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_479),
.B(n_229),
.Y(n_543)
);

INVxp33_ASAP7_75t_L g544 ( 
.A(n_505),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_481),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_441),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_490),
.A2(n_413),
.B1(n_417),
.B2(n_390),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_481),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_442),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_446),
.B(n_432),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_491),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_442),
.B(n_230),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_487),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_440),
.B(n_424),
.Y(n_554)
);

BUFx12f_ASAP7_75t_SL g555 ( 
.A(n_506),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_485),
.B(n_413),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_445),
.B(n_426),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_442),
.B(n_232),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_487),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_444),
.B(n_413),
.Y(n_560)
);

BUFx8_ASAP7_75t_L g561 ( 
.A(n_476),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_489),
.B(n_427),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_449),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_493),
.B(n_429),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_494),
.B(n_417),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_460),
.B(n_233),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_436),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_466),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_467),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_461),
.A2(n_417),
.B1(n_236),
.B2(n_269),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_495),
.B(n_433),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_437),
.B(n_237),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_L g573 ( 
.A(n_497),
.B(n_500),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_506),
.B(n_287),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_501),
.B(n_467),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_501),
.B(n_469),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_469),
.B(n_431),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_471),
.B(n_431),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_474),
.B(n_242),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_471),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_523),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_538),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_567),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_525),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_516),
.B(n_436),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_568),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_526),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_572),
.B(n_443),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_538),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_555),
.Y(n_591)
);

O2A1O1Ixp33_ASAP7_75t_L g592 ( 
.A1(n_510),
.A2(n_478),
.B(n_492),
.C(n_490),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_517),
.B(n_488),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_572),
.B(n_443),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_533),
.A2(n_478),
.B1(n_492),
.B2(n_390),
.Y(n_595)
);

BUFx4f_ASAP7_75t_L g596 ( 
.A(n_560),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_523),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_518),
.B(n_488),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_533),
.A2(n_518),
.B1(n_514),
.B2(n_510),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_571),
.B(n_496),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_526),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_542),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_519),
.B(n_473),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_561),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_523),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_569),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_580),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_522),
.B(n_473),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_535),
.Y(n_609)
);

OR2x2_ASAP7_75t_SL g610 ( 
.A(n_574),
.B(n_470),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_561),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_514),
.A2(n_499),
.B1(n_468),
.B2(n_444),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_508),
.B(n_475),
.Y(n_613)
);

INVxp67_ASAP7_75t_SL g614 ( 
.A(n_523),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_527),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_563),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_550),
.B(n_444),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_537),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_521),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_528),
.B(n_531),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_545),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_524),
.B(n_457),
.Y(n_622)
);

A2O1A1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_565),
.A2(n_317),
.B(n_455),
.C(n_449),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_521),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_551),
.B(n_457),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_548),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_537),
.Y(n_627)
);

INVxp67_ASAP7_75t_SL g628 ( 
.A(n_575),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_553),
.B(n_475),
.Y(n_629)
);

AND2x4_ASAP7_75t_SL g630 ( 
.A(n_560),
.B(n_470),
.Y(n_630)
);

BUFx4f_ASAP7_75t_SL g631 ( 
.A(n_552),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_R g632 ( 
.A(n_515),
.B(n_463),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_559),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_556),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_540),
.B(n_463),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_579),
.B(n_565),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_563),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_579),
.A2(n_552),
.B1(n_558),
.B2(n_543),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_560),
.Y(n_639)
);

OA22x2_ASAP7_75t_L g640 ( 
.A1(n_602),
.A2(n_570),
.B1(n_544),
.B2(n_554),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_615),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_636),
.B(n_547),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_621),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_600),
.B(n_544),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_583),
.Y(n_645)
);

BUFx8_ASAP7_75t_L g646 ( 
.A(n_604),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_635),
.B(n_547),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_635),
.B(n_557),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_618),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_597),
.Y(n_650)
);

AOI221xp5_ASAP7_75t_L g651 ( 
.A1(n_622),
.A2(n_609),
.B1(n_595),
.B2(n_539),
.C(n_593),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_585),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_593),
.B(n_562),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_622),
.B(n_634),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_618),
.B(n_549),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_617),
.B(n_564),
.Y(n_656)
);

O2A1O1Ixp5_ASAP7_75t_L g657 ( 
.A1(n_598),
.A2(n_529),
.B(n_558),
.C(n_534),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_639),
.B(n_536),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_597),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_595),
.A2(n_529),
.B1(n_509),
.B2(n_576),
.Y(n_660)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_614),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_586),
.A2(n_573),
.B(n_575),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_590),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_599),
.A2(n_576),
.B1(n_530),
.B2(n_534),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_617),
.A2(n_566),
.B1(n_543),
.B2(n_530),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_589),
.A2(n_594),
.B(n_592),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_625),
.B(n_610),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_581),
.B(n_511),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_592),
.A2(n_578),
.B(n_577),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_614),
.A2(n_513),
.B(n_512),
.Y(n_670)
);

O2A1O1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_598),
.A2(n_546),
.B(n_541),
.C(n_520),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_582),
.A2(n_498),
.B(n_484),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_626),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_633),
.Y(n_674)
);

CKINVDCx8_ASAP7_75t_R g675 ( 
.A(n_591),
.Y(n_675)
);

O2A1O1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_620),
.A2(n_456),
.B(n_451),
.C(n_452),
.Y(n_676)
);

O2A1O1Ixp5_ASAP7_75t_SL g677 ( 
.A1(n_587),
.A2(n_502),
.B(n_433),
.C(n_245),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_581),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_603),
.B(n_451),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_582),
.A2(n_498),
.B(n_484),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_597),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_631),
.B(n_612),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_606),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_661),
.Y(n_684)
);

OA21x2_ASAP7_75t_L g685 ( 
.A1(n_666),
.A2(n_623),
.B(n_638),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_652),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_657),
.A2(n_623),
.B(n_608),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_669),
.A2(n_629),
.B(n_613),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_662),
.A2(n_582),
.B(n_628),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_664),
.A2(n_628),
.B(n_607),
.Y(n_690)
);

OAI21x1_ASAP7_75t_L g691 ( 
.A1(n_672),
.A2(n_584),
.B(n_588),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_644),
.B(n_619),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_641),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_651),
.B(n_632),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_643),
.Y(n_695)
);

AO31x2_ASAP7_75t_L g696 ( 
.A1(n_660),
.A2(n_637),
.A3(n_616),
.B(n_458),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_675),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_673),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_677),
.A2(n_455),
.B(n_452),
.Y(n_699)
);

CKINVDCx11_ASAP7_75t_R g700 ( 
.A(n_649),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_656),
.A2(n_582),
.B(n_588),
.Y(n_701)
);

AND3x4_ASAP7_75t_L g702 ( 
.A(n_658),
.B(n_611),
.C(n_624),
.Y(n_702)
);

AOI221x1_ASAP7_75t_L g703 ( 
.A1(n_682),
.A2(n_605),
.B1(n_601),
.B2(n_597),
.C(n_458),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_642),
.B(n_630),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_646),
.Y(n_705)
);

AO32x2_ASAP7_75t_L g706 ( 
.A1(n_647),
.A2(n_640),
.A3(n_653),
.B1(n_631),
.B2(n_648),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_658),
.B(n_618),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_665),
.A2(n_601),
.B(n_596),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_674),
.B(n_605),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_654),
.B(n_678),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_667),
.Y(n_711)
);

OAI21x1_ASAP7_75t_L g712 ( 
.A1(n_680),
.A2(n_462),
.B(n_456),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_646),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_683),
.B(n_618),
.Y(n_714)
);

CKINVDCx11_ASAP7_75t_R g715 ( 
.A(n_649),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_649),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_668),
.B(n_627),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_671),
.A2(n_596),
.B(n_627),
.C(n_464),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_650),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_679),
.A2(n_627),
.B(n_464),
.Y(n_720)
);

OAI22x1_ASAP7_75t_L g721 ( 
.A1(n_645),
.A2(n_632),
.B1(n_268),
.B2(n_267),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_663),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_670),
.A2(n_462),
.B(n_502),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_681),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_650),
.B(n_627),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_676),
.A2(n_502),
.B(n_248),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_690),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_697),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_693),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_695),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_698),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_707),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_694),
.A2(n_681),
.B1(n_659),
.B2(n_655),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_684),
.B(n_659),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_692),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_704),
.B(n_247),
.Y(n_736)
);

BUFx2_ASAP7_75t_SL g737 ( 
.A(n_710),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_696),
.Y(n_738)
);

OAI21x1_ASAP7_75t_L g739 ( 
.A1(n_689),
.A2(n_433),
.B(n_395),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_711),
.A2(n_276),
.B1(n_303),
.B2(n_302),
.Y(n_740)
);

OAI21x1_ASAP7_75t_L g741 ( 
.A1(n_688),
.A2(n_395),
.B(n_28),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_717),
.B(n_251),
.Y(n_742)
);

OAI21x1_ASAP7_75t_SL g743 ( 
.A1(n_708),
.A2(n_0),
.B(n_2),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_722),
.Y(n_744)
);

OAI21x1_ASAP7_75t_L g745 ( 
.A1(n_712),
.A2(n_29),
.B(n_27),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_686),
.B(n_702),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_714),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_747)
);

AOI221xp5_ASAP7_75t_L g748 ( 
.A1(n_721),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.C(n_261),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_709),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_723),
.A2(n_103),
.B(n_195),
.Y(n_750)
);

OAI21x1_ASAP7_75t_SL g751 ( 
.A1(n_708),
.A2(n_2),
.B(n_3),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_685),
.A2(n_293),
.B1(n_301),
.B2(n_298),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_709),
.Y(n_753)
);

BUFx2_ASAP7_75t_R g754 ( 
.A(n_705),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_687),
.A2(n_262),
.B(n_297),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_714),
.Y(n_756)
);

AO31x2_ASAP7_75t_L g757 ( 
.A1(n_703),
.A2(n_431),
.A3(n_4),
.B(n_5),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_691),
.A2(n_100),
.B(n_193),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_687),
.A2(n_99),
.B(n_192),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_707),
.B(n_30),
.Y(n_760)
);

INVx3_ASAP7_75t_SL g761 ( 
.A(n_713),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_719),
.Y(n_762)
);

OAI21x1_ASAP7_75t_L g763 ( 
.A1(n_720),
.A2(n_95),
.B(n_190),
.Y(n_763)
);

OAI21x1_ASAP7_75t_L g764 ( 
.A1(n_720),
.A2(n_94),
.B(n_189),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_719),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_725),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_699),
.A2(n_92),
.B(n_188),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_699),
.A2(n_90),
.B(n_186),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_685),
.B(n_280),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_701),
.A2(n_89),
.B(n_183),
.Y(n_770)
);

AO21x2_ASAP7_75t_L g771 ( 
.A1(n_718),
.A2(n_431),
.B(n_290),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_726),
.A2(n_281),
.B(n_4),
.C(n_6),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_716),
.B(n_31),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_766),
.B(n_696),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_735),
.B(n_706),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_752),
.A2(n_706),
.B1(n_724),
.B2(n_726),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_756),
.B(n_700),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_SL g778 ( 
.A1(n_773),
.A2(n_715),
.B(n_706),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_729),
.Y(n_779)
);

AOI21x1_ASAP7_75t_SL g780 ( 
.A1(n_769),
.A2(n_734),
.B(n_760),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_SL g781 ( 
.A1(n_773),
.A2(n_88),
.B(n_181),
.Y(n_781)
);

NAND2x1p5_ASAP7_75t_L g782 ( 
.A(n_762),
.B(n_696),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_752),
.A2(n_87),
.B(n_179),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_744),
.Y(n_784)
);

AOI21x1_ASAP7_75t_SL g785 ( 
.A1(n_769),
.A2(n_3),
.B(n_7),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_737),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_732),
.B(n_32),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_772),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_SL g789 ( 
.A1(n_773),
.A2(n_104),
.B(n_176),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_765),
.Y(n_790)
);

OA21x2_ASAP7_75t_L g791 ( 
.A1(n_767),
.A2(n_9),
.B(n_10),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_730),
.B(n_731),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_746),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_793)
);

AOI21x1_ASAP7_75t_SL g794 ( 
.A1(n_734),
.A2(n_11),
.B(n_12),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_732),
.B(n_35),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_760),
.B(n_36),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_SL g797 ( 
.A1(n_742),
.A2(n_108),
.B(n_174),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_740),
.A2(n_748),
.B1(n_736),
.B2(n_733),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_749),
.B(n_753),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_SL g800 ( 
.A1(n_748),
.A2(n_107),
.B(n_172),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_755),
.A2(n_106),
.B(n_166),
.Y(n_801)
);

AND2x6_ASAP7_75t_L g802 ( 
.A(n_743),
.B(n_37),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_738),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_761),
.Y(n_804)
);

OA21x2_ASAP7_75t_L g805 ( 
.A1(n_768),
.A2(n_15),
.B(n_16),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_755),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_738),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_740),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_757),
.B(n_20),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_747),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_754),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_774),
.Y(n_812)
);

AO21x1_ASAP7_75t_SL g813 ( 
.A1(n_809),
.A2(n_727),
.B(n_757),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_804),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_784),
.B(n_727),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_775),
.B(n_741),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_780),
.A2(n_739),
.B(n_758),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_782),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_782),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_807),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_792),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_779),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_803),
.Y(n_823)
);

NOR2x1_ASAP7_75t_R g824 ( 
.A(n_804),
.B(n_796),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_790),
.B(n_757),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_799),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_804),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_791),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_791),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_805),
.Y(n_830)
);

OAI21x1_ASAP7_75t_L g831 ( 
.A1(n_776),
.A2(n_750),
.B(n_764),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_805),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_776),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_802),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_778),
.B(n_759),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_SL g836 ( 
.A1(n_806),
.A2(n_771),
.B(n_747),
.Y(n_836)
);

OA21x2_ASAP7_75t_L g837 ( 
.A1(n_801),
.A2(n_751),
.B(n_745),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_820),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_821),
.B(n_777),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_820),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_821),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_822),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_821),
.B(n_771),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_816),
.B(n_786),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_818),
.B(n_819),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_822),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_823),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_822),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_826),
.B(n_798),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_823),
.B(n_810),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_826),
.B(n_810),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_818),
.B(n_763),
.Y(n_852)
);

AO21x2_ASAP7_75t_L g853 ( 
.A1(n_828),
.A2(n_783),
.B(n_800),
.Y(n_853)
);

NAND5xp2_ASAP7_75t_SL g854 ( 
.A(n_844),
.B(n_814),
.C(n_835),
.D(n_788),
.E(n_825),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_838),
.Y(n_855)
);

AOI221xp5_ASAP7_75t_L g856 ( 
.A1(n_849),
.A2(n_811),
.B1(n_793),
.B2(n_808),
.C(n_836),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_838),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_841),
.B(n_823),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_842),
.Y(n_859)
);

AOI31xp33_ASAP7_75t_L g860 ( 
.A1(n_844),
.A2(n_824),
.A3(n_835),
.B(n_851),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_839),
.Y(n_861)
);

AO21x2_ASAP7_75t_L g862 ( 
.A1(n_846),
.A2(n_830),
.B(n_828),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_SL g863 ( 
.A1(n_853),
.A2(n_834),
.B1(n_833),
.B2(n_825),
.Y(n_863)
);

OAI33xp33_ASAP7_75t_L g864 ( 
.A1(n_850),
.A2(n_830),
.A3(n_812),
.B1(n_833),
.B2(n_832),
.B3(n_829),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_839),
.B(n_816),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_855),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_858),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_857),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_862),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_861),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_865),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_867),
.B(n_861),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_868),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_870),
.B(n_863),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_871),
.B(n_850),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_869),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_866),
.B(n_863),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_876),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_875),
.B(n_866),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_874),
.B(n_860),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_876),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_877),
.A2(n_856),
.B1(n_834),
.B2(n_854),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_879),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_878),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_882),
.A2(n_872),
.B1(n_834),
.B2(n_873),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_880),
.B(n_827),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_881),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_884),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_883),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_887),
.A2(n_827),
.B(n_832),
.C(n_829),
.Y(n_890)
);

OAI221xp5_ASAP7_75t_L g891 ( 
.A1(n_885),
.A2(n_761),
.B1(n_797),
.B2(n_836),
.C(n_781),
.Y(n_891)
);

OAI32xp33_ASAP7_75t_L g892 ( 
.A1(n_886),
.A2(n_829),
.A3(n_832),
.B1(n_864),
.B2(n_819),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_889),
.B(n_888),
.Y(n_893)
);

NOR2x1p5_ASAP7_75t_L g894 ( 
.A(n_891),
.B(n_754),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_890),
.B(n_862),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_892),
.B(n_728),
.Y(n_896)
);

NOR2x1_ASAP7_75t_L g897 ( 
.A(n_888),
.B(n_789),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_889),
.A2(n_853),
.B1(n_864),
.B2(n_843),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_889),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_889),
.B(n_859),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_L g901 ( 
.A(n_899),
.B(n_26),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_893),
.B(n_859),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_900),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_896),
.Y(n_904)
);

OAI21xp33_ASAP7_75t_L g905 ( 
.A1(n_897),
.A2(n_843),
.B(n_845),
.Y(n_905)
);

AOI211xp5_ASAP7_75t_L g906 ( 
.A1(n_895),
.A2(n_824),
.B(n_796),
.C(n_787),
.Y(n_906)
);

AOI221xp5_ASAP7_75t_L g907 ( 
.A1(n_898),
.A2(n_853),
.B1(n_840),
.B2(n_847),
.C(n_841),
.Y(n_907)
);

AOI221xp5_ASAP7_75t_L g908 ( 
.A1(n_894),
.A2(n_840),
.B1(n_847),
.B2(n_846),
.C(n_845),
.Y(n_908)
);

OAI221xp5_ASAP7_75t_SL g909 ( 
.A1(n_898),
.A2(n_818),
.B1(n_819),
.B2(n_812),
.C(n_842),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_897),
.A2(n_802),
.B(n_831),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_SL g911 ( 
.A1(n_904),
.A2(n_794),
.B(n_785),
.C(n_848),
.Y(n_911)
);

OAI221xp5_ASAP7_75t_L g912 ( 
.A1(n_906),
.A2(n_837),
.B1(n_848),
.B2(n_795),
.C(n_802),
.Y(n_912)
);

XNOR2xp5_ASAP7_75t_L g913 ( 
.A(n_901),
.B(n_852),
.Y(n_913)
);

AOI221xp5_ASAP7_75t_L g914 ( 
.A1(n_903),
.A2(n_845),
.B1(n_852),
.B2(n_816),
.C(n_815),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_908),
.A2(n_802),
.B1(n_845),
.B2(n_852),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_SL g916 ( 
.A1(n_910),
.A2(n_816),
.B(n_815),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_902),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_905),
.Y(n_918)
);

AOI221x1_ASAP7_75t_L g919 ( 
.A1(n_909),
.A2(n_815),
.B1(n_40),
.B2(n_41),
.C(n_42),
.Y(n_919)
);

OAI22xp33_ASAP7_75t_L g920 ( 
.A1(n_907),
.A2(n_837),
.B1(n_815),
.B2(n_813),
.Y(n_920)
);

NOR3xp33_ASAP7_75t_L g921 ( 
.A(n_917),
.B(n_770),
.C(n_831),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_918),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_913),
.B(n_837),
.Y(n_923)
);

NOR2xp67_ASAP7_75t_SL g924 ( 
.A(n_912),
.B(n_916),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_911),
.Y(n_925)
);

NOR2x1p5_ASAP7_75t_L g926 ( 
.A(n_919),
.B(n_39),
.Y(n_926)
);

OAI31xp33_ASAP7_75t_SL g927 ( 
.A1(n_920),
.A2(n_817),
.A3(n_813),
.B(n_837),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_915),
.B(n_43),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_914),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_918),
.B(n_44),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_922),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_SL g932 ( 
.A1(n_925),
.A2(n_817),
.B1(n_49),
.B2(n_55),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_929),
.B(n_48),
.Y(n_933)
);

OAI211xp5_ASAP7_75t_SL g934 ( 
.A1(n_930),
.A2(n_928),
.B(n_927),
.C(n_923),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_926),
.Y(n_935)
);

NOR2x1_ASAP7_75t_L g936 ( 
.A(n_924),
.B(n_56),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_921),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_922),
.Y(n_938)
);

NAND2x1p5_ASAP7_75t_L g939 ( 
.A(n_936),
.B(n_60),
.Y(n_939)
);

NOR2x1_ASAP7_75t_L g940 ( 
.A(n_938),
.B(n_62),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_935),
.Y(n_941)
);

NOR3x1_ASAP7_75t_L g942 ( 
.A(n_931),
.B(n_63),
.C(n_66),
.Y(n_942)
);

AOI21x1_ASAP7_75t_L g943 ( 
.A1(n_937),
.A2(n_69),
.B(n_71),
.Y(n_943)
);

NOR2x1_ASAP7_75t_L g944 ( 
.A(n_940),
.B(n_933),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_939),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_942),
.Y(n_946)
);

NOR3x1_ASAP7_75t_L g947 ( 
.A(n_941),
.B(n_934),
.C(n_943),
.Y(n_947)
);

AOI221xp5_ASAP7_75t_L g948 ( 
.A1(n_946),
.A2(n_932),
.B1(n_76),
.B2(n_80),
.C(n_81),
.Y(n_948)
);

OAI221xp5_ASAP7_75t_L g949 ( 
.A1(n_944),
.A2(n_74),
.B1(n_102),
.B2(n_109),
.C(n_113),
.Y(n_949)
);

XNOR2x1_ASAP7_75t_L g950 ( 
.A(n_948),
.B(n_947),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_949),
.B(n_945),
.Y(n_951)
);

XNOR2xp5_ASAP7_75t_L g952 ( 
.A(n_950),
.B(n_114),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_951),
.A2(n_115),
.B1(n_117),
.B2(n_122),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_953),
.A2(n_123),
.B1(n_125),
.B2(n_128),
.Y(n_954)
);

OR3x2_ASAP7_75t_L g955 ( 
.A(n_952),
.B(n_129),
.C(n_131),
.Y(n_955)
);

XOR2xp5_ASAP7_75t_L g956 ( 
.A(n_955),
.B(n_133),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_954),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_R g958 ( 
.A1(n_957),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_958),
.B(n_956),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_959),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_960),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_961)
);

AOI211xp5_ASAP7_75t_L g962 ( 
.A1(n_961),
.A2(n_150),
.B(n_152),
.C(n_153),
.Y(n_962)
);


endmodule