module fake_jpeg_26293_n_108 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp67_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_24),
.Y(n_48)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_22),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_37),
.C(n_28),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_53),
.C(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_42),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_17),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_15),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_15),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_35),
.B1(n_29),
.B2(n_33),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_68),
.Y(n_74)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_23),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_23),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_21),
.B1(n_35),
.B2(n_3),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_1),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_61),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_67),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_41),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_56),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_54),
.B(n_40),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_68),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_74),
.B(n_78),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_81),
.C(n_70),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_73),
.B1(n_74),
.B2(n_41),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_49),
.B1(n_62),
.B2(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_86),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_43),
.B(n_49),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_79),
.C(n_72),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_91),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_10),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_80),
.B(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_97),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_2),
.B(n_6),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_9),
.B(n_10),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_101),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_99),
.B(n_96),
.CI(n_93),
.CON(n_102),
.SN(n_102)
);

NAND2xp33_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_46),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_104),
.B(n_103),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_104),
.Y(n_108)
);


endmodule