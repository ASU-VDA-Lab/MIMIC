module real_aes_17648_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_887;
wire n_187;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
wire n_862;
AND2x4_ASAP7_75t_L g880 ( .A(n_0), .B(n_881), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_1), .A2(n_3), .B1(n_216), .B2(n_217), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_2), .A2(n_46), .B1(n_181), .B2(n_199), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_4), .A2(n_25), .B1(n_199), .B2(n_255), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_5), .A2(n_17), .B1(n_512), .B2(n_541), .Y(n_540) );
AOI22x1_ASAP7_75t_SL g845 ( .A1(n_6), .A2(n_78), .B1(n_846), .B2(n_847), .Y(n_845) );
INVxp67_ASAP7_75t_SL g847 ( .A(n_6), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_7), .A2(n_63), .B1(n_145), .B2(n_146), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_8), .A2(n_18), .B1(n_181), .B2(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g881 ( .A(n_9), .Y(n_881) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_10), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_11), .Y(n_553) );
AOI22x1_ASAP7_75t_L g110 ( .A1(n_12), .A2(n_111), .B1(n_112), .B2(n_115), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_12), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_13), .A2(n_19), .B1(n_530), .B2(n_531), .Y(n_529) );
OR2x2_ASAP7_75t_L g835 ( .A(n_14), .B(n_40), .Y(n_835) );
BUFx2_ASAP7_75t_L g884 ( .A(n_14), .Y(n_884) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_15), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_16), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_20), .A2(n_102), .B1(n_217), .B2(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_21), .A2(n_39), .B1(n_138), .B2(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_22), .B(n_136), .Y(n_554) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_23), .A2(n_60), .B(n_151), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_24), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_26), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_27), .B(n_133), .Y(n_227) );
INVx4_ASAP7_75t_R g168 ( .A(n_28), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_29), .A2(n_49), .B1(n_185), .B2(n_214), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_30), .A2(n_55), .B1(n_185), .B2(n_512), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_31), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_32), .B(n_539), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_33), .Y(n_566) );
INVx1_ASAP7_75t_L g222 ( .A(n_34), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_35), .B(n_199), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_SL g269 ( .A1(n_36), .A2(n_132), .B(n_181), .C(n_270), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_37), .A2(n_56), .B1(n_181), .B2(n_185), .Y(n_256) );
XOR2xp5_ASAP7_75t_L g841 ( .A(n_38), .B(n_188), .Y(n_841) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_40), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g108 ( .A1(n_41), .A2(n_109), .B1(n_110), .B2(n_116), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_41), .Y(n_109) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_41), .A2(n_109), .B1(n_110), .B2(n_116), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_42), .A2(n_90), .B1(n_181), .B2(n_582), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g862 ( .A(n_43), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_44), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_45), .A2(n_48), .B1(n_181), .B2(n_182), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_47), .A2(n_61), .B1(n_512), .B2(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g231 ( .A(n_50), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_51), .B(n_181), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_52), .Y(n_197) );
INVx2_ASAP7_75t_L g830 ( .A(n_53), .Y(n_830) );
BUFx3_ASAP7_75t_L g833 ( .A(n_54), .Y(n_833) );
INVx1_ASAP7_75t_L g855 ( .A(n_54), .Y(n_855) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_57), .A2(n_861), .B(n_866), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_58), .A2(n_91), .B1(n_181), .B2(n_185), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_59), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_62), .A2(n_105), .B1(n_873), .B2(n_887), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_64), .A2(n_79), .B1(n_214), .B2(n_514), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_65), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_66), .A2(n_82), .B1(n_181), .B2(n_182), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_67), .A2(n_100), .B1(n_512), .B2(n_531), .Y(n_563) );
INVx1_ASAP7_75t_L g151 ( .A(n_68), .Y(n_151) );
AND2x4_ASAP7_75t_L g154 ( .A(n_69), .B(n_155), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_70), .A2(n_93), .B1(n_185), .B2(n_214), .Y(n_213) );
AO22x1_ASAP7_75t_L g134 ( .A1(n_71), .A2(n_80), .B1(n_135), .B2(n_138), .Y(n_134) );
OAI22x1_ASAP7_75t_SL g112 ( .A1(n_72), .A2(n_74), .B1(n_113), .B2(n_114), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_72), .Y(n_113) );
INVx1_ASAP7_75t_L g155 ( .A(n_73), .Y(n_155) );
INVx1_ASAP7_75t_L g114 ( .A(n_74), .Y(n_114) );
AND2x2_ASAP7_75t_L g272 ( .A(n_75), .B(n_193), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_76), .B(n_145), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_77), .Y(n_265) );
INVx1_ASAP7_75t_L g846 ( .A(n_78), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_81), .B(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_84), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_85), .B(n_193), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_86), .A2(n_101), .B1(n_145), .B2(n_185), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_87), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_88), .B(n_149), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_89), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_92), .B(n_193), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_94), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_95), .B(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g122 ( .A(n_96), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_96), .B(n_854), .Y(n_853) );
NAND2xp33_ASAP7_75t_L g557 ( .A(n_97), .B(n_136), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g162 ( .A1(n_98), .A2(n_145), .B(n_163), .C(n_165), .Y(n_162) );
AND2x2_ASAP7_75t_L g175 ( .A(n_99), .B(n_176), .Y(n_175) );
NAND2xp33_ASAP7_75t_L g203 ( .A(n_103), .B(n_169), .Y(n_203) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_836), .Y(n_105) );
AOI21xp33_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_825), .B(n_827), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_117), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_110), .Y(n_116) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g825 ( .A(n_118), .B(n_826), .Y(n_825) );
OA22x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_123), .B1(n_500), .B2(n_822), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx8_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g871 ( .A(n_121), .B(n_872), .Y(n_871) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g824 ( .A(n_122), .Y(n_824) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_399), .Y(n_123) );
AND3x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_317), .C(n_376), .Y(n_124) );
AOI221xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_208), .B1(n_236), .B2(n_289), .C(n_292), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_189), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_156), .Y(n_128) );
INVx2_ASAP7_75t_L g247 ( .A(n_129), .Y(n_247) );
AND2x2_ASAP7_75t_L g304 ( .A(n_129), .B(n_246), .Y(n_304) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g397 ( .A(n_130), .B(n_332), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_130), .B(n_178), .Y(n_461) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_134), .B(n_140), .C(n_152), .Y(n_131) );
INVx6_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_132), .A2(n_203), .B(n_204), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_132), .B(n_134), .Y(n_286) );
O2A1O1Ixp5_ASAP7_75t_L g552 ( .A1(n_132), .A2(n_182), .B(n_553), .C(n_554), .Y(n_552) );
BUFx8_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g143 ( .A(n_133), .Y(n_143) );
INVx1_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
INVx1_ASAP7_75t_L g230 ( .A(n_133), .Y(n_230) );
INVxp67_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
INVx3_ASAP7_75t_L g512 ( .A(n_136), .Y(n_512) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g139 ( .A(n_137), .Y(n_139) );
INVx1_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_137), .Y(n_147) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
INVx3_ASAP7_75t_L g181 ( .A(n_137), .Y(n_181) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_137), .Y(n_185) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_137), .Y(n_199) );
INVx1_ASAP7_75t_L g218 ( .A(n_137), .Y(n_218) );
INVx2_ASAP7_75t_L g255 ( .A(n_137), .Y(n_255) );
OAI21xp33_ASAP7_75t_SL g226 ( .A1(n_138), .A2(n_227), .B(n_228), .Y(n_226) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g285 ( .A(n_140), .Y(n_285) );
OAI21x1_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_144), .B(n_148), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_141), .A2(n_233), .B(n_234), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_141), .A2(n_183), .B1(n_254), .B2(n_256), .Y(n_253) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g515 ( .A(n_142), .Y(n_515) );
BUFx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g201 ( .A(n_143), .Y(n_201) );
INVx1_ASAP7_75t_L g530 ( .A(n_146), .Y(n_530) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_147), .B(n_164), .Y(n_163) );
OAI21xp33_ASAP7_75t_L g152 ( .A1(n_148), .A2(n_149), .B(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
INVx2_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
INVx2_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
INVx1_ASAP7_75t_L g287 ( .A(n_152), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_153), .A2(n_263), .B(n_269), .Y(n_262) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx10_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
BUFx10_ASAP7_75t_L g207 ( .A(n_154), .Y(n_207) );
INVx1_ASAP7_75t_L g220 ( .A(n_154), .Y(n_220) );
INVx2_ASAP7_75t_L g336 ( .A(n_156), .Y(n_336) );
OR2x2_ASAP7_75t_L g425 ( .A(n_156), .B(n_342), .Y(n_425) );
OR2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_178), .Y(n_156) );
INVx1_ASAP7_75t_L g240 ( .A(n_157), .Y(n_240) );
INVx2_ASAP7_75t_L g327 ( .A(n_157), .Y(n_327) );
AND2x2_ASAP7_75t_L g351 ( .A(n_157), .B(n_178), .Y(n_351) );
AND2x4_ASAP7_75t_L g364 ( .A(n_157), .B(n_284), .Y(n_364) );
AND2x2_ASAP7_75t_L g381 ( .A(n_157), .B(n_243), .Y(n_381) );
AND2x2_ASAP7_75t_L g391 ( .A(n_157), .B(n_283), .Y(n_391) );
AND2x2_ASAP7_75t_L g419 ( .A(n_157), .B(n_191), .Y(n_419) );
AO21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_161), .B(n_175), .Y(n_157) );
AO31x2_ASAP7_75t_L g508 ( .A1(n_158), .A2(n_509), .A3(n_510), .B(n_516), .Y(n_508) );
AO31x2_ASAP7_75t_L g519 ( .A1(n_158), .A2(n_219), .A3(n_520), .B(n_523), .Y(n_519) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_SL g534 ( .A(n_160), .B(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_160), .B(n_585), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_166), .B(n_173), .Y(n_161) );
INVx1_ASAP7_75t_L g172 ( .A(n_165), .Y(n_172) );
INVx1_ASAP7_75t_SL g533 ( .A(n_165), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_167), .B(n_172), .Y(n_166) );
OAI22xp33_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_167) );
INVx2_ASAP7_75t_L g214 ( .A(n_169), .Y(n_214) );
INVx1_ASAP7_75t_L g539 ( .A(n_169), .Y(n_539) );
INVx1_ASAP7_75t_L g541 ( .A(n_170), .Y(n_541) );
OAI22x1_ASAP7_75t_L g179 ( .A1(n_172), .A2(n_180), .B1(n_183), .B2(n_184), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_172), .A2(n_183), .B1(n_213), .B2(n_215), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_172), .A2(n_183), .B1(n_581), .B2(n_583), .Y(n_580) );
INVx1_ASAP7_75t_L g509 ( .A(n_173), .Y(n_509) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AO31x2_ASAP7_75t_L g178 ( .A1(n_174), .A2(n_179), .A3(n_186), .B(n_187), .Y(n_178) );
AO31x2_ASAP7_75t_L g527 ( .A1(n_174), .A2(n_211), .A3(n_528), .B(n_534), .Y(n_527) );
AO31x2_ASAP7_75t_L g536 ( .A1(n_174), .A2(n_537), .A3(n_542), .B(n_543), .Y(n_536) );
AO31x2_ASAP7_75t_L g596 ( .A1(n_174), .A2(n_257), .A3(n_597), .B(n_600), .Y(n_596) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_177), .B(n_188), .Y(n_187) );
BUFx2_ASAP7_75t_L g211 ( .A(n_177), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_177), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_177), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g246 ( .A(n_178), .Y(n_246) );
AND2x2_ASAP7_75t_L g288 ( .A(n_178), .B(n_191), .Y(n_288) );
INVx2_ASAP7_75t_L g332 ( .A(n_178), .Y(n_332) );
AND2x2_ASAP7_75t_L g464 ( .A(n_178), .B(n_327), .Y(n_464) );
INVx4_ASAP7_75t_L g182 ( .A(n_181), .Y(n_182) );
INVx1_ASAP7_75t_L g514 ( .A(n_181), .Y(n_514) );
INVx1_ASAP7_75t_L g531 ( .A(n_181), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_182), .A2(n_197), .B(n_198), .C(n_200), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_183), .A2(n_511), .B1(n_513), .B2(n_515), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_183), .A2(n_515), .B1(n_521), .B2(n_522), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_183), .A2(n_529), .B1(n_532), .B2(n_533), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_183), .A2(n_515), .B1(n_538), .B2(n_540), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_183), .A2(n_556), .B(n_557), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_183), .A2(n_533), .B1(n_563), .B2(n_564), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_183), .A2(n_515), .B1(n_598), .B2(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g216 ( .A(n_185), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_185), .B(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_186), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_186), .B(n_524), .Y(n_523) );
AND3x1_ASAP7_75t_L g300 ( .A(n_189), .B(n_240), .C(n_301), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_189), .B(n_304), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_189), .B(n_464), .Y(n_481) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
BUFx2_ASAP7_75t_L g385 ( .A(n_190), .Y(n_385) );
AND2x2_ASAP7_75t_L g494 ( .A(n_190), .B(n_276), .Y(n_494) );
BUFx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g243 ( .A(n_191), .Y(n_243) );
AND2x2_ASAP7_75t_L g245 ( .A(n_191), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g333 ( .A(n_191), .Y(n_333) );
NAND2x1p5_ASAP7_75t_L g191 ( .A(n_192), .B(n_195), .Y(n_191) );
NOR2x1_ASAP7_75t_L g205 ( .A(n_193), .B(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g257 ( .A(n_193), .Y(n_257) );
INVx4_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g235 ( .A(n_194), .B(n_207), .Y(n_235) );
BUFx3_ASAP7_75t_L g542 ( .A(n_194), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_194), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g550 ( .A(n_194), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_194), .B(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_194), .B(n_601), .Y(n_600) );
OAI21x1_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_202), .B(n_205), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_199), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AO31x2_ASAP7_75t_L g252 ( .A1(n_207), .A2(n_253), .A3(n_257), .B(n_258), .Y(n_252) );
BUFx2_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g360 ( .A(n_209), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g467 ( .A(n_209), .B(n_357), .Y(n_467) );
AND2x2_ASAP7_75t_L g474 ( .A(n_209), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_223), .Y(n_209) );
INVx1_ASAP7_75t_L g291 ( .A(n_210), .Y(n_291) );
INVx1_ASAP7_75t_L g309 ( .A(n_210), .Y(n_309) );
OR2x2_ASAP7_75t_L g313 ( .A(n_210), .B(n_252), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_210), .B(n_252), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_210), .B(n_278), .Y(n_339) );
INVx1_ASAP7_75t_L g411 ( .A(n_210), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_210), .B(n_260), .Y(n_470) );
AO31x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .A3(n_219), .B(n_221), .Y(n_210) );
AOI21x1_ASAP7_75t_L g261 ( .A1(n_211), .A2(n_262), .B(n_272), .Y(n_261) );
AO31x2_ASAP7_75t_L g561 ( .A1(n_211), .A2(n_509), .A3(n_562), .B(n_565), .Y(n_561) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_218), .B(n_267), .Y(n_266) );
AO31x2_ASAP7_75t_L g579 ( .A1(n_219), .A2(n_542), .A3(n_580), .B(n_584), .Y(n_579) );
INVx2_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_SL g558 ( .A(n_220), .Y(n_558) );
OR2x2_ASAP7_75t_L g308 ( .A(n_223), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_223), .B(n_276), .Y(n_315) );
INVx3_ASAP7_75t_L g323 ( .A(n_223), .Y(n_323) );
NAND2x1p5_ASAP7_75t_SL g348 ( .A(n_223), .B(n_322), .Y(n_348) );
BUFx2_ASAP7_75t_L g370 ( .A(n_223), .Y(n_370) );
INVx1_ASAP7_75t_L g375 ( .A(n_223), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_223), .B(n_411), .Y(n_428) );
AND2x4_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_232), .B(n_235), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
BUFx4f_ASAP7_75t_L g268 ( .A(n_230), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_273), .Y(n_236) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_244), .B(n_248), .Y(n_237) );
INVxp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g306 ( .A(n_240), .Y(n_306) );
INVx1_ASAP7_75t_L g398 ( .A(n_240), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_241), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g434 ( .A(n_241), .B(n_351), .Y(n_434) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g446 ( .A(n_242), .B(n_364), .Y(n_446) );
BUFx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g350 ( .A(n_243), .B(n_283), .Y(n_350) );
AND2x2_ASAP7_75t_L g390 ( .A(n_243), .B(n_332), .Y(n_390) );
AND2x4_ASAP7_75t_SL g244 ( .A(n_245), .B(n_247), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_245), .B(n_326), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_245), .B(n_364), .Y(n_373) );
AND2x2_ASAP7_75t_L g413 ( .A(n_245), .B(n_406), .Y(n_413) );
INVx1_ASAP7_75t_L g430 ( .A(n_246), .Y(n_430) );
OAI322xp33_ASAP7_75t_L g292 ( .A1(n_247), .A2(n_293), .A3(n_299), .B1(n_302), .B2(n_307), .C1(n_311), .C2(n_316), .Y(n_292) );
AOI32xp33_ASAP7_75t_L g383 ( .A1(n_247), .A2(n_343), .A3(n_384), .B1(n_386), .B2(n_388), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_247), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g471 ( .A(n_247), .B(n_390), .Y(n_471) );
INVxp67_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g310 ( .A(n_251), .Y(n_310) );
AND2x2_ASAP7_75t_L g374 ( .A(n_251), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g448 ( .A(n_251), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_251), .B(n_410), .Y(n_449) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_260), .Y(n_251) );
INVx2_ASAP7_75t_SL g278 ( .A(n_252), .Y(n_278) );
BUFx2_ASAP7_75t_L g296 ( .A(n_252), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_255), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_SL g582 ( .A(n_255), .Y(n_582) );
INVx2_ASAP7_75t_L g322 ( .A(n_260), .Y(n_322) );
OR2x2_ASAP7_75t_L g358 ( .A(n_260), .B(n_278), .Y(n_358) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g276 ( .A(n_261), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_266), .B(n_268), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_279), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g475 ( .A(n_275), .Y(n_475) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_276), .B(n_323), .Y(n_338) );
INVxp67_ASAP7_75t_L g345 ( .A(n_276), .Y(n_345) );
OR2x2_ASAP7_75t_L g415 ( .A(n_277), .B(n_322), .Y(n_415) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_288), .Y(n_280) );
AND2x2_ASAP7_75t_L g335 ( .A(n_281), .B(n_336), .Y(n_335) );
NOR2x1_ASAP7_75t_L g498 ( .A(n_281), .B(n_333), .Y(n_498) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g406 ( .A(n_282), .Y(n_406) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g326 ( .A(n_283), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g431 ( .A(n_284), .B(n_327), .Y(n_431) );
AOI21x1_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B(n_287), .Y(n_284) );
INVx2_ASAP7_75t_L g367 ( .A(n_288), .Y(n_367) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g298 ( .A(n_291), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
INVx1_ASAP7_75t_L g371 ( .A(n_294), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_294), .B(n_410), .Y(n_479) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_295), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g438 ( .A(n_295), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g347 ( .A(n_298), .B(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_298), .B(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g343 ( .A(n_308), .Y(n_343) );
INVx1_ASAP7_75t_L g439 ( .A(n_308), .Y(n_439) );
INVx1_ASAP7_75t_L g489 ( .A(n_308), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_312), .B(n_362), .Y(n_394) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g379 ( .A(n_313), .Y(n_379) );
OR2x2_ASAP7_75t_L g387 ( .A(n_313), .B(n_348), .Y(n_387) );
OR2x2_ASAP7_75t_L g455 ( .A(n_313), .B(n_362), .Y(n_455) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g403 ( .A(n_315), .B(n_320), .Y(n_403) );
INVx1_ASAP7_75t_L g486 ( .A(n_316), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_352), .Y(n_317) );
OAI321xp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_324), .A3(n_328), .B1(n_334), .B2(n_337), .C(n_340), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_319), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g362 ( .A(n_322), .Y(n_362) );
AND2x4_ASAP7_75t_L g410 ( .A(n_323), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g414 ( .A(n_323), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_325), .B(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI211xp5_ASAP7_75t_L g420 ( .A1(n_329), .A2(n_421), .B(n_424), .C(n_426), .Y(n_420) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g418 ( .A(n_331), .Y(n_418) );
INVx1_ASAP7_75t_L g452 ( .A(n_331), .Y(n_452) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g342 ( .A(n_333), .Y(n_342) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g341 ( .A(n_336), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_337), .B(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_338), .Y(n_442) );
AOI32xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .A3(n_344), .B1(n_346), .B2(n_349), .Y(n_340) );
OR2x2_ASAP7_75t_L g496 ( .A(n_342), .B(n_397), .Y(n_496) );
AND2x2_ASAP7_75t_L g377 ( .A(n_344), .B(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g422 ( .A(n_345), .B(n_423), .Y(n_422) );
NAND2x1_ASAP7_75t_L g488 ( .A(n_345), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
AND2x2_ASAP7_75t_L g468 ( .A(n_350), .B(n_464), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_351), .B(n_406), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_351), .A2(n_378), .B1(n_474), .B2(n_476), .Y(n_473) );
OAI221xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_359), .B2(n_363), .C(n_365), .Y(n_352) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g409 ( .A(n_357), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g499 ( .A(n_361), .B(n_378), .Y(n_499) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx3_ASAP7_75t_L g369 ( .A(n_364), .Y(n_369) );
AND2x2_ASAP7_75t_L g476 ( .A(n_364), .B(n_418), .Y(n_476) );
AOI32xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_370), .A3(n_371), .B1(n_372), .B2(n_374), .Y(n_365) );
NOR2xp33_ASAP7_75t_SL g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g378 ( .A(n_375), .B(n_379), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_380), .B(n_382), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g392 ( .A1(n_378), .A2(n_393), .B(n_395), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g491 ( .A1(n_378), .A2(n_492), .B(n_495), .Y(n_491) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_392), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AND2x2_ASAP7_75t_L g490 ( .A(n_391), .B(n_452), .Y(n_490) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
NOR4xp75_ASAP7_75t_L g399 ( .A(n_400), .B(n_432), .C(n_456), .D(n_482), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_420), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B(n_407), .Y(n_401) );
INVx2_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_405), .A2(n_445), .B1(n_447), .B2(n_449), .Y(n_444) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_412), .B1(n_414), .B2(n_416), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_408), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g423 ( .A(n_410), .Y(n_423) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_417), .A2(n_498), .B(n_499), .Y(n_497) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_425), .A2(n_451), .B(n_453), .Y(n_450) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
OR2x2_ASAP7_75t_L g447 ( .A(n_428), .B(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g443 ( .A(n_429), .Y(n_443) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B(n_440), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI211xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_443), .B(n_444), .C(n_450), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g465 ( .A(n_447), .Y(n_465) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2x1_ASAP7_75t_SL g456 ( .A(n_457), .B(n_472), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_466), .Y(n_457) );
OAI21xp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_462), .B(n_465), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B1(n_469), .B2(n_471), .Y(n_466) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_477), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_474), .A2(n_486), .B1(n_487), .B2(n_490), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_497), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_491), .Y(n_484) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_500), .A2(n_844), .B1(n_845), .B2(n_848), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_500), .Y(n_844) );
AND3x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_719), .C(n_797), .Y(n_500) );
NOR2x1_ASAP7_75t_L g501 ( .A(n_502), .B(n_662), .Y(n_501) );
NAND3xp33_ASAP7_75t_L g502 ( .A(n_503), .B(n_609), .C(n_632), .Y(n_502) );
AOI221x1_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_545), .B1(n_567), .B2(n_576), .C(n_586), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_525), .Y(n_504) );
AND2x4_ASAP7_75t_L g699 ( .A(n_505), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
INVx2_ASAP7_75t_L g658 ( .A(n_507), .Y(n_658) );
INVx1_ASAP7_75t_L g685 ( .A(n_507), .Y(n_685) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g570 ( .A(n_508), .Y(n_570) );
AND2x4_ASAP7_75t_L g636 ( .A(n_508), .B(n_571), .Y(n_636) );
INVx1_ASAP7_75t_L g718 ( .A(n_518), .Y(n_718) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g571 ( .A(n_519), .Y(n_571) );
AND2x4_ASAP7_75t_L g607 ( .A(n_519), .B(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g627 ( .A(n_519), .B(n_536), .Y(n_627) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_519), .Y(n_679) );
INVx1_ASAP7_75t_L g772 ( .A(n_519), .Y(n_772) );
AND2x2_ASAP7_75t_L g818 ( .A(n_519), .B(n_527), .Y(n_818) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_526), .B(n_684), .Y(n_683) );
NAND2x1_ASAP7_75t_L g688 ( .A(n_526), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g812 ( .A(n_526), .B(n_710), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_526), .B(n_766), .Y(n_816) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_536), .Y(n_526) );
INVx4_ASAP7_75t_SL g573 ( .A(n_527), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_527), .B(n_575), .Y(n_620) );
BUFx2_ASAP7_75t_L g704 ( .A(n_527), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_527), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g575 ( .A(n_536), .Y(n_575) );
INVx2_ASAP7_75t_L g608 ( .A(n_536), .Y(n_608) );
AND2x2_ASAP7_75t_L g610 ( .A(n_536), .B(n_570), .Y(n_610) );
INVx1_ASAP7_75t_L g635 ( .A(n_536), .Y(n_635) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_536), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_536), .B(n_718), .Y(n_749) );
INVxp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g793 ( .A(n_547), .B(n_794), .Y(n_793) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_560), .Y(n_547) );
AND2x4_ASAP7_75t_L g590 ( .A(n_548), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g650 ( .A(n_548), .B(n_595), .Y(n_650) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx2_ASAP7_75t_L g736 ( .A(n_549), .Y(n_736) );
OAI21x1_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B(n_559), .Y(n_549) );
OAI21x1_ASAP7_75t_L g623 ( .A1(n_550), .A2(n_551), .B(n_559), .Y(n_623) );
OAI21x1_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_555), .B(n_558), .Y(n_551) );
AND2x4_ASAP7_75t_L g648 ( .A(n_560), .B(n_579), .Y(n_648) );
INVx3_ASAP7_75t_L g671 ( .A(n_560), .Y(n_671) );
INVx2_ASAP7_75t_L g692 ( .A(n_560), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_560), .B(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_560), .B(n_594), .Y(n_786) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g578 ( .A(n_561), .B(n_579), .Y(n_578) );
BUFx2_ASAP7_75t_L g589 ( .A(n_561), .Y(n_589) );
AND2x2_ASAP7_75t_L g665 ( .A(n_561), .B(n_591), .Y(n_665) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx3_ASAP7_75t_L g643 ( .A(n_570), .Y(n_643) );
AND2x2_ASAP7_75t_L g678 ( .A(n_570), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g747 ( .A(n_570), .B(n_573), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_571), .B(n_573), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g709 ( .A(n_572), .B(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx2_ASAP7_75t_L g606 ( .A(n_573), .Y(n_606) );
AND2x2_ASAP7_75t_L g634 ( .A(n_573), .B(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g652 ( .A(n_573), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g694 ( .A(n_573), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_573), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g755 ( .A(n_573), .Y(n_755) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_578), .B(n_622), .Y(n_621) );
AND2x4_ASAP7_75t_SL g629 ( .A(n_578), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g708 ( .A(n_578), .B(n_593), .Y(n_708) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_578), .Y(n_743) );
INVx2_ASAP7_75t_L g760 ( .A(n_578), .Y(n_760) );
INVx2_ASAP7_75t_L g591 ( .A(n_579), .Y(n_591) );
OR2x2_ASAP7_75t_L g640 ( .A(n_579), .B(n_631), .Y(n_640) );
INVx1_ASAP7_75t_L g661 ( .A(n_579), .Y(n_661) );
BUFx2_ASAP7_75t_L g676 ( .A(n_579), .Y(n_676) );
OR2x2_ASAP7_75t_L g745 ( .A(n_579), .B(n_596), .Y(n_745) );
AOI21xp5_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_592), .B(n_603), .Y(n_586) );
O2A1O1Ixp33_ASAP7_75t_L g711 ( .A1(n_587), .A2(n_667), .B(n_712), .C(n_715), .Y(n_711) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g611 ( .A(n_588), .B(n_612), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_588), .A2(n_645), .B1(n_811), .B2(n_812), .Y(n_810) );
AND2x4_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g602 ( .A(n_590), .Y(n_602) );
AND2x4_ASAP7_75t_L g730 ( .A(n_590), .B(n_639), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_590), .B(n_785), .Y(n_784) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_602), .Y(n_592) );
INVx1_ASAP7_75t_L g612 ( .A(n_593), .Y(n_612) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g630 ( .A(n_594), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_595), .B(n_623), .Y(n_673) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g622 ( .A(n_596), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g639 ( .A(n_596), .Y(n_639) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_596), .Y(n_714) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
AND2x2_ASAP7_75t_L g625 ( .A(n_605), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_606), .B(n_685), .Y(n_724) );
INVx2_ASAP7_75t_L g616 ( .A(n_607), .Y(n_616) );
AND2x2_ASAP7_75t_L g693 ( .A(n_607), .B(n_694), .Y(n_693) );
NAND2x1p5_ASAP7_75t_L g738 ( .A(n_607), .B(n_657), .Y(n_738) );
AND2x2_ASAP7_75t_L g775 ( .A(n_607), .B(n_747), .Y(n_775) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B(n_613), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_621), .B1(n_624), .B2(n_628), .Y(n_613) );
NOR2x1_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g819 ( .A(n_616), .Y(n_819) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g659 ( .A(n_622), .Y(n_659) );
AND2x2_ASAP7_75t_L g686 ( .A(n_622), .B(n_671), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_622), .B(n_665), .Y(n_756) );
AND2x4_ASAP7_75t_L g802 ( .A(n_622), .B(n_648), .Y(n_802) );
INVx1_ASAP7_75t_L g631 ( .A(n_623), .Y(n_631) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x4_ASAP7_75t_L g808 ( .A(n_626), .B(n_704), .Y(n_808) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g741 ( .A(n_627), .B(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g769 ( .A(n_627), .B(n_643), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_628), .B(n_801), .Y(n_800) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g750 ( .A(n_630), .B(n_751), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_637), .B1(n_641), .B2(n_645), .C(n_651), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g667 ( .A(n_634), .Y(n_667) );
AND2x2_ASAP7_75t_L g791 ( .A(n_634), .B(n_657), .Y(n_791) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_635), .Y(n_655) );
INVx3_ASAP7_75t_L g653 ( .A(n_636), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_636), .B(n_703), .Y(n_702) );
AND2x4_ASAP7_75t_L g725 ( .A(n_636), .B(n_726), .Y(n_725) );
NOR2xp67_ASAP7_75t_SL g637 ( .A(n_638), .B(n_640), .Y(n_637) );
AND2x2_ASAP7_75t_L g664 ( .A(n_638), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_638), .B(n_671), .Y(n_733) );
AOI322xp5_ASAP7_75t_L g739 ( .A1(n_638), .A2(n_725), .A3(n_740), .B1(n_743), .B2(n_744), .C1(n_746), .C2(n_750), .Y(n_739) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g681 ( .A(n_639), .B(n_648), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_640), .B(n_692), .Y(n_691) );
NOR2x1_ASAP7_75t_L g789 ( .A(n_640), .B(n_790), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_641), .A2(n_783), .B1(n_787), .B2(n_791), .Y(n_782) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx4_ASAP7_75t_L g766 ( .A(n_643), .Y(n_766) );
OR2x2_ASAP7_75t_L g796 ( .A(n_643), .B(n_771), .Y(n_796) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g809 ( .A(n_648), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_649), .B(n_675), .Y(n_696) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI211x1_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B(n_659), .C(n_660), .Y(n_651) );
INVx2_ASAP7_75t_L g689 ( .A(n_653), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g716 ( .A(n_657), .Y(n_716) );
NAND2x1_ASAP7_75t_L g807 ( .A(n_657), .B(n_808), .Y(n_807) );
INVx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g713 ( .A(n_658), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g778 ( .A(n_660), .Y(n_778) );
BUFx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_680), .C(n_695), .Y(n_662) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B(n_668), .C(n_678), .Y(n_663) );
INVx1_ASAP7_75t_L g677 ( .A(n_664), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_665), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g735 ( .A(n_665), .B(n_736), .Y(n_735) );
NAND2xp33_ASAP7_75t_L g758 ( .A(n_665), .B(n_706), .Y(n_758) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_677), .Y(n_668) );
INVx1_ASAP7_75t_L g804 ( .A(n_669), .Y(n_804) );
NAND2x1p5_ASAP7_75t_L g669 ( .A(n_670), .B(n_674), .Y(n_669) );
AND2x4_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx2_ASAP7_75t_L g751 ( .A(n_671), .Y(n_751) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g706 ( .A(n_673), .Y(n_706) );
INVxp67_ASAP7_75t_SL g781 ( .A(n_673), .Y(n_781) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g710 ( .A(n_679), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B1(n_686), .B2(n_687), .C(n_690), .Y(n_680) );
INVxp67_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g742 ( .A(n_685), .Y(n_742) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g728 ( .A(n_692), .Y(n_728) );
NOR2x1p5_ASAP7_75t_L g744 ( .A(n_692), .B(n_745), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_693), .A2(n_732), .B(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g700 ( .A(n_694), .Y(n_700) );
AOI211xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_701), .C(n_711), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_705), .B1(n_707), .B2(n_709), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g790 ( .A(n_714), .Y(n_790) );
OR2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_752), .C(n_773), .Y(n_719) );
NAND3xp33_ASAP7_75t_SL g720 ( .A(n_721), .B(n_731), .C(n_739), .Y(n_720) );
OAI21xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_725), .B(n_727), .Y(n_721) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
AND2x2_ASAP7_75t_L g821 ( .A(n_728), .B(n_789), .Y(n_821) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g767 ( .A1(n_730), .A2(n_768), .B(n_770), .Y(n_767) );
INVxp67_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_737), .Y(n_734) );
OR2x2_ASAP7_75t_L g759 ( .A(n_736), .B(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g794 ( .A(n_745), .Y(n_794) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_748), .Y(n_811) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g754 ( .A(n_749), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g764 ( .A(n_749), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_756), .B1(n_757), .B2(n_761), .C(n_767), .Y(n_752) );
OAI21xp5_ASAP7_75t_L g798 ( .A1(n_753), .A2(n_799), .B(n_803), .Y(n_798) );
BUFx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AOI32xp33_ASAP7_75t_L g792 ( .A1(n_755), .A2(n_766), .A3(n_793), .B1(n_794), .B2(n_795), .Y(n_792) );
AND2x2_ASAP7_75t_SL g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_768), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OAI211xp5_ASAP7_75t_SL g773 ( .A1(n_774), .A2(n_776), .B(n_782), .C(n_792), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AND2x4_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NOR3xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_805), .C(n_813), .Y(n_797) );
INVxp33_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OAI21xp33_ASAP7_75t_SL g805 ( .A1(n_806), .A2(n_809), .B(n_810), .Y(n_805) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_817), .B(n_820), .Y(n_813) );
INVxp67_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NOR2xp33_ASAP7_75t_SL g817 ( .A(n_818), .B(n_819), .Y(n_817) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_823), .Y(n_822) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
AND3x2_ASAP7_75t_L g858 ( .A(n_824), .B(n_834), .C(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_824), .B(n_880), .Y(n_879) );
INVx4_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AND2x6_ASAP7_75t_SL g828 ( .A(n_829), .B(n_831), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx3_ASAP7_75t_L g840 ( .A(n_830), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_830), .B(n_870), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_832), .B(n_834), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NOR2x1_ASAP7_75t_L g872 ( .A(n_833), .B(n_835), .Y(n_872) );
AND2x6_ASAP7_75t_SL g852 ( .A(n_834), .B(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
OAI21xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_842), .B(n_856), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_841), .Y(n_837) );
AOI21xp33_ASAP7_75t_L g856 ( .A1(n_838), .A2(n_857), .B(n_864), .Y(n_856) );
CKINVDCx11_ASAP7_75t_R g838 ( .A(n_839), .Y(n_838) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI31xp33_ASAP7_75t_SL g857 ( .A1(n_841), .A2(n_843), .A3(n_858), .B(n_860), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_849), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_845), .Y(n_848) );
BUFx3_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
BUFx12f_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx4_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx3_ASAP7_75t_L g863 ( .A(n_852), .Y(n_863) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_855), .Y(n_859) );
NOR2x1p5_ASAP7_75t_L g878 ( .A(n_859), .B(n_879), .Y(n_878) );
INVxp67_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_865), .Y(n_864) );
INVx3_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx6_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
BUFx10_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_874), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_875), .Y(n_874) );
CKINVDCx11_ASAP7_75t_R g875 ( .A(n_876), .Y(n_875) );
OR2x6_ASAP7_75t_L g876 ( .A(n_877), .B(n_882), .Y(n_876) );
OR2x6_ASAP7_75t_L g889 ( .A(n_877), .B(n_882), .Y(n_889) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .Y(n_883) );
INVxp33_ASAP7_75t_SL g885 ( .A(n_886), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_888), .Y(n_887) );
INVx4_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
endmodule