module fake_jpeg_5990_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_67;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx12_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_18),
.B1(n_16),
.B2(n_19),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_21),
.A2(n_22),
.B1(n_20),
.B2(n_17),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_13),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_10),
.Y(n_33)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_34),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_0),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_21),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_23),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_41),
.B1(n_29),
.B2(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_33),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_31),
.C(n_37),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_40),
.C(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_29),
.B1(n_47),
.B2(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_30),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_33),
.B1(n_47),
.B2(n_24),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_58),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

AOI31xp67_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_57),
.A3(n_50),
.B(n_62),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_68),
.A2(n_55),
.B(n_66),
.C(n_61),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_64),
.B1(n_53),
.B2(n_56),
.Y(n_71)
);

AOI321xp33_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_7),
.A3(n_9),
.B1(n_34),
.B2(n_69),
.C(n_55),
.Y(n_72)
);


endmodule