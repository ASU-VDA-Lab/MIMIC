module fake_jpeg_16256_n_92 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_92);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_92;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_3),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_4),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx2_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_7),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_0),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_23),
.A2(n_26),
.B(n_5),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_27),
.B(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_1),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_16),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_4),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_13),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_34),
.A2(n_41),
.B1(n_45),
.B2(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_33),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_23),
.A2(n_14),
.B1(n_22),
.B2(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_23),
.B(n_10),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_25),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_12),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_50),
.B(n_52),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_51),
.B1(n_5),
.B2(n_6),
.Y(n_57)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_12),
.C(n_17),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_54),
.C(n_58),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_12),
.C(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_64),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_6),
.C(n_7),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_7),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_65),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_8),
.C(n_11),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_46),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_67),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_34),
.B1(n_43),
.B2(n_44),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_43),
.B1(n_52),
.B2(n_44),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_70),
.B(n_37),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_60),
.B1(n_55),
.B2(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_56),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_72),
.A2(n_75),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_58),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_35),
.C(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_80),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_81),
.C(n_82),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_48),
.C(n_37),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_11),
.B(n_38),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_70),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_84),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_71),
.C(n_66),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_87),
.B1(n_86),
.B2(n_73),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_91),
.C(n_69),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_84),
.A3(n_85),
.B1(n_77),
.B2(n_67),
.C(n_69),
.Y(n_91)
);


endmodule