module fake_aes_5043_n_32 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AND2x4_ASAP7_75t_L g9 ( .A(n_7), .B(n_0), .Y(n_9) );
CKINVDCx20_ASAP7_75t_R g10 ( .A(n_0), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_1), .Y(n_11) );
AND2x2_ASAP7_75t_SL g12 ( .A(n_5), .B(n_8), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx2_ASAP7_75t_SL g15 ( .A(n_9), .Y(n_15) );
INVxp67_ASAP7_75t_SL g16 ( .A(n_9), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_13), .B(n_2), .Y(n_17) );
OAI21x1_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_14), .B(n_12), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_15), .B(n_11), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_19), .B(n_16), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_18), .B(n_15), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_18), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_22), .B(n_10), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
AOI21xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_23), .B(n_12), .Y(n_27) );
NOR2x1_ASAP7_75t_L g28 ( .A(n_26), .B(n_10), .Y(n_28) );
AND2x4_ASAP7_75t_L g29 ( .A(n_27), .B(n_2), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
AO22x2_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_28), .B1(n_3), .B2(n_6), .Y(n_31) );
INVxp67_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
endmodule