module real_jpeg_33610_n_23 (n_17, n_8, n_0, n_21, n_2, n_180, n_10, n_175, n_9, n_178, n_12, n_170, n_176, n_6, n_171, n_177, n_179, n_11, n_14, n_172, n_7, n_22, n_18, n_3, n_174, n_5, n_4, n_173, n_1, n_20, n_19, n_16, n_15, n_13, n_23);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_180;
input n_10;
input n_175;
input n_9;
input n_178;
input n_12;
input n_170;
input n_176;
input n_6;
input n_171;
input n_177;
input n_179;
input n_11;
input n_14;
input n_172;
input n_7;
input n_22;
input n_18;
input n_3;
input n_174;
input n_5;
input n_4;
input n_173;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_23;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_139;
wire n_33;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_150;
wire n_41;
wire n_74;
wire n_32;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AOI221xp5_ASAP7_75t_L g82 ( 
.A1(n_0),
.A2(n_15),
.B1(n_83),
.B2(n_89),
.C(n_90),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_0),
.B(n_83),
.C(n_89),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_1),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_2),
.B(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_2),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_4),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_4),
.Y(n_127)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_6),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_6),
.B(n_71),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_7),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_8),
.Y(n_61)
);

AOI322xp5_ASAP7_75t_L g123 ( 
.A1(n_8),
.A2(n_54),
.A3(n_56),
.B1(n_63),
.B2(n_124),
.C1(n_126),
.C2(n_180),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_9),
.B(n_65),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_10),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_11),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_14),
.Y(n_136)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_15),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_16),
.B(n_36),
.Y(n_156)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_17),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_17),
.B(n_116),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_18),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_18),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_22),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_31),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_129),
.B(n_151),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_42),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_41),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_39),
.B(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI31xp33_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_76),
.A3(n_114),
.B(n_119),
.Y(n_44)
);

NOR3xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_62),
.C(n_70),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_46),
.A2(n_120),
.B(n_123),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_54),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR3xp33_ASAP7_75t_L g124 ( 
.A(n_48),
.B(n_70),
.C(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_171),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_176),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

OA21x2_ASAP7_75t_SL g120 ( 
.A1(n_62),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_104),
.C(n_105),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_94),
.B(n_103),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_92),
.B2(n_93),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_102),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_137),
.C(n_141),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_155),
.C(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_136),
.Y(n_160)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_154),
.B(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI221xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_143),
.B1(n_152),
.B2(n_158),
.C(n_165),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.Y(n_142)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_170),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_172),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_173),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_174),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_175),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_177),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_178),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_179),
.Y(n_117)
);


endmodule