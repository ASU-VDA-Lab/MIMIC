module real_jpeg_17110_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_464),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_0),
.B(n_465),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_1),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_1),
.B(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_1),
.B(n_31),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g203 ( 
.A(n_1),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g334 ( 
.A(n_1),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_1),
.B(n_61),
.Y(n_385)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_2),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_2),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_3),
.B(n_83),
.Y(n_82)
);

NAND2xp67_ASAP7_75t_L g132 ( 
.A(n_3),
.B(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_3),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_3),
.B(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_3),
.B(n_436),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_4),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_4),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_4),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_5),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_6),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_6),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_6),
.B(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_6),
.B(n_137),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_6),
.B(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_SL g342 ( 
.A(n_6),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_6),
.B(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_7),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_7),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_7),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_7),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_7),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_7),
.B(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_7),
.Y(n_372)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_8),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_8),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_9),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_9),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_9),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_10),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_10),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_10),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_10),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_10),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_10),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_10),
.B(n_125),
.Y(n_298)
);

AND2x2_ASAP7_75t_SL g454 ( 
.A(n_10),
.B(n_455),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_11),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_11),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_11),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_11),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_12),
.Y(n_77)
);

NAND2x1_ASAP7_75t_L g96 ( 
.A(n_12),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_12),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_12),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_12),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_12),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_12),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_12),
.B(n_291),
.Y(n_290)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_13),
.Y(n_159)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_13),
.Y(n_242)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_14),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_14),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_14),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_14),
.B(n_129),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_14),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_14),
.B(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g336 ( 
.A(n_14),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_14),
.B(n_377),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_16),
.Y(n_116)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_17),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g293 ( 
.A(n_17),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_427),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_314),
.Y(n_21)
);

A2O1A1O1Ixp25_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_219),
.B(n_275),
.C(n_276),
.D(n_313),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_24),
.B(n_277),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_183),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_25),
.B(n_183),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_104),
.Y(n_25)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_26),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_68),
.C(n_92),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_28),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_42),
.C(n_54),
.Y(n_28)
);

XNOR2x1_ASAP7_75t_SL g243 ( 
.A(n_29),
.B(n_244),
.Y(n_243)
);

XNOR2x2_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_30),
.B(n_35),
.C(n_39),
.Y(n_94)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_32),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_38),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_39),
.B(n_161),
.Y(n_393)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_42),
.A2(n_43),
.B1(n_54),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_43),
.A2(n_44),
.B(n_49),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_46),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_47),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_48),
.B(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_52),
.Y(n_459)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_53),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_54),
.Y(n_245)
);

MAJx3_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.C(n_64),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_55),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_59),
.B(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_60),
.B(n_64),
.Y(n_191)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_63),
.Y(n_163)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_69),
.A2(n_92),
.B1(n_93),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_69),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_82),
.C(n_86),
.Y(n_69)
);

XNOR2x2_ASAP7_75t_SL g210 ( 
.A(n_70),
.B(n_211),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.C(n_78),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_71),
.B(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_74),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_74),
.A2(n_208),
.B1(n_228),
.B2(n_264),
.Y(n_438)
);

OR2x2_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_78),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_78),
.Y(n_227)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_81),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_82),
.B(n_86),
.Y(n_211)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_85),
.Y(n_209)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_101),
.C(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_96),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_98),
.Y(n_270)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_99),
.Y(n_235)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_102),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_155),
.B1(n_181),
.B2(n_182),
.Y(n_104)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_141),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_106),
.B(n_142),
.C(n_154),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_120),
.C(n_131),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_107),
.B(n_120),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_108),
.A2(n_113),
.B(n_117),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_119),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_112),
.A2(n_113),
.B1(n_194),
.B2(n_195),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_113),
.B(n_117),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_113),
.B(n_194),
.Y(n_193)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_117),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_119),
.B1(n_161),
.B2(n_164),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_117),
.B(n_157),
.C(n_164),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_117),
.B(n_385),
.Y(n_384)
);

BUFx12f_ASAP7_75t_L g358 ( 
.A(n_118),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_119),
.B(n_385),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.C(n_128),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_121),
.A2(n_122),
.B1(n_128),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_126),
.A2(n_213),
.B1(n_214),
.B2(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_126),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_126),
.A2(n_216),
.B1(n_300),
.B2(n_303),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_126),
.B(n_303),
.C(n_442),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_127),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_128),
.Y(n_215)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2x2_ASAP7_75t_L g217 ( 
.A(n_131),
.B(n_218),
.Y(n_217)
);

XNOR2x1_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_134),
.C(n_140),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_133)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_135),
.Y(n_437)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_140),
.B(n_458),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_154),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_153),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_148),
.B(n_152),
.C(n_153),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_148),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_148),
.B(n_290),
.C(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_155),
.B(n_181),
.C(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_156),
.B(n_166),
.C(n_169),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_161),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_161),
.A2(n_164),
.B1(n_208),
.B2(n_264),
.Y(n_305)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_163),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_SL g440 ( 
.A(n_164),
.B(n_208),
.C(n_306),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_168),
.A2(n_231),
.B1(n_412),
.B2(n_413),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_175),
.B1(n_179),
.B2(n_180),
.Y(n_170)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_175),
.B(n_180),
.C(n_227),
.Y(n_296)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_217),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_184),
.A2(n_185),
.B1(n_217),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_188),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_210),
.C(n_212),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_223),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_201),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_190),
.B(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_192),
.A2(n_193),
.B1(n_201),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.C(n_208),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_202),
.A2(n_208),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_202),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_203),
.B(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_207),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_208),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_217),
.Y(n_248)
);

AOI21x1_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_249),
.B(n_274),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_246),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_221),
.B(n_246),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.C(n_243),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_243),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.C(n_230),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_229),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.C(n_236),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_232),
.A2(n_236),
.B1(n_237),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_232),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_250),
.B(n_252),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.C(n_260),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_253),
.A2(n_254),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_256),
.A2(n_257),
.B1(n_260),
.B2(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_260),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.C(n_266),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_261),
.B(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_265),
.B(n_266),
.Y(n_417)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.C(n_273),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_267),
.A2(n_268),
.B1(n_273),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_271),
.B(n_405),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_273),
.Y(n_406)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_280),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_281),
.B(n_283),
.C(n_294),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_294),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_284),
.B(n_286),
.C(n_287),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_288),
.Y(n_450)
);

INVx3_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_304),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_296),
.B(n_304),
.C(n_446),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_297),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_298),
.Y(n_442)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_302),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND4xp25_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.C(n_317),
.D(n_318),
.Y(n_314)
);

OAI21x1_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_420),
.B(n_426),
.Y(n_318)
);

AOI21x1_ASAP7_75t_SL g319 ( 
.A1(n_320),
.A2(n_408),
.B(n_419),
.Y(n_319)
);

OAI21x1_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_387),
.B(n_407),
.Y(n_320)
);

AOI21x1_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_361),
.B(n_386),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_348),
.B(n_360),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_332),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_324),
.B(n_332),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_329),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_357),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_340),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_342),
.C(n_344),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_334),
.B(n_336),
.Y(n_382)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_344),
.B2(n_345),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_356),
.B(n_359),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_355),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_355),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_363),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_380),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_382),
.C(n_383),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_370),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_365),
.B(n_376),
.C(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_376),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_389),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_401),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_390),
.B(n_402),
.C(n_404),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_394),
.C(n_399),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_393),
.A2(n_394),
.B1(n_399),
.B2(n_400),
.Y(n_392)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_393),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_394),
.Y(n_400)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx8_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_418),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_SL g419 ( 
.A(n_409),
.B(n_418),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_416),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_415),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_415),
.C(n_416),
.Y(n_425)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_425),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_421),
.B(n_425),
.Y(n_426)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_462),
.Y(n_427)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_461),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_430),
.B(n_461),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_460),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_443),
.B2(n_444),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XNOR2x2_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_439),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_438),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_447),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_448),
.A2(n_449),
.B1(n_451),
.B2(n_452),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_454),
.B1(n_456),
.B2(n_457),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);


endmodule