module fake_netlist_1_12121_n_39 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_10), .B(n_0), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
INVx4_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_12), .B(n_2), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
INVxp67_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
OAI21x1_ASAP7_75t_SL g23 ( .A1(n_18), .A2(n_14), .B(n_15), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_22), .B(n_21), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
OAI33xp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_17), .A3(n_15), .B1(n_12), .B2(n_13), .B3(n_23), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
OAI21xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_18), .B(n_20), .Y(n_28) );
AOI221xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_21), .B1(n_18), .B2(n_16), .C(n_20), .Y(n_29) );
OAI211xp5_ASAP7_75t_SL g30 ( .A1(n_29), .A2(n_21), .B(n_3), .C(n_4), .Y(n_30) );
AOI211xp5_ASAP7_75t_SL g31 ( .A1(n_28), .A2(n_2), .B(n_3), .C(n_4), .Y(n_31) );
AOI22x1_ASAP7_75t_SL g32 ( .A1(n_29), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_32) );
AND4x1_ASAP7_75t_L g33 ( .A(n_31), .B(n_5), .C(n_6), .D(n_7), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_30), .A2(n_16), .B1(n_8), .B2(n_11), .Y(n_34) );
AND2x2_ASAP7_75t_L g35 ( .A(n_32), .B(n_16), .Y(n_35) );
HB1xp67_ASAP7_75t_L g36 ( .A(n_35), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_33), .Y(n_37) );
AO22x1_ASAP7_75t_L g38 ( .A1(n_36), .A2(n_32), .B1(n_34), .B2(n_37), .Y(n_38) );
INVx4_ASAP7_75t_L g39 ( .A(n_38), .Y(n_39) );
endmodule