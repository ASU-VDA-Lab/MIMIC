module fake_jpeg_9087_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_10),
.B(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_38),
.Y(n_72)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_25),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_8),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_35),
.Y(n_55)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_18),
.B1(n_30),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_53),
.B1(n_31),
.B2(n_22),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_62),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_18),
.B1(n_30),
.B2(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_55),
.B(n_63),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_44),
.B1(n_30),
.B2(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_58),
.A2(n_65),
.B1(n_17),
.B2(n_31),
.Y(n_100)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_47),
.B1(n_44),
.B2(n_38),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_30),
.B1(n_16),
.B2(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_74),
.Y(n_135)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_80),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_76),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_72),
.A2(n_40),
.B(n_31),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_103),
.B(n_21),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_78),
.A2(n_94),
.B1(n_111),
.B2(n_33),
.Y(n_128)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_38),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_87),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_84),
.B(n_91),
.Y(n_140)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_89),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_39),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_93),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_60),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_32),
.B1(n_46),
.B2(n_34),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_23),
.B(n_19),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_20),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_20),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_46),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_61),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_24),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_17),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_19),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_24),
.B1(n_22),
.B2(n_17),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_28),
.B1(n_25),
.B2(n_21),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g109 ( 
.A1(n_73),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_109),
.A2(n_22),
.B1(n_24),
.B2(n_19),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_120),
.B1(n_89),
.B2(n_112),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_117),
.B(n_127),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_119),
.B(n_103),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_41),
.B(n_33),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_124),
.A2(n_130),
.B(n_103),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_134),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_41),
.B(n_33),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_29),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_77),
.C(n_105),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_43),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_74),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_29),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_142),
.B(n_76),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_95),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_144),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_87),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_145),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_92),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_149),
.Y(n_188)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_111),
.B1(n_75),
.B2(n_85),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_163),
.B1(n_135),
.B2(n_141),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_130),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_156),
.C(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_154),
.A2(n_169),
.B(n_173),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_161),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_108),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_109),
.B1(n_86),
.B2(n_92),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_167),
.B(n_121),
.Y(n_197)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g162 ( 
.A(n_135),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_165),
.B1(n_133),
.B2(n_139),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_176),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_137),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_97),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_174),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_97),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_172),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_137),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_117),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_120),
.B1(n_140),
.B2(n_116),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_177),
.A2(n_192),
.B1(n_193),
.B2(n_204),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_163),
.A2(n_140),
.B1(n_120),
.B2(n_138),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_178),
.A2(n_206),
.B1(n_173),
.B2(n_164),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_123),
.B1(n_149),
.B2(n_159),
.Y(n_220)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_185),
.B(n_202),
.Y(n_235)
);

O2A1O1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_132),
.B(n_115),
.C(n_120),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_187),
.A2(n_197),
.B(n_209),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_115),
.B1(n_124),
.B2(n_119),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_139),
.B1(n_131),
.B2(n_133),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_175),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_195),
.A2(n_205),
.B1(n_208),
.B2(n_161),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_131),
.C(n_110),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_174),
.C(n_170),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_125),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_192),
.Y(n_218)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_148),
.A2(n_90),
.B1(n_106),
.B2(n_123),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_160),
.A2(n_90),
.B1(n_106),
.B2(n_98),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_153),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_125),
.B(n_117),
.Y(n_209)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_220),
.B1(n_230),
.B2(n_218),
.Y(n_242)
);

NOR2x1_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_152),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_219),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_223),
.Y(n_251)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_225),
.C(n_228),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_147),
.C(n_143),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_147),
.C(n_162),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_187),
.A2(n_88),
.B1(n_96),
.B2(n_81),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_230),
.A2(n_205),
.B1(n_208),
.B2(n_199),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_21),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_234),
.C(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_233),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_29),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_177),
.A2(n_191),
.B1(n_204),
.B2(n_197),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_236),
.A2(n_178),
.B1(n_191),
.B2(n_185),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_28),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_258),
.B1(n_220),
.B2(n_212),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_247),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_256),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_236),
.B1(n_215),
.B2(n_220),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_201),
.C(n_209),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_257),
.C(n_259),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_260),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_225),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_189),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_222),
.A2(n_180),
.B1(n_189),
.B2(n_203),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_212),
.B(n_198),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_263),
.Y(n_290)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_215),
.B1(n_220),
.B2(n_213),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_267),
.B1(n_271),
.B2(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_211),
.B(n_180),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_261),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_224),
.C(n_237),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_256),
.C(n_241),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_238),
.A2(n_203),
.B(n_186),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_10),
.B(n_15),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_2),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_96),
.B1(n_216),
.B2(n_28),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_279),
.B1(n_280),
.B2(n_1),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_259),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_266),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_25),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_257),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_253),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_243),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_274),
.Y(n_281)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_266),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_289),
.C(n_291),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_283),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_267),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_296),
.Y(n_304)
);

AO221x1_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_239),
.B1(n_250),
.B2(n_244),
.C(n_249),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_287),
.A2(n_295),
.B(n_283),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_288),
.B(n_292),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_241),
.C(n_252),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_10),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_264),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_268),
.B1(n_274),
.B2(n_269),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_285),
.B(n_276),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_307),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_278),
.C(n_272),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_306),
.C(n_308),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_286),
.B(n_294),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_9),
.C(n_14),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_286),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_313)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_281),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_313),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_316),
.B(n_317),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_293),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_282),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_300),
.A2(n_6),
.B(n_7),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_6),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_309),
.B1(n_302),
.B2(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_324),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_306),
.B(n_308),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_319),
.B(n_315),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_303),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_303),
.C(n_312),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_320),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_329),
.B(n_330),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_332),
.B(n_318),
.Y(n_334)
);

AOI321xp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_326),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_15),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_11),
.B(n_13),
.Y(n_337)
);


endmodule