module fake_netlist_6_3106_n_1751 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1751);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1751;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_65),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_62),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_61),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_44),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_91),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_30),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_42),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_94),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_27),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_129),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_74),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_27),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_40),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_88),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_21),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_60),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_114),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_157),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_29),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_87),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_52),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_69),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_100),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_95),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_51),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_63),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_4),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_93),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_89),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_109),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_84),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_119),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_96),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_139),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_143),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_50),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_108),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_18),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_16),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_136),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_36),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_64),
.Y(n_225)
);

BUFx2_ASAP7_75t_R g226 ( 
.A(n_172),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_5),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_39),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_24),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_141),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_72),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_16),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_59),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_86),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_111),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_162),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_150),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_121),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_97),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_40),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_106),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_145),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_137),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_23),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_104),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_0),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_12),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_82),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_71),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_152),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_120),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_3),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_22),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_155),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_13),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_90),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_66),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_133),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_134),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_19),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_47),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_70),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_116),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_53),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_127),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_12),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_103),
.Y(n_267)
);

HB1xp67_ASAP7_75t_SL g268 ( 
.A(n_13),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_124),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_30),
.Y(n_270)
);

BUFx8_ASAP7_75t_SL g271 ( 
.A(n_9),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_22),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_123),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_92),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_17),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_19),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_142),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_38),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_118),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_149),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_6),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_166),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_38),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_79),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_57),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_3),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_164),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_81),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_33),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_130),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_171),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_35),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_36),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_101),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_2),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_67),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_85),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_14),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_54),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_76),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_99),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_33),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_35),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_20),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_25),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_170),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_107),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_2),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_122),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_105),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_9),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_148),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_126),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_32),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_43),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_21),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_6),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_77),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_117),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_5),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_18),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_140),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_17),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_42),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_169),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_68),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_31),
.Y(n_327)
);

BUFx10_ASAP7_75t_L g328 ( 
.A(n_146),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_113),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_156),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_7),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_8),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_24),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_75),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_78),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_159),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_20),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_102),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_55),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_112),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_167),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_165),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_4),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_160),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_260),
.B(n_0),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_268),
.B(n_1),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_260),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_271),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_176),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_260),
.Y(n_350)
);

INVxp33_ASAP7_75t_SL g351 ( 
.A(n_272),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_260),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_260),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_260),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_224),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_173),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_229),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_260),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_260),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_343),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_179),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_244),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_219),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_219),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_343),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_312),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_343),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_178),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_343),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_343),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_184),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_252),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_189),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_316),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g377 ( 
.A(n_256),
.B(n_163),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_316),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_190),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_R g380 ( 
.A(n_200),
.B(n_161),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_194),
.B(n_1),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_253),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_235),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_233),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_191),
.B(n_7),
.Y(n_385)
);

INVxp33_ASAP7_75t_SL g386 ( 
.A(n_182),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_201),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_221),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_255),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_307),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_183),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_222),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_228),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_234),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_266),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_287),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_183),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_319),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_232),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_240),
.Y(n_400)
);

INVxp33_ASAP7_75t_L g401 ( 
.A(n_320),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_247),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_261),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_270),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_264),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_276),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_278),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_293),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_336),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_295),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_281),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_302),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_312),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_216),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_193),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_304),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_308),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_315),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_249),
.B(n_10),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_323),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_327),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_341),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_249),
.B(n_10),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_256),
.B(n_11),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_217),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_256),
.B(n_11),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_337),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_283),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_192),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_192),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_175),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_286),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_180),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_187),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_188),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_361),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_361),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_349),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_347),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_414),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_426),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_352),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_353),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_362),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_348),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_354),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_373),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_348),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_366),
.Y(n_453)
);

OA21x2_ASAP7_75t_L g454 ( 
.A1(n_345),
.A2(n_214),
.B(n_208),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_369),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_208),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_377),
.Y(n_457)
);

AND3x2_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_385),
.C(n_419),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_425),
.A2(n_215),
.B(n_214),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_377),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_377),
.Y(n_461)
);

AND2x2_ASAP7_75t_SL g462 ( 
.A(n_423),
.B(n_215),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_397),
.Y(n_463)
);

OA21x2_ASAP7_75t_L g464 ( 
.A1(n_431),
.A2(n_230),
.B(n_218),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_369),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_356),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_375),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_415),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_401),
.B(n_203),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_371),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_359),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_351),
.A2(n_209),
.B1(n_199),
.B2(n_188),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_355),
.B(n_209),
.C(n_199),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_360),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_R g475 ( 
.A(n_358),
.B(n_174),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g477 ( 
.A(n_415),
.B(n_218),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_372),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_372),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_437),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_377),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_431),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_384),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_409),
.B(n_195),
.Y(n_484)
);

NOR2xp67_ASAP7_75t_L g485 ( 
.A(n_432),
.B(n_198),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_432),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_367),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_367),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_367),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_363),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_367),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_374),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_374),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_382),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_387),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_388),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_413),
.B(n_203),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_436),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_396),
.B(n_213),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_390),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_435),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_392),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_382),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_428),
.B(n_230),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g505 ( 
.A1(n_393),
.A2(n_284),
.B(n_279),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_399),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

AND2x2_ASAP7_75t_SL g508 ( 
.A(n_381),
.B(n_279),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_402),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_L g510 ( 
.A(n_389),
.B(n_298),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_457),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_487),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_499),
.B(n_394),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_508),
.B(n_497),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_455),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_457),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_455),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_468),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_508),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_441),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_441),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_508),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_472),
.B(n_391),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_442),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_442),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_497),
.B(n_422),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_442),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_445),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_462),
.B(n_428),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_468),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_468),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_445),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_462),
.B(n_357),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_487),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_446),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_446),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_488),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_446),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_449),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_449),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_449),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_490),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_471),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_462),
.B(n_383),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_471),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_484),
.B(n_386),
.Y(n_548)
);

BUFx4f_ASAP7_75t_L g549 ( 
.A(n_457),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_457),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_456),
.B(n_398),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_471),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_488),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_457),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_440),
.Y(n_555)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_473),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_474),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_474),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_458),
.B(n_377),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_481),
.B(n_377),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_474),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_438),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_468),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_438),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_456),
.B(n_364),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_454),
.A2(n_377),
.B1(n_351),
.B2(n_368),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_439),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_439),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_457),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_489),
.B(n_395),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_450),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_466),
.B(n_395),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_463),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_450),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_453),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_469),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_480),
.B(n_386),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_456),
.B(n_365),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_453),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_510),
.B(n_404),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_454),
.A2(n_381),
.B1(n_391),
.B2(n_313),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_465),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_456),
.B(n_378),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_460),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_447),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_460),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_492),
.B(n_406),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_498),
.B(n_376),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_465),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_504),
.B(n_376),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_L g591 ( 
.A(n_460),
.B(n_380),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_470),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_460),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_470),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_476),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_493),
.B(n_407),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_460),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_475),
.A2(n_275),
.B1(n_303),
.B2(n_227),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_490),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_479),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_494),
.B(n_407),
.Y(n_601)
);

BUFx4f_ASAP7_75t_L g602 ( 
.A(n_460),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_461),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_479),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_489),
.B(n_411),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_503),
.B(n_411),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_467),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_467),
.B(n_430),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_495),
.B(n_430),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_476),
.Y(n_610)
);

HAxp5_ASAP7_75t_SL g611 ( 
.A(n_451),
.B(n_346),
.CON(n_611),
.SN(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_454),
.A2(n_313),
.B1(n_284),
.B2(n_416),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_478),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_461),
.B(n_434),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_478),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_498),
.B(n_434),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_454),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_505),
.A2(n_410),
.B1(n_421),
.B2(n_420),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_496),
.A2(n_207),
.B1(n_185),
.B2(n_311),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_479),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_491),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_461),
.B(n_205),
.Y(n_622)
);

NAND2x1p5_ASAP7_75t_L g623 ( 
.A(n_461),
.B(n_206),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_505),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_479),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_501),
.B(n_370),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_461),
.B(n_203),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_483),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_505),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_443),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_505),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_502),
.B(n_403),
.C(n_379),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_461),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_486),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_464),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_481),
.B(n_243),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_464),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_486),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_481),
.B(n_243),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_486),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_464),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_464),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_444),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_482),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_507),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_502),
.B(n_405),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_481),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_459),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_506),
.B(n_424),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_507),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_482),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_646),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_646),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_562),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_562),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_567),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_L g657 ( 
.A(n_637),
.B(n_193),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_565),
.B(n_506),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_519),
.B(n_477),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_519),
.B(n_477),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_577),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_523),
.A2(n_477),
.B1(n_459),
.B2(n_210),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_523),
.B(n_477),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_514),
.B(n_477),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_514),
.B(n_477),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_549),
.A2(n_485),
.B(n_507),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_548),
.B(n_448),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_567),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_530),
.B(n_477),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_560),
.B(n_511),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_564),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_556),
.B(n_580),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_560),
.B(n_193),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_534),
.A2(n_254),
.B1(n_265),
.B2(n_263),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_566),
.A2(n_477),
.B1(n_325),
.B2(n_297),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_574),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_564),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_590),
.B(n_452),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_574),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_568),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_560),
.B(n_193),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_549),
.A2(n_485),
.B(n_509),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_599),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_530),
.B(n_220),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_568),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_575),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_637),
.B(n_223),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_534),
.A2(n_246),
.B(n_509),
.C(n_418),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_575),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_637),
.B(n_237),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_637),
.B(n_241),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_579),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_579),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_637),
.B(n_248),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_571),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_571),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_R g697 ( 
.A(n_630),
.B(n_500),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_549),
.A2(n_285),
.B(n_282),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_576),
.B(n_573),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_588),
.B(n_346),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_582),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_582),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_590),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_595),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_546),
.B(n_267),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_635),
.A2(n_269),
.B(n_280),
.Y(n_706)
);

OAI221xp5_ASAP7_75t_L g707 ( 
.A1(n_581),
.A2(n_408),
.B1(n_412),
.B2(n_417),
.C(n_288),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_616),
.B(n_309),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_589),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_589),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_624),
.B(n_631),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_511),
.B(n_516),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_624),
.B(n_310),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_559),
.A2(n_291),
.B1(n_258),
.B2(n_257),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_511),
.B(n_193),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_612),
.A2(n_340),
.B1(n_344),
.B2(n_342),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_595),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_599),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_651),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_631),
.B(n_225),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_635),
.B(n_231),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_651),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_555),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_511),
.B(n_193),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_641),
.B(n_236),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_544),
.B(n_226),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_641),
.B(n_238),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_592),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_565),
.B(n_424),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_630),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_511),
.B(n_193),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_592),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_544),
.B(n_429),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_629),
.A2(n_429),
.B(n_339),
.C(n_333),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_551),
.A2(n_296),
.B1(n_294),
.B2(n_290),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_651),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_644),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_587),
.B(n_174),
.Y(n_738)
);

AND2x4_ASAP7_75t_SL g739 ( 
.A(n_607),
.B(n_243),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_551),
.A2(n_277),
.B1(n_274),
.B2(n_273),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_527),
.A2(n_328),
.B1(n_333),
.B2(n_332),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_609),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_642),
.B(n_239),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_644),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_642),
.B(n_242),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_642),
.B(n_245),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_527),
.B(n_250),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_594),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_614),
.A2(n_639),
.B1(n_636),
.B2(n_570),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_516),
.B(n_251),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_596),
.B(n_177),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_594),
.B(n_262),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_601),
.B(n_177),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_606),
.B(n_181),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_610),
.B(n_181),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_613),
.B(n_186),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_516),
.B(n_186),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_643),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_609),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_578),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_605),
.A2(n_344),
.B1(n_342),
.B2(n_196),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_629),
.A2(n_339),
.B(n_298),
.C(n_305),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_513),
.B(n_289),
.C(n_292),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_613),
.B(n_196),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_516),
.B(n_569),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_578),
.B(n_305),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_615),
.B(n_197),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_634),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_615),
.B(n_197),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_602),
.A2(n_338),
.B(n_335),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_512),
.B(n_202),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_634),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_638),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_572),
.B(n_334),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_638),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_600),
.B(n_334),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_600),
.B(n_204),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_604),
.B(n_204),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_583),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_622),
.A2(n_328),
.B1(n_317),
.B2(n_324),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_516),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_L g782 ( 
.A(n_569),
.B(n_211),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_604),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_L g784 ( 
.A(n_524),
.B(n_211),
.C(n_330),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_536),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_640),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_604),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_591),
.B(n_322),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_569),
.B(n_322),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_640),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_536),
.B(n_212),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_569),
.B(n_212),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_569),
.B(n_584),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_622),
.A2(n_331),
.B1(n_317),
.B2(n_321),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_602),
.A2(n_330),
.B(n_329),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_515),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_536),
.B(n_329),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_584),
.B(n_259),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_L g799 ( 
.A(n_626),
.B(n_300),
.C(n_326),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_627),
.A2(n_301),
.B1(n_326),
.B2(n_306),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_675),
.A2(n_749),
.B1(n_672),
.B2(n_705),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_711),
.B(n_617),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_661),
.B(n_598),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_664),
.A2(n_648),
.B(n_623),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_706),
.A2(n_647),
.B(n_597),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_667),
.B(n_598),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_760),
.B(n_539),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_738),
.B(n_628),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_737),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_737),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_671),
.B(n_518),
.Y(n_811)
);

AOI22x1_ASAP7_75t_SL g812 ( 
.A1(n_730),
.A2(n_758),
.B1(n_643),
.B2(n_585),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_793),
.A2(n_647),
.B(n_597),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_793),
.A2(n_647),
.B(n_554),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_751),
.B(n_608),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_670),
.A2(n_550),
.B(n_593),
.Y(n_816)
);

BUFx2_ASAP7_75t_SL g817 ( 
.A(n_723),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_670),
.A2(n_550),
.B(n_593),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_779),
.B(n_553),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_687),
.A2(n_550),
.B(n_593),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_690),
.A2(n_550),
.B(n_593),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_785),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_691),
.A2(n_554),
.B(n_597),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_744),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_699),
.B(n_584),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_694),
.A2(n_554),
.B(n_597),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_712),
.A2(n_554),
.B(n_603),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_703),
.B(n_619),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_708),
.B(n_553),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_734),
.A2(n_650),
.B(n_645),
.C(n_649),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_753),
.B(n_621),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_781),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_734),
.A2(n_650),
.B(n_645),
.C(n_618),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_765),
.A2(n_603),
.B(n_633),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_765),
.A2(n_586),
.B(n_584),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_697),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_759),
.A2(n_648),
.B1(n_633),
.B2(n_584),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_677),
.B(n_621),
.Y(n_838)
);

OR2x6_ASAP7_75t_SL g839 ( 
.A(n_730),
.B(n_758),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_669),
.A2(n_603),
.B(n_586),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_754),
.B(n_632),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_680),
.B(n_586),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_713),
.A2(n_633),
.B(n_586),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_743),
.A2(n_622),
.B(n_526),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_685),
.B(n_603),
.Y(n_845)
);

O2A1O1Ixp5_ASAP7_75t_L g846 ( 
.A1(n_750),
.A2(n_620),
.B(n_625),
.C(n_520),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_684),
.A2(n_623),
.B1(n_532),
.B2(n_518),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_652),
.B(n_623),
.Y(n_848)
);

AOI21x1_ASAP7_75t_L g849 ( 
.A1(n_745),
.A2(n_535),
.B(n_526),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_744),
.Y(n_850)
);

BUFx4f_ASAP7_75t_L g851 ( 
.A(n_683),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_659),
.A2(n_541),
.B(n_520),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_781),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_660),
.A2(n_541),
.B(n_521),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_658),
.A2(n_532),
.B1(n_531),
.B2(n_528),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_718),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_796),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_723),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_796),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_695),
.B(n_531),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_781),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_729),
.B(n_625),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_746),
.A2(n_620),
.B1(n_533),
.B2(n_535),
.Y(n_863)
);

NOR2xp67_ASAP7_75t_L g864 ( 
.A(n_678),
.B(n_515),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_654),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_654),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_696),
.B(n_558),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_701),
.B(n_558),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_742),
.B(n_318),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_774),
.A2(n_533),
.B(n_538),
.C(n_543),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_762),
.A2(n_538),
.B(n_543),
.C(n_547),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_663),
.A2(n_666),
.B(n_657),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_702),
.B(n_547),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_657),
.A2(n_537),
.B(n_521),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_655),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_762),
.A2(n_537),
.B(n_522),
.C(n_561),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_720),
.A2(n_540),
.B(n_522),
.Y(n_877)
);

AND2x4_ASAP7_75t_SL g878 ( 
.A(n_733),
.B(n_517),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_709),
.B(n_542),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_682),
.A2(n_542),
.B(n_525),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_710),
.B(n_545),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_728),
.B(n_540),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_656),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_662),
.A2(n_732),
.B1(n_748),
.B2(n_721),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_673),
.A2(n_557),
.B(n_552),
.Y(n_885)
);

AO21x1_ASAP7_75t_L g886 ( 
.A1(n_750),
.A2(n_681),
.B(n_673),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_653),
.B(n_306),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_747),
.B(n_557),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_700),
.B(n_517),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_697),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_688),
.B(n_529),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_725),
.A2(n_563),
.B(n_301),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_788),
.A2(n_563),
.B(n_154),
.Y(n_893)
);

NOR2xp67_ASAP7_75t_L g894 ( 
.A(n_799),
.B(n_153),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_729),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_656),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_727),
.A2(n_611),
.B1(n_131),
.B2(n_128),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_726),
.B(n_14),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_783),
.A2(n_125),
.B(n_115),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_729),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_688),
.B(n_15),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_715),
.A2(n_83),
.B(n_80),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_787),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_668),
.B(n_58),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_766),
.B(n_15),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_776),
.A2(n_25),
.B(n_26),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_791),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_739),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_763),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_714),
.B(n_26),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_668),
.B(n_28),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_777),
.A2(n_28),
.B(n_31),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_676),
.B(n_32),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_784),
.B(n_34),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_739),
.B(n_34),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_676),
.B(n_37),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_778),
.A2(n_37),
.B(n_39),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_679),
.B(n_41),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_761),
.B(n_41),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_679),
.B(n_43),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_752),
.A2(n_44),
.B(n_45),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_719),
.A2(n_46),
.B(n_47),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_797),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_686),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_686),
.B(n_46),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_689),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_692),
.B(n_48),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_674),
.B(n_740),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_692),
.B(n_48),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_782),
.A2(n_49),
.B(n_50),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_693),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_693),
.B(n_49),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_707),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_704),
.B(n_717),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_715),
.A2(n_56),
.B(n_724),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_704),
.B(n_717),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_771),
.A2(n_735),
.B1(n_789),
.B2(n_757),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_719),
.A2(n_736),
.B(n_722),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_757),
.A2(n_792),
.B1(n_789),
.B2(n_798),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_722),
.B(n_736),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_768),
.B(n_772),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_724),
.A2(n_792),
.B(n_798),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_768),
.B(n_772),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_731),
.A2(n_773),
.B(n_790),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_731),
.A2(n_773),
.B(n_790),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_775),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_755),
.B(n_767),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_775),
.B(n_786),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_756),
.B(n_769),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_764),
.A2(n_698),
.B(n_795),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_L g951 ( 
.A(n_716),
.B(n_800),
.C(n_770),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_780),
.A2(n_741),
.B(n_794),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_706),
.A2(n_602),
.B(n_549),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_706),
.A2(n_602),
.B(n_549),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_734),
.A2(n_762),
.B(n_688),
.C(n_519),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_661),
.B(n_672),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_654),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_661),
.B(n_672),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_706),
.A2(n_602),
.B(n_549),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_672),
.A2(n_523),
.B(n_519),
.C(n_514),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_781),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_711),
.A2(n_665),
.B(n_664),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_734),
.A2(n_762),
.B(n_688),
.C(n_519),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_711),
.A2(n_665),
.B(n_664),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_928),
.A2(n_806),
.B1(n_841),
.B2(n_831),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_866),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_956),
.B(n_958),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_836),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_889),
.Y(n_969)
);

AOI221xp5_ASAP7_75t_SL g970 ( 
.A1(n_952),
.A2(n_963),
.B1(n_955),
.B2(n_933),
.C(n_922),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_900),
.B(n_895),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_947),
.B(n_907),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_803),
.B(n_808),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_895),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_852),
.A2(n_854),
.B(n_874),
.Y(n_975)
);

CKINVDCx11_ASAP7_75t_R g976 ( 
.A(n_839),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_962),
.A2(n_964),
.B(n_960),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_802),
.A2(n_801),
.B(n_833),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_805),
.A2(n_954),
.B(n_953),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_856),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_851),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_840),
.A2(n_938),
.B(n_821),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_959),
.A2(n_814),
.B(n_813),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_851),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_817),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_923),
.B(n_878),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_900),
.B(n_819),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_822),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_802),
.A2(n_804),
.B(n_884),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_890),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_949),
.B(n_807),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_820),
.A2(n_826),
.B(n_823),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_950),
.A2(n_818),
.B(n_816),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_875),
.Y(n_994)
);

NAND2x1p5_ASAP7_75t_L g995 ( 
.A(n_822),
.B(n_832),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_858),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_819),
.B(n_807),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_924),
.Y(n_998)
);

OAI22x1_ASAP7_75t_L g999 ( 
.A1(n_919),
.A2(n_914),
.B1(n_898),
.B2(n_909),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_822),
.Y(n_1000)
);

OR2x6_ASAP7_75t_L g1001 ( 
.A(n_929),
.B(n_862),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_812),
.Y(n_1002)
);

O2A1O1Ixp5_ASAP7_75t_L g1003 ( 
.A1(n_892),
.A2(n_937),
.B(n_939),
.C(n_849),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_844),
.A2(n_942),
.B(n_863),
.Y(n_1004)
);

OAI22x1_ASAP7_75t_L g1005 ( 
.A1(n_915),
.A2(n_908),
.B1(n_869),
.B2(n_887),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_888),
.A2(n_843),
.B(n_829),
.Y(n_1006)
);

OR2x6_ASAP7_75t_L g1007 ( 
.A(n_929),
.B(n_862),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_883),
.Y(n_1008)
);

OR2x6_ASAP7_75t_L g1009 ( 
.A(n_910),
.B(n_864),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_905),
.A2(n_871),
.B(n_899),
.C(n_830),
.Y(n_1010)
);

O2A1O1Ixp5_ASAP7_75t_L g1011 ( 
.A1(n_886),
.A2(n_825),
.B(n_870),
.C(n_848),
.Y(n_1011)
);

AO31x2_ASAP7_75t_L g1012 ( 
.A1(n_837),
.A2(n_913),
.A3(n_927),
.B(n_925),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_876),
.A2(n_846),
.B(n_885),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_903),
.B(n_897),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_827),
.A2(n_835),
.B(n_834),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_838),
.B(n_881),
.Y(n_1016)
);

AOI21x1_ASAP7_75t_L g1017 ( 
.A1(n_904),
.A2(n_891),
.B(n_934),
.Y(n_1017)
);

NAND3xp33_ASAP7_75t_L g1018 ( 
.A(n_901),
.B(n_921),
.C(n_930),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_924),
.Y(n_1019)
);

AO31x2_ASAP7_75t_L g1020 ( 
.A1(n_911),
.A2(n_913),
.A3(n_932),
.B(n_916),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_944),
.A2(n_945),
.B(n_940),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_935),
.B(n_917),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_936),
.A2(n_941),
.B(n_948),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_853),
.B(n_861),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_853),
.B(n_961),
.Y(n_1025)
);

NAND2x1p5_ASAP7_75t_L g1026 ( 
.A(n_832),
.B(n_961),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_842),
.A2(n_845),
.B(n_948),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_911),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_943),
.A2(n_881),
.B(n_904),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_811),
.A2(n_867),
.B(n_868),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_847),
.A2(n_912),
.B(n_906),
.C(n_855),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_811),
.A2(n_916),
.B(n_918),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_918),
.A2(n_920),
.B(n_882),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_SL g1034 ( 
.A1(n_873),
.A2(n_860),
.B(n_879),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_931),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_861),
.A2(n_957),
.B1(n_926),
.B2(n_896),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_865),
.B(n_809),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_810),
.B(n_824),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_893),
.A2(n_850),
.B(n_857),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_859),
.B(n_946),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_894),
.B(n_902),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_841),
.B(n_831),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_962),
.A2(n_964),
.B(n_960),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_851),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_956),
.B(n_700),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_805),
.A2(n_602),
.B(n_549),
.Y(n_1046)
);

AOI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_806),
.A2(n_841),
.B(n_815),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_841),
.B(n_831),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_SL g1049 ( 
.A1(n_886),
.A2(n_922),
.B(n_955),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_851),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_822),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_841),
.B(n_831),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_956),
.B(n_700),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_SL g1054 ( 
.A1(n_901),
.A2(n_559),
.B(n_911),
.Y(n_1054)
);

OAI22x1_ASAP7_75t_L g1055 ( 
.A1(n_806),
.A2(n_619),
.B1(n_815),
.B2(n_598),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_962),
.A2(n_964),
.B(n_960),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_924),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_960),
.A2(n_884),
.A3(n_870),
.B(n_939),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_895),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_956),
.B(n_700),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_828),
.B(n_700),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_841),
.A2(n_806),
.B(n_815),
.C(n_928),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_805),
.A2(n_602),
.B(n_549),
.Y(n_1063)
);

OAI21xp33_ASAP7_75t_L g1064 ( 
.A1(n_841),
.A2(n_806),
.B(n_815),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_SL g1065 ( 
.A1(n_806),
.A2(n_841),
.B(n_952),
.Y(n_1065)
);

AOI21xp33_ASAP7_75t_L g1066 ( 
.A1(n_806),
.A2(n_841),
.B(n_815),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_828),
.B(n_700),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_841),
.B(n_831),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_962),
.A2(n_964),
.B(n_960),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_SL g1070 ( 
.A1(n_886),
.A2(n_922),
.B(n_955),
.Y(n_1070)
);

NOR2xp67_ASAP7_75t_SL g1071 ( 
.A(n_895),
.B(n_817),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_962),
.A2(n_964),
.B(n_960),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_924),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_866),
.Y(n_1074)
);

AOI221x1_ASAP7_75t_L g1075 ( 
.A1(n_951),
.A2(n_939),
.B1(n_937),
.B2(n_960),
.C(n_801),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_895),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_828),
.B(n_700),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_877),
.A2(n_872),
.B(n_880),
.Y(n_1078)
);

AO21x2_ASAP7_75t_L g1079 ( 
.A1(n_953),
.A2(n_959),
.B(n_954),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_841),
.B(n_831),
.Y(n_1080)
);

AOI21xp33_ASAP7_75t_L g1081 ( 
.A1(n_806),
.A2(n_841),
.B(n_815),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_851),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_895),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_828),
.B(n_700),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_841),
.B(n_831),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_962),
.A2(n_964),
.B(n_960),
.Y(n_1086)
);

NAND2x1p5_ASAP7_75t_L g1087 ( 
.A(n_900),
.B(n_822),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_962),
.A2(n_964),
.B(n_960),
.Y(n_1088)
);

BUFx4_ASAP7_75t_SL g1089 ( 
.A(n_858),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_956),
.B(n_700),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_924),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_924),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_815),
.B(n_672),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_841),
.B(n_831),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_806),
.A2(n_841),
.B1(n_815),
.B2(n_928),
.Y(n_1095)
);

CKINVDCx8_ASAP7_75t_R g1096 ( 
.A(n_817),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_965),
.B(n_1042),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_997),
.B(n_987),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_973),
.B(n_1045),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_SL g1100 ( 
.A1(n_1048),
.A2(n_1068),
.B1(n_1094),
.B2(n_1085),
.Y(n_1100)
);

INVx6_ASAP7_75t_L g1101 ( 
.A(n_1059),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_980),
.Y(n_1102)
);

AO21x1_ASAP7_75t_L g1103 ( 
.A1(n_1065),
.A2(n_1066),
.B(n_1047),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_969),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_1089),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_996),
.Y(n_1106)
);

OAI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1095),
.A2(n_1080),
.B1(n_1052),
.B2(n_1081),
.Y(n_1107)
);

INVx6_ASAP7_75t_L g1108 ( 
.A(n_1059),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1064),
.B(n_1062),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1037),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_988),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_1082),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1053),
.B(n_1060),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_966),
.Y(n_1114)
);

OA22x2_ASAP7_75t_L g1115 ( 
.A1(n_1055),
.A2(n_1065),
.B1(n_999),
.B2(n_967),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_985),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1093),
.B(n_1028),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_981),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_994),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_969),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_997),
.B(n_987),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1008),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_983),
.A2(n_979),
.B(n_993),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1090),
.B(n_1061),
.Y(n_1124)
);

BUFx12f_ASAP7_75t_L g1125 ( 
.A(n_976),
.Y(n_1125)
);

OAI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_972),
.A2(n_1084),
.B1(n_1077),
.B2(n_1067),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1001),
.B(n_1007),
.Y(n_1127)
);

NAND2x1_ASAP7_75t_L g1128 ( 
.A(n_1000),
.B(n_1001),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_968),
.Y(n_1129)
);

AOI21xp33_ASAP7_75t_SL g1130 ( 
.A1(n_1005),
.A2(n_986),
.B(n_984),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1016),
.B(n_1023),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_991),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_988),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_992),
.A2(n_978),
.B(n_1006),
.Y(n_1134)
);

OA21x2_ASAP7_75t_L g1135 ( 
.A1(n_1075),
.A2(n_970),
.B(n_989),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1074),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1079),
.A2(n_1046),
.B(n_1063),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1044),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1049),
.A2(n_1070),
.B1(n_1018),
.B2(n_1014),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1038),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1096),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1001),
.B(n_1007),
.Y(n_1142)
);

AO21x2_ASAP7_75t_L g1143 ( 
.A1(n_989),
.A2(n_1056),
.B(n_1088),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1050),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1040),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_998),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_1007),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_988),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1009),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1010),
.A2(n_970),
.B(n_1018),
.C(n_1031),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1009),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1019),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1059),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1023),
.B(n_1030),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1035),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1057),
.Y(n_1156)
);

O2A1O1Ixp5_ASAP7_75t_L g1157 ( 
.A1(n_1004),
.A2(n_1015),
.B(n_1011),
.C(n_1056),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_990),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1073),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_977),
.A2(n_1072),
.B(n_1069),
.C(n_1043),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1091),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1002),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1051),
.B(n_1076),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_971),
.B(n_974),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_974),
.B(n_1076),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1092),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1083),
.B(n_1000),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1083),
.B(n_1024),
.Y(n_1168)
);

NOR2xp67_ASAP7_75t_L g1169 ( 
.A(n_971),
.B(n_1025),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1032),
.B(n_1033),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_977),
.A2(n_1043),
.B1(n_1088),
.B2(n_1069),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1024),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1025),
.B(n_1071),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1022),
.B(n_1041),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1032),
.B(n_1033),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1087),
.B(n_1020),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_995),
.A2(n_1086),
.B1(n_1034),
.B2(n_1026),
.Y(n_1177)
);

CKINVDCx16_ASAP7_75t_R g1178 ( 
.A(n_1022),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1026),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1041),
.B(n_1029),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1086),
.A2(n_1021),
.B(n_1078),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1022),
.B(n_1036),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_982),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1021),
.A2(n_1027),
.B1(n_1013),
.B2(n_1039),
.Y(n_1184)
);

AOI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1017),
.A2(n_1013),
.B(n_975),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1020),
.B(n_1058),
.Y(n_1186)
);

OAI221xp5_ASAP7_75t_L g1187 ( 
.A1(n_1054),
.A2(n_1095),
.B1(n_1064),
.B2(n_1081),
.C(n_1066),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1012),
.A2(n_1095),
.B1(n_1062),
.B2(n_965),
.Y(n_1188)
);

BUFx10_ASAP7_75t_L g1189 ( 
.A(n_1058),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1012),
.A2(n_983),
.B(n_979),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_980),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_983),
.A2(n_979),
.B(n_805),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1095),
.A2(n_1062),
.B1(n_965),
.B2(n_1048),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1095),
.A2(n_1062),
.B1(n_965),
.B2(n_1048),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1061),
.B(n_1067),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_997),
.B(n_987),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_965),
.A2(n_1095),
.B1(n_806),
.B2(n_1064),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1047),
.A2(n_1066),
.B1(n_1081),
.B2(n_1064),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_965),
.B(n_1042),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1095),
.A2(n_1062),
.B1(n_965),
.B2(n_1048),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_973),
.B(n_1045),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_965),
.B(n_1042),
.Y(n_1202)
);

INVx6_ASAP7_75t_L g1203 ( 
.A(n_1059),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_988),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1037),
.Y(n_1205)
);

INVx3_ASAP7_75t_SL g1206 ( 
.A(n_985),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1037),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_973),
.B(n_1045),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_973),
.B(n_1045),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_983),
.A2(n_979),
.B(n_805),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_988),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_973),
.B(n_1045),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_983),
.A2(n_979),
.B(n_805),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_983),
.A2(n_979),
.B(n_805),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1061),
.B(n_1067),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1047),
.A2(n_1066),
.B1(n_1081),
.B2(n_1064),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1075),
.A2(n_1003),
.B(n_978),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1061),
.B(n_1067),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_973),
.B(n_1045),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_969),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1061),
.B(n_1067),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_966),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_973),
.B(n_1045),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_965),
.B(n_1042),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1037),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_996),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_983),
.A2(n_979),
.B(n_805),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_980),
.Y(n_1228)
);

AOI222xp33_ASAP7_75t_L g1229 ( 
.A1(n_1064),
.A2(n_1055),
.B1(n_806),
.B2(n_965),
.C1(n_1062),
.C2(n_973),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_997),
.B(n_987),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_965),
.B(n_1042),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1095),
.A2(n_1062),
.B1(n_965),
.B2(n_1048),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_980),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_965),
.B(n_1042),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1047),
.A2(n_1066),
.B1(n_1081),
.B2(n_1064),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1197),
.A2(n_1235),
.B1(n_1216),
.B2(n_1198),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1206),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1153),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1206),
.Y(n_1239)
);

OR2x6_ASAP7_75t_L g1240 ( 
.A(n_1174),
.B(n_1177),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1193),
.A2(n_1232),
.B1(n_1200),
.B2(n_1194),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1122),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1119),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1097),
.A2(n_1224),
.B1(n_1234),
.B2(n_1202),
.Y(n_1244)
);

AOI222xp33_ASAP7_75t_L g1245 ( 
.A1(n_1107),
.A2(n_1109),
.B1(n_1219),
.B2(n_1099),
.C1(n_1212),
.C2(n_1223),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1136),
.Y(n_1246)
);

AOI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1181),
.A2(n_1134),
.B(n_1190),
.Y(n_1247)
);

INVx6_ASAP7_75t_L g1248 ( 
.A(n_1164),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1201),
.B(n_1208),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1105),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1120),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1209),
.B(n_1107),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1102),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1097),
.A2(n_1234),
.B1(n_1202),
.B2(n_1231),
.Y(n_1254)
);

CKINVDCx11_ASAP7_75t_R g1255 ( 
.A(n_1125),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1222),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1127),
.B(n_1142),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1110),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1199),
.A2(n_1231),
.B1(n_1224),
.B2(n_1100),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1180),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1169),
.B(n_1164),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_SL g1262 ( 
.A1(n_1100),
.A2(n_1109),
.B1(n_1124),
.B2(n_1199),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1188),
.B(n_1170),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1229),
.B(n_1103),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1106),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1187),
.A2(n_1150),
.B(n_1182),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1205),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1115),
.B(n_1132),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1117),
.A2(n_1126),
.B1(n_1104),
.B2(n_1132),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1115),
.B(n_1186),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1140),
.B(n_1145),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1113),
.B(n_1126),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1180),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1187),
.A2(n_1221),
.B1(n_1195),
.B2(n_1218),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1207),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1225),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1226),
.Y(n_1277)
);

INVx8_ASAP7_75t_L g1278 ( 
.A(n_1098),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1120),
.B(n_1220),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1152),
.Y(n_1280)
);

INVx6_ASAP7_75t_L g1281 ( 
.A(n_1098),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1156),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1220),
.B(n_1176),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1143),
.B(n_1171),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1166),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1146),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1155),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1159),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1172),
.B(n_1147),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_1158),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1189),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1161),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1129),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1215),
.A2(n_1171),
.B1(n_1143),
.B2(n_1151),
.Y(n_1294)
);

BUFx10_ASAP7_75t_L g1295 ( 
.A(n_1168),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1112),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1104),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1189),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1116),
.B(n_1131),
.Y(n_1299)
);

AO21x1_ASAP7_75t_L g1300 ( 
.A1(n_1160),
.A2(n_1134),
.B(n_1154),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1131),
.B(n_1230),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1178),
.A2(n_1191),
.B1(n_1139),
.B2(n_1118),
.Y(n_1302)
);

INVx5_ASAP7_75t_L g1303 ( 
.A(n_1183),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1228),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1192),
.A2(n_1214),
.B(n_1213),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1157),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1183),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1147),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1135),
.B(n_1139),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1233),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1135),
.B(n_1175),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1141),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1170),
.B(n_1175),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1217),
.B(n_1163),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1121),
.B(n_1230),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1149),
.A2(n_1196),
.B1(n_1121),
.B2(n_1191),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_SL g1317 ( 
.A1(n_1138),
.A2(n_1196),
.B1(n_1173),
.B2(n_1154),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1144),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1165),
.B(n_1130),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1184),
.A2(n_1128),
.B1(n_1167),
.B2(n_1179),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1111),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1153),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1153),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1111),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1111),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1148),
.B(n_1204),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1184),
.A2(n_1101),
.B1(n_1108),
.B2(n_1203),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1181),
.B(n_1123),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1133),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1210),
.A2(n_1227),
.B(n_1214),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1101),
.A2(n_1108),
.B1(n_1203),
.B2(n_1148),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1211),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1101),
.A2(n_1108),
.B1(n_1203),
.B2(n_1204),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1211),
.B(n_1162),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1185),
.A2(n_992),
.B(n_1137),
.Y(n_1335)
);

BUFx4f_ASAP7_75t_SL g1336 ( 
.A(n_1158),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1109),
.B(n_1197),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1114),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1193),
.A2(n_1047),
.B1(n_1081),
.B2(n_1066),
.Y(n_1339)
);

NAND2x1p5_ASAP7_75t_L g1340 ( 
.A(n_1179),
.B(n_1071),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1193),
.A2(n_1047),
.B1(n_1081),
.B2(n_1066),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1105),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1153),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1153),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1197),
.A2(n_1095),
.B1(n_806),
.B2(n_965),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1109),
.B(n_1197),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1125),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1099),
.B(n_973),
.Y(n_1348)
);

AOI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1247),
.A2(n_1330),
.B(n_1305),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1251),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1251),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1279),
.Y(n_1352)
);

AO21x2_ASAP7_75t_L g1353 ( 
.A1(n_1335),
.A2(n_1300),
.B(n_1306),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1270),
.B(n_1283),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1311),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1303),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1311),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1284),
.Y(n_1358)
);

OR2x6_ASAP7_75t_L g1359 ( 
.A(n_1240),
.B(n_1328),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1266),
.A2(n_1254),
.B(n_1244),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1263),
.B(n_1272),
.Y(n_1361)
);

NAND2x1_ASAP7_75t_L g1362 ( 
.A(n_1240),
.B(n_1260),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1309),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1309),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1313),
.B(n_1337),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1263),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1345),
.A2(n_1236),
.B(n_1259),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1313),
.B(n_1337),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1314),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1339),
.A2(n_1341),
.B(n_1241),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1314),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1346),
.B(n_1264),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1346),
.B(n_1264),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1246),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1237),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1256),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1298),
.A2(n_1268),
.B(n_1294),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1256),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1237),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1268),
.A2(n_1252),
.B(n_1307),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1308),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1269),
.B(n_1274),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1240),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1253),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1295),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1295),
.Y(n_1386)
);

NOR2x1_ASAP7_75t_SL g1387 ( 
.A(n_1320),
.B(n_1307),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1249),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1243),
.Y(n_1389)
);

BUFx12f_ASAP7_75t_L g1390 ( 
.A(n_1255),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1291),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1273),
.B(n_1291),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1291),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1301),
.A2(n_1285),
.B(n_1280),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1257),
.B(n_1271),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1257),
.B(n_1245),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1282),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1242),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1293),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1338),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1286),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1299),
.B(n_1348),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1319),
.A2(n_1292),
.B(n_1288),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1295),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1302),
.A2(n_1317),
.B(n_1327),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1287),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1258),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1262),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1257),
.B(n_1289),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1267),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1318),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1275),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1276),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1297),
.B(n_1289),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1332),
.B(n_1310),
.Y(n_1415)
);

CKINVDCx6p67_ASAP7_75t_R g1416 ( 
.A(n_1293),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1359),
.B(n_1261),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1363),
.B(n_1329),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1383),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1364),
.B(n_1304),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1370),
.A2(n_1281),
.B1(n_1316),
.B2(n_1310),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1380),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1359),
.B(n_1261),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1364),
.B(n_1239),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1359),
.B(n_1261),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1358),
.B(n_1323),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1403),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1366),
.B(n_1324),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1358),
.B(n_1325),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1359),
.B(n_1322),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1389),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1380),
.Y(n_1432)
);

OR2x2_ASAP7_75t_SL g1433 ( 
.A(n_1382),
.B(n_1334),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1408),
.A2(n_1281),
.B1(n_1312),
.B2(n_1278),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1383),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_1403),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1369),
.B(n_1238),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1361),
.B(n_1340),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1380),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1371),
.B(n_1238),
.Y(n_1440)
);

AOI21xp33_ASAP7_75t_L g1441 ( 
.A1(n_1360),
.A2(n_1315),
.B(n_1340),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1355),
.B(n_1334),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1359),
.B(n_1343),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1380),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1408),
.A2(n_1281),
.B1(n_1312),
.B2(n_1278),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1372),
.B(n_1238),
.Y(n_1446)
);

AOI322xp5_ASAP7_75t_L g1447 ( 
.A1(n_1373),
.A2(n_1290),
.A3(n_1333),
.B1(n_1296),
.B2(n_1265),
.C1(n_1277),
.C2(n_1342),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1357),
.B(n_1344),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1357),
.B(n_1344),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1354),
.B(n_1344),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1392),
.B(n_1277),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1403),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1352),
.B(n_1296),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1365),
.B(n_1326),
.Y(n_1454)
);

OAI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1382),
.A2(n_1248),
.B1(n_1336),
.B2(n_1278),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1403),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1353),
.B(n_1248),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1368),
.B(n_1248),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1447),
.A2(n_1405),
.B(n_1396),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1448),
.B(n_1377),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1421),
.A2(n_1367),
.B1(n_1416),
.B2(n_1388),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1438),
.B(n_1384),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1449),
.B(n_1368),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1441),
.B(n_1367),
.C(n_1411),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1449),
.B(n_1395),
.Y(n_1465)
);

NOR3xp33_ASAP7_75t_L g1466 ( 
.A(n_1441),
.B(n_1402),
.C(n_1362),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1438),
.B(n_1360),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1450),
.B(n_1395),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1454),
.B(n_1360),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1455),
.B(n_1409),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_L g1471 ( 
.A(n_1447),
.B(n_1394),
.C(n_1391),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1434),
.A2(n_1362),
.B(n_1396),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1431),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1424),
.B(n_1394),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1417),
.B(n_1409),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1427),
.A2(n_1452),
.B(n_1436),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1420),
.B(n_1394),
.Y(n_1477)
);

OAI221xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1445),
.A2(n_1416),
.B1(n_1414),
.B2(n_1379),
.C(n_1375),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1417),
.B(n_1409),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1420),
.B(n_1394),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1430),
.A2(n_1423),
.B1(n_1417),
.B2(n_1425),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1442),
.B(n_1350),
.Y(n_1482)
);

NOR3xp33_ASAP7_75t_L g1483 ( 
.A(n_1428),
.B(n_1349),
.C(n_1331),
.Y(n_1483)
);

OAI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1453),
.A2(n_1375),
.B1(n_1379),
.B2(n_1386),
.C(n_1385),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1418),
.B(n_1428),
.Y(n_1485)
);

NOR3xp33_ASAP7_75t_L g1486 ( 
.A(n_1458),
.B(n_1349),
.C(n_1255),
.Y(n_1486)
);

OAI21xp33_ASAP7_75t_L g1487 ( 
.A1(n_1422),
.A2(n_1414),
.B(n_1398),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1430),
.A2(n_1407),
.B(n_1413),
.Y(n_1488)
);

AND2x2_ASAP7_75t_SL g1489 ( 
.A(n_1417),
.B(n_1409),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_1432),
.B(n_1393),
.C(n_1397),
.Y(n_1490)
);

AND2x2_ASAP7_75t_SL g1491 ( 
.A(n_1423),
.B(n_1356),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1437),
.B(n_1440),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_L g1493 ( 
.A(n_1432),
.B(n_1393),
.C(n_1376),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1439),
.B(n_1393),
.C(n_1376),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1426),
.B(n_1351),
.Y(n_1495)
);

OAI31xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1423),
.A2(n_1415),
.A3(n_1400),
.B(n_1387),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1439),
.B(n_1378),
.C(n_1374),
.Y(n_1497)
);

OAI221xp5_ASAP7_75t_L g1498 ( 
.A1(n_1453),
.A2(n_1379),
.B1(n_1375),
.B2(n_1386),
.C(n_1385),
.Y(n_1498)
);

AOI221x1_ASAP7_75t_SL g1499 ( 
.A1(n_1446),
.A2(n_1406),
.B1(n_1401),
.B2(n_1410),
.C(n_1412),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1429),
.B(n_1381),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1476),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1473),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1473),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1491),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1476),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1469),
.B(n_1444),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1476),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1476),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1460),
.B(n_1456),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1467),
.B(n_1419),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1474),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1477),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1480),
.B(n_1427),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1497),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1475),
.B(n_1423),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1475),
.B(n_1425),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1499),
.B(n_1452),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1492),
.B(n_1457),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1490),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1493),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1494),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1489),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1485),
.B(n_1466),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1462),
.B(n_1399),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1500),
.B(n_1435),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1487),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1463),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1487),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1482),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1502),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1502),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1503),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1522),
.B(n_1491),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1522),
.B(n_1489),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1503),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1515),
.B(n_1479),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1504),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1504),
.B(n_1489),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1525),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1523),
.B(n_1465),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1504),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1510),
.B(n_1495),
.Y(n_1542)
);

INVxp33_ASAP7_75t_L g1543 ( 
.A(n_1523),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1504),
.B(n_1464),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1501),
.Y(n_1545)
);

NAND3xp33_ASAP7_75t_L g1546 ( 
.A(n_1514),
.B(n_1486),
.C(n_1459),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1517),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1525),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1529),
.B(n_1468),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1517),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1527),
.Y(n_1551)
);

OAI21xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1526),
.A2(n_1496),
.B(n_1479),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1515),
.B(n_1488),
.Y(n_1553)
);

OR2x6_ASAP7_75t_L g1554 ( 
.A(n_1514),
.B(n_1470),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1515),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1527),
.B(n_1433),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1501),
.Y(n_1557)
);

OR2x6_ASAP7_75t_L g1558 ( 
.A(n_1515),
.B(n_1470),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1527),
.B(n_1433),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1526),
.A2(n_1461),
.B1(n_1451),
.B2(n_1425),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1520),
.Y(n_1561)
);

INVxp67_ASAP7_75t_SL g1562 ( 
.A(n_1505),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1516),
.B(n_1481),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1516),
.B(n_1425),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1529),
.B(n_1483),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1520),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1547),
.Y(n_1567)
);

XNOR2xp5_ASAP7_75t_L g1568 ( 
.A(n_1546),
.B(n_1290),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1530),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1531),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1550),
.B(n_1519),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1545),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1532),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1545),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1538),
.B(n_1516),
.Y(n_1575)
);

AO21x1_ASAP7_75t_L g1576 ( 
.A1(n_1543),
.A2(n_1519),
.B(n_1521),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1541),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1538),
.B(n_1516),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1534),
.B(n_1516),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1535),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1537),
.B(n_1505),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1557),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1562),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1536),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1534),
.B(n_1536),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1562),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1536),
.B(n_1518),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1557),
.Y(n_1588)
);

AND2x2_ASAP7_75t_SL g1589 ( 
.A(n_1565),
.B(n_1521),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1554),
.A2(n_1471),
.B1(n_1478),
.B2(n_1528),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1537),
.B(n_1555),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1537),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1561),
.B(n_1566),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1543),
.A2(n_1528),
.B(n_1472),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1551),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1549),
.Y(n_1596)
);

NOR2x1_ASAP7_75t_L g1597 ( 
.A(n_1554),
.B(n_1508),
.Y(n_1597)
);

INVxp67_ASAP7_75t_SL g1598 ( 
.A(n_1540),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1556),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1559),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1558),
.B(n_1518),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1558),
.B(n_1518),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1539),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1548),
.B(n_1511),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1555),
.B(n_1508),
.Y(n_1605)
);

OR2x6_ASAP7_75t_L g1606 ( 
.A(n_1544),
.B(n_1554),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_SL g1607 ( 
.A(n_1544),
.B(n_1390),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1553),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1544),
.A2(n_1387),
.B(n_1506),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1558),
.B(n_1509),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1585),
.B(n_1533),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1605),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1589),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1571),
.B(n_1506),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1568),
.B(n_1390),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1577),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1589),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1571),
.B(n_1513),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1568),
.B(n_1347),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1585),
.B(n_1533),
.Y(n_1620)
);

AND2x4_ASAP7_75t_SL g1621 ( 
.A(n_1606),
.B(n_1584),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1589),
.B(n_1552),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1569),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1590),
.A2(n_1560),
.B(n_1563),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1597),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1569),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1605),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1601),
.B(n_1564),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1605),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1570),
.Y(n_1630)
);

INVxp67_ASAP7_75t_L g1631 ( 
.A(n_1607),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1567),
.B(n_1511),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1605),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1567),
.B(n_1513),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1587),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1570),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1590),
.A2(n_1563),
.B1(n_1553),
.B2(n_1443),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1573),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_SL g1639 ( 
.A(n_1607),
.B(n_1484),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1573),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1594),
.A2(n_1553),
.B1(n_1443),
.B2(n_1430),
.Y(n_1641)
);

OR2x6_ASAP7_75t_L g1642 ( 
.A(n_1606),
.B(n_1386),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1580),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1577),
.B(n_1599),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1599),
.B(n_1600),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1606),
.Y(n_1646)
);

AOI31xp33_ASAP7_75t_L g1647 ( 
.A1(n_1622),
.A2(n_1576),
.A3(n_1597),
.B(n_1594),
.Y(n_1647)
);

OAI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1639),
.A2(n_1606),
.B1(n_1609),
.B2(n_1584),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1616),
.B(n_1603),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1645),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1624),
.A2(n_1576),
.B1(n_1606),
.B2(n_1603),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1645),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1637),
.A2(n_1606),
.B1(n_1609),
.B2(n_1598),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1611),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1644),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_SL g1656 ( 
.A(n_1613),
.B(n_1608),
.C(n_1600),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1617),
.B(n_1598),
.Y(n_1657)
);

AO22x1_ASAP7_75t_L g1658 ( 
.A1(n_1625),
.A2(n_1592),
.B1(n_1591),
.B2(n_1586),
.Y(n_1658)
);

AOI21xp33_ASAP7_75t_L g1659 ( 
.A1(n_1625),
.A2(n_1586),
.B(n_1583),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1621),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1644),
.B(n_1599),
.Y(n_1661)
);

AOI211xp5_ASAP7_75t_L g1662 ( 
.A1(n_1631),
.A2(n_1583),
.B(n_1608),
.C(n_1600),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1636),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1646),
.B(n_1604),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1636),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1635),
.B(n_1596),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1611),
.B(n_1596),
.Y(n_1667)
);

NAND3xp33_ASAP7_75t_SL g1668 ( 
.A(n_1641),
.B(n_1620),
.C(n_1615),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1638),
.Y(n_1669)
);

AOI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1619),
.A2(n_1608),
.B(n_1593),
.C(n_1592),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1620),
.B(n_1593),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1628),
.B(n_1635),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1651),
.A2(n_1621),
.B1(n_1642),
.B2(n_1584),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1647),
.A2(n_1632),
.B(n_1642),
.Y(n_1674)
);

AOI222xp33_ASAP7_75t_L g1675 ( 
.A1(n_1656),
.A2(n_1626),
.B1(n_1623),
.B2(n_1630),
.C1(n_1638),
.C2(n_1643),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1655),
.B(n_1662),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1653),
.A2(n_1642),
.B1(n_1584),
.B2(n_1601),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1661),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1649),
.B(n_1654),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1650),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1670),
.B(n_1628),
.Y(n_1681)
);

NOR2x1_ASAP7_75t_L g1682 ( 
.A(n_1647),
.B(n_1642),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1648),
.B(n_1618),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1672),
.B(n_1652),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1668),
.B(n_1660),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1663),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1658),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1660),
.B(n_1575),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1664),
.B(n_1634),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1657),
.B(n_1634),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1665),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1671),
.B(n_1347),
.Y(n_1692)
);

AOI211xp5_ASAP7_75t_L g1693 ( 
.A1(n_1673),
.A2(n_1653),
.B(n_1659),
.C(n_1667),
.Y(n_1693)
);

OAI211xp5_ASAP7_75t_L g1694 ( 
.A1(n_1682),
.A2(n_1659),
.B(n_1669),
.C(n_1666),
.Y(n_1694)
);

A2O1A1Ixp33_ASAP7_75t_L g1695 ( 
.A1(n_1674),
.A2(n_1618),
.B(n_1591),
.C(n_1592),
.Y(n_1695)
);

OAI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1676),
.A2(n_1643),
.B1(n_1640),
.B2(n_1633),
.C(n_1629),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1687),
.A2(n_1640),
.B1(n_1633),
.B2(n_1629),
.C(n_1627),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1685),
.B(n_1587),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1687),
.A2(n_1627),
.B(n_1612),
.Y(n_1699)
);

AOI21xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1675),
.A2(n_1342),
.B(n_1250),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1677),
.A2(n_1612),
.B(n_1591),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1692),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1683),
.A2(n_1591),
.B1(n_1614),
.B2(n_1581),
.C(n_1580),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1692),
.B(n_1250),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1702),
.B(n_1678),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1699),
.B(n_1681),
.Y(n_1706)
);

NOR2x1p5_ASAP7_75t_SL g1707 ( 
.A(n_1694),
.B(n_1679),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1698),
.B(n_1689),
.Y(n_1708)
);

XOR2x2_ASAP7_75t_L g1709 ( 
.A(n_1704),
.B(n_1684),
.Y(n_1709)
);

NAND2x1_ASAP7_75t_SL g1710 ( 
.A(n_1700),
.B(n_1688),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1697),
.Y(n_1711)
);

XNOR2xp5_ASAP7_75t_L g1712 ( 
.A(n_1693),
.B(n_1690),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1696),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_L g1714 ( 
.A(n_1703),
.B(n_1680),
.C(n_1686),
.Y(n_1714)
);

INVx2_ASAP7_75t_SL g1715 ( 
.A(n_1701),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1695),
.B(n_1575),
.Y(n_1716)
);

NOR3xp33_ASAP7_75t_L g1717 ( 
.A(n_1705),
.B(n_1691),
.C(n_1524),
.Y(n_1717)
);

NOR4xp25_ASAP7_75t_L g1718 ( 
.A(n_1711),
.B(n_1614),
.C(n_1588),
.D(n_1582),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1708),
.B(n_1604),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1707),
.B(n_1610),
.Y(n_1720)
);

NOR3xp33_ASAP7_75t_L g1721 ( 
.A(n_1706),
.B(n_1321),
.C(n_1581),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1715),
.B(n_1581),
.Y(n_1722)
);

NAND3xp33_ASAP7_75t_SL g1723 ( 
.A(n_1711),
.B(n_1610),
.C(n_1602),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1719),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_L g1725 ( 
.A(n_1720),
.B(n_1723),
.Y(n_1725)
);

INVxp67_ASAP7_75t_L g1726 ( 
.A(n_1722),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1718),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1717),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1721),
.A2(n_1712),
.B1(n_1716),
.B2(n_1713),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1719),
.Y(n_1730)
);

NOR2xp67_ASAP7_75t_L g1731 ( 
.A(n_1726),
.B(n_1714),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1725),
.B(n_1728),
.Y(n_1732)
);

OAI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1729),
.A2(n_1710),
.B1(n_1709),
.B2(n_1602),
.C(n_1572),
.Y(n_1733)
);

NOR3xp33_ASAP7_75t_L g1734 ( 
.A(n_1724),
.B(n_1321),
.C(n_1581),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1727),
.A2(n_1595),
.B1(n_1588),
.B2(n_1582),
.Y(n_1735)
);

AND4x1_ASAP7_75t_L g1736 ( 
.A(n_1730),
.B(n_1578),
.C(n_1579),
.D(n_1595),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1732),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1731),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1733),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1737),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1740),
.B(n_1738),
.C(n_1739),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1741),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1741),
.A2(n_1734),
.B1(n_1739),
.B2(n_1735),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1743),
.A2(n_1736),
.B1(n_1588),
.B2(n_1582),
.Y(n_1744)
);

AOI21xp33_ASAP7_75t_SL g1745 ( 
.A1(n_1742),
.A2(n_1574),
.B(n_1572),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1744),
.A2(n_1574),
.B(n_1572),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1745),
.B(n_1578),
.Y(n_1747)
);

OA21x2_ASAP7_75t_L g1748 ( 
.A1(n_1746),
.A2(n_1574),
.B(n_1579),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1747),
.B1(n_1507),
.B2(n_1501),
.Y(n_1749)
);

OAI221xp5_ASAP7_75t_R g1750 ( 
.A1(n_1749),
.A2(n_1507),
.B1(n_1278),
.B2(n_1498),
.C(n_1542),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1507),
.B(n_1404),
.C(n_1512),
.Y(n_1751)
);


endmodule