module fake_netlist_6_4157_n_2159 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_422, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2159);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_422;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2159;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1371;
wire n_1285;
wire n_461;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_1815;
wire n_659;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1605;
wire n_1413;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_928;
wire n_835;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_437;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_458;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_623;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_527;
wire n_683;
wire n_1207;
wire n_474;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_1092;
wire n_441;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2052;
wire n_1847;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_621;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_1642;
wire n_711;
wire n_1352;
wire n_579;
wire n_937;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_523;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_611;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_1737;
wire n_653;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_1028;
wire n_576;
wire n_2106;
wire n_472;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_924;
wire n_475;
wire n_1582;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1888;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_1322;
wire n_640;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_629;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_1025;
wire n_2116;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_1742;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_411),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_271),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g427 ( 
.A(n_156),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_319),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_277),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_350),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_153),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_160),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_383),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_34),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_114),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_41),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_420),
.Y(n_437)
);

BUFx5_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_176),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_3),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_8),
.Y(n_441)
);

BUFx5_ASAP7_75t_L g442 ( 
.A(n_408),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_140),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_400),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_385),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_276),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_399),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_13),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_78),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_397),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_173),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_216),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_327),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_222),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_72),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_101),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_310),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_121),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_170),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_177),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_105),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_183),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_387),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_45),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_7),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_370),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_118),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_320),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_28),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_417),
.Y(n_470)
);

BUFx4f_ASAP7_75t_SL g471 ( 
.A(n_169),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_81),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_326),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_334),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_412),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_287),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_114),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_262),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_421),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_164),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_274),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_172),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_414),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_366),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_9),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_188),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_65),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_410),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_209),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_224),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_120),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_290),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_18),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_226),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_192),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_265),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_126),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_130),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_416),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_375),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_357),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_51),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_73),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_419),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_390),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_159),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_344),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_382),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_188),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_106),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_294),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_377),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_130),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_314),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_315),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_104),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_39),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_339),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_61),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_398),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_278),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_203),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_14),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_337),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_168),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_313),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_353),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_346),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_361),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_152),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_172),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_193),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_86),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_378),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_345),
.Y(n_535)
);

BUFx5_ASAP7_75t_L g536 ( 
.A(n_71),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_422),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_219),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_58),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_405),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_325),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_272),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_20),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_354),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_175),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_137),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_379),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_247),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_312),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_365),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_128),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_39),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_54),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_311),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_181),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_57),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_121),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_289),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_15),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_49),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_369),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_248),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_233),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_156),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_388),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_262),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_51),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_214),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_415),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_6),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_367),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_309),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_371),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_186),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_44),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_275),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_195),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_98),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_183),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_26),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_391),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_241),
.Y(n_582)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_360),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_259),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_324),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_396),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_393),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_84),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_47),
.Y(n_589)
);

CKINVDCx16_ASAP7_75t_R g590 ( 
.A(n_205),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_331),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_243),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_100),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_112),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_373),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_280),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_189),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_313),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_177),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_347),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_418),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_368),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_49),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_119),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_66),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_122),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_340),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_233),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_128),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_364),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_56),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_212),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_230),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_189),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_1),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_348),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_261),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_424),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_25),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_402),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_94),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_118),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_104),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_90),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_305),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_279),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_253),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_318),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_5),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_26),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_242),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_240),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_363),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_423),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_352),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_7),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_29),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_332),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_376),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_34),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_21),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_106),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_166),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_20),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_72),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_137),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_264),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_146),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_335),
.Y(n_649)
);

INVxp33_ASAP7_75t_SL g650 ( 
.A(n_342),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_161),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_292),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_209),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_92),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_374),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_236),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_90),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_1),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_317),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_351),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_24),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_358),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_27),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_401),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_386),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_322),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_270),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_292),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_273),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_142),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_86),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_349),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_329),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_151),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_355),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_101),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_343),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_89),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_143),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_275),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_91),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_305),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_151),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_48),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_73),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_171),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_333),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_381),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_253),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_50),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_55),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_237),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_47),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_409),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_301),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_228),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_234),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_389),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_323),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_68),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_321),
.Y(n_701)
);

BUFx8_ASAP7_75t_SL g702 ( 
.A(n_71),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_359),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_296),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_336),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_247),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_229),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_111),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_175),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_164),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_301),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_107),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_356),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_395),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_372),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_330),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_4),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_403),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_59),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_105),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_302),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_404),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_143),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_41),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_380),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_338),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_145),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_413),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_394),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_85),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_328),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_286),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_3),
.Y(n_733)
);

CKINVDCx12_ASAP7_75t_R g734 ( 
.A(n_5),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_269),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_97),
.Y(n_736)
);

CKINVDCx14_ASAP7_75t_R g737 ( 
.A(n_46),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_36),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_392),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_407),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_75),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_19),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_12),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_308),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_265),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_147),
.Y(n_746)
);

INVxp33_ASAP7_75t_SL g747 ( 
.A(n_88),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_170),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_362),
.Y(n_749)
);

BUFx10_ASAP7_75t_L g750 ( 
.A(n_384),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_406),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_213),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_13),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_244),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_258),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_702),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_536),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_658),
.Y(n_758)
);

INVxp33_ASAP7_75t_L g759 ( 
.A(n_456),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_427),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_470),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_536),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_564),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_462),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_536),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_564),
.Y(n_766)
);

CKINVDCx16_ASAP7_75t_R g767 ( 
.A(n_542),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_591),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_536),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_536),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_536),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_737),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_734),
.Y(n_773)
);

INVxp33_ASAP7_75t_SL g774 ( 
.A(n_429),
.Y(n_774)
);

CKINVDCx16_ASAP7_75t_R g775 ( 
.A(n_580),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_590),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_536),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_536),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_564),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_688),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_509),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_498),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_509),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_429),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_489),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_549),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_490),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_436),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_492),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_549),
.Y(n_790)
);

INVxp33_ASAP7_75t_SL g791 ( 
.A(n_431),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_652),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_652),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_684),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_595),
.Y(n_795)
);

INVxp67_ASAP7_75t_SL g796 ( 
.A(n_587),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_684),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_431),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_709),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_709),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_493),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_436),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_436),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_436),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_587),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_494),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_636),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_436),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_496),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_568),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_568),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_568),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_716),
.B(n_0),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_568),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_568),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_614),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_614),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_614),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_614),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_510),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_614),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_619),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_619),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_497),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_619),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_619),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_663),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_503),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_663),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_795),
.Y(n_830)
);

BUFx12f_ASAP7_75t_L g831 ( 
.A(n_760),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_788),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_795),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_788),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_795),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_802),
.B(n_620),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_795),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_803),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_760),
.B(n_583),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_772),
.B(n_750),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_795),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_768),
.A2(n_434),
.B1(n_435),
.B2(n_432),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_757),
.A2(n_534),
.B(n_518),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_804),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_808),
.B(n_620),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_780),
.A2(n_434),
.B1(n_435),
.B2(n_432),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_810),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_811),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_796),
.B(n_665),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_812),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_814),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_772),
.B(n_650),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_815),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_816),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_817),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_SL g856 ( 
.A(n_764),
.B(n_672),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_813),
.B(n_716),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_818),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_819),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_756),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_776),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_821),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_822),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_823),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_825),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_SL g866 ( 
.A1(n_782),
.A2(n_558),
.B1(n_559),
.B2(n_530),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_805),
.B(n_761),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_826),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_827),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_829),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_758),
.A2(n_643),
.B1(n_661),
.B2(n_592),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_781),
.B(n_665),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_762),
.A2(n_534),
.B(n_518),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_783),
.B(n_449),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_765),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_769),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_770),
.B(n_713),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_771),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_SL g879 ( 
.A1(n_782),
.A2(n_710),
.B1(n_719),
.B2(n_689),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_777),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_778),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_799),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_786),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_790),
.Y(n_884)
);

OA21x2_ASAP7_75t_L g885 ( 
.A1(n_792),
.A2(n_586),
.B(n_581),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_793),
.B(n_713),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_794),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_797),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_800),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_756),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_860),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_834),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_860),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_834),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_831),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_866),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_R g897 ( 
.A(n_890),
.B(n_785),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_875),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_890),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_831),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_833),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_875),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_838),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_877),
.B(n_878),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_838),
.Y(n_905)
);

CKINVDCx16_ASAP7_75t_R g906 ( 
.A(n_856),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_866),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_833),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_861),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_878),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_844),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_882),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_852),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_844),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_881),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_867),
.B(n_774),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_882),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_R g918 ( 
.A(n_849),
.B(n_785),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_848),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_R g920 ( 
.A(n_881),
.B(n_787),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_879),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_879),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_871),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_871),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_839),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_863),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_833),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_848),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_840),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_833),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_863),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_842),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_874),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_846),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_833),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_857),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_863),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_850),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_857),
.Y(n_939)
);

XOR2xp5_ASAP7_75t_L g940 ( 
.A(n_877),
.B(n_820),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_857),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_R g942 ( 
.A(n_888),
.B(n_787),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_876),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_857),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_857),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_876),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_874),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_884),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_892),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_912),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_916),
.B(n_913),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_926),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_898),
.B(n_877),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_933),
.B(n_774),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_931),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_937),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_902),
.B(n_877),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_904),
.B(n_595),
.Y(n_958)
);

BUFx10_ASAP7_75t_L g959 ( 
.A(n_895),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_910),
.Y(n_960)
);

NOR2x1_ASAP7_75t_L g961 ( 
.A(n_947),
.B(n_468),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_915),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_948),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_947),
.B(n_791),
.Y(n_964)
);

INVx5_ASAP7_75t_L g965 ( 
.A(n_901),
.Y(n_965)
);

INVx3_ASAP7_75t_R g966 ( 
.A(n_900),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_943),
.B(n_886),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_917),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_892),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_903),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_891),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_946),
.B(n_880),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_903),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_920),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_905),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_905),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_893),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_901),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_894),
.Y(n_979)
);

INVxp67_ASAP7_75t_SL g980 ( 
.A(n_901),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_911),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_894),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_929),
.A2(n_504),
.B1(n_602),
.B2(n_529),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_911),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_901),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_940),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_908),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_914),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_918),
.B(n_880),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_942),
.B(n_936),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_914),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_939),
.B(n_595),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_908),
.B(n_927),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_919),
.Y(n_994)
);

INVx5_ASAP7_75t_L g995 ( 
.A(n_908),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_909),
.B(n_789),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_932),
.B(n_791),
.Y(n_997)
);

AND2x6_ASAP7_75t_L g998 ( 
.A(n_919),
.B(n_581),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_927),
.B(n_836),
.Y(n_999)
);

AND2x6_ASAP7_75t_L g1000 ( 
.A(n_928),
.B(n_586),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_928),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_897),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_899),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_925),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_938),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_938),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_927),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_930),
.B(n_836),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_930),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_930),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_935),
.B(n_836),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_935),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_935),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_923),
.A2(n_885),
.B1(n_747),
.B2(n_553),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_941),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_945),
.Y(n_1016)
);

INVx4_ASAP7_75t_SL g1017 ( 
.A(n_944),
.Y(n_1017)
);

AND2x6_ASAP7_75t_SL g1018 ( 
.A(n_896),
.B(n_426),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_934),
.B(n_789),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_925),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_906),
.B(n_801),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_944),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_924),
.B(n_595),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_895),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_921),
.A2(n_885),
.B1(n_747),
.B2(n_553),
.Y(n_1025)
);

AND2x6_ASAP7_75t_L g1026 ( 
.A(n_922),
.B(n_638),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_1014),
.A2(n_650),
.B1(n_715),
.B2(n_638),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_951),
.B(n_801),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_963),
.B(n_951),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_954),
.A2(n_635),
.B1(n_749),
.B2(n_677),
.Y(n_1030)
);

AO22x2_ASAP7_75t_L g1031 ( 
.A1(n_1023),
.A2(n_472),
.B1(n_556),
.B2(n_449),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1001),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1001),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_979),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_962),
.B(n_886),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_960),
.B(n_806),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_1025),
.A2(n_731),
.B1(n_751),
.B2(n_715),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_970),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_962),
.B(n_886),
.Y(n_1039)
);

AND2x6_ASAP7_75t_L g1040 ( 
.A(n_952),
.B(n_731),
.Y(n_1040)
);

AND2x6_ASAP7_75t_L g1041 ( 
.A(n_955),
.B(n_751),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_954),
.Y(n_1042)
);

NAND2x1p5_ASAP7_75t_L g1043 ( 
.A(n_963),
.B(n_888),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_979),
.Y(n_1044)
);

NAND2x1p5_ASAP7_75t_L g1045 ( 
.A(n_950),
.B(n_888),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_973),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_975),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_976),
.Y(n_1048)
);

BUFx8_ASAP7_75t_L g1049 ( 
.A(n_1002),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_989),
.B(n_806),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_981),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_950),
.B(n_784),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_982),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_988),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_994),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_956),
.B(n_809),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1005),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_1020),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_984),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_967),
.B(n_886),
.Y(n_1060)
);

BUFx8_ASAP7_75t_L g1061 ( 
.A(n_968),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_967),
.B(n_883),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_994),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1016),
.B(n_883),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_991),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1025),
.B(n_809),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1006),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_953),
.B(n_824),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_949),
.Y(n_1069)
);

AND2x2_ASAP7_75t_SL g1070 ( 
.A(n_997),
.B(n_767),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1019),
.B(n_798),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_974),
.B(n_775),
.Y(n_1072)
);

OR2x6_ASAP7_75t_SL g1073 ( 
.A(n_1022),
.B(n_776),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_949),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_957),
.B(n_824),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1019),
.A2(n_845),
.B1(n_836),
.B2(n_828),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_969),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_969),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_980),
.B(n_828),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1012),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_1016),
.B(n_887),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1012),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_996),
.B(n_884),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_1004),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_997),
.B(n_884),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1009),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1010),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_961),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_985),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_1015),
.B(n_887),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1013),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_983),
.B(n_820),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_972),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_999),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_1015),
.B(n_889),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1008),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1011),
.Y(n_1097)
);

INVxp67_ASAP7_75t_L g1098 ( 
.A(n_964),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1026),
.A2(n_845),
.B1(n_699),
.B2(n_610),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_993),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1017),
.B(n_889),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_964),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_980),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_971),
.B(n_759),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_971),
.B(n_759),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1014),
.B(n_884),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_1023),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_987),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_987),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1007),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1007),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_985),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_1021),
.B(n_884),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1026),
.B(n_845),
.Y(n_1114)
);

OAI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_992),
.A2(n_896),
.B1(n_907),
.B2(n_872),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_985),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_985),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1017),
.B(n_990),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1017),
.B(n_990),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_978),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_965),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_1026),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_992),
.B(n_845),
.Y(n_1123)
);

NAND2x1p5_ASAP7_75t_L g1124 ( 
.A(n_977),
.B(n_1003),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_998),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_978),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1026),
.A2(n_466),
.B1(n_473),
.B2(n_444),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_977),
.B(n_1003),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1093),
.B(n_1026),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1094),
.A2(n_958),
.B(n_873),
.Y(n_1130)
);

NOR3xp33_ASAP7_75t_L g1131 ( 
.A(n_1092),
.B(n_1021),
.C(n_1028),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1108),
.A2(n_965),
.B(n_958),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1096),
.A2(n_873),
.B(n_843),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1093),
.B(n_995),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1042),
.B(n_1024),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1079),
.B(n_959),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1071),
.B(n_763),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1098),
.B(n_986),
.Y(n_1138)
);

O2A1O1Ixp5_ASAP7_75t_L g1139 ( 
.A1(n_1113),
.A2(n_499),
.B(n_527),
.C(n_505),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1107),
.B(n_995),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1068),
.B(n_995),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1126),
.A2(n_965),
.B(n_885),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1126),
.A2(n_885),
.B(n_841),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1082),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1097),
.A2(n_841),
.B(n_835),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_SL g1146 ( 
.A(n_1128),
.B(n_959),
.Y(n_1146)
);

OAI21xp33_ASAP7_75t_L g1147 ( 
.A1(n_1027),
.A2(n_1066),
.B(n_1037),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1125),
.A2(n_843),
.B(n_865),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1075),
.B(n_447),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1050),
.B(n_701),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1100),
.B(n_847),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1123),
.A2(n_907),
.B1(n_714),
.B2(n_541),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1076),
.A2(n_528),
.B(n_561),
.C(n_550),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1036),
.B(n_1102),
.C(n_1029),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_1128),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1103),
.B(n_847),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1106),
.A2(n_1000),
.B(n_998),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_1089),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1030),
.A2(n_986),
.B1(n_484),
.B2(n_488),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1114),
.A2(n_841),
.B(n_835),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_1089),
.B(n_837),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1111),
.A2(n_841),
.B(n_835),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1109),
.A2(n_841),
.B(n_835),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1035),
.B(n_854),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1056),
.A2(n_556),
.B(n_567),
.C(n_472),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1110),
.A2(n_835),
.B(n_830),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1082),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1035),
.B(n_425),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1032),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1039),
.B(n_854),
.Y(n_1170)
);

NOR3xp33_ASAP7_75t_L g1171 ( 
.A(n_1115),
.B(n_779),
.C(n_766),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_1121),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1122),
.A2(n_1099),
.B1(n_1046),
.B2(n_1047),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1084),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1032),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1085),
.A2(n_567),
.B(n_679),
.C(n_593),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1039),
.B(n_858),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1031),
.B(n_858),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1031),
.B(n_862),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1121),
.A2(n_1060),
.B(n_1120),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1038),
.B(n_862),
.Y(n_1181)
);

OAI21xp33_ASAP7_75t_L g1182 ( 
.A1(n_1127),
.A2(n_446),
.B(n_443),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1048),
.B(n_865),
.Y(n_1183)
);

AO32x1_ASAP7_75t_L g1184 ( 
.A1(n_1086),
.A2(n_593),
.A3(n_745),
.B1(n_679),
.B2(n_603),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1121),
.A2(n_830),
.B(n_837),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1104),
.B(n_807),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1051),
.B(n_868),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1033),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1033),
.Y(n_1189)
);

O2A1O1Ixp5_ASAP7_75t_L g1190 ( 
.A1(n_1083),
.A2(n_565),
.B(n_601),
.C(n_600),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1101),
.B(n_1064),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1086),
.A2(n_832),
.B(n_868),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1123),
.A2(n_714),
.B1(n_616),
.B2(n_628),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1058),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1070),
.A2(n_500),
.B1(n_501),
.B2(n_483),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1089),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1054),
.B(n_869),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1116),
.A2(n_1062),
.B(n_1117),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1116),
.A2(n_830),
.B(n_607),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_SL g1200 ( 
.A(n_1124),
.B(n_966),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1062),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1057),
.B(n_869),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1064),
.B(n_1000),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1081),
.B(n_425),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1112),
.B(n_595),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1077),
.A2(n_662),
.B(n_607),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1081),
.B(n_998),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1077),
.A2(n_662),
.B(n_607),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1034),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1044),
.A2(n_662),
.B(n_607),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1101),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1105),
.B(n_799),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1052),
.B(n_1018),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1053),
.A2(n_662),
.B(n_607),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1059),
.B(n_998),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1080),
.A2(n_687),
.B(n_662),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1087),
.Y(n_1217)
);

INVx4_ASAP7_75t_L g1218 ( 
.A(n_1118),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1088),
.A2(n_508),
.B1(n_512),
.B2(n_507),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1049),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1055),
.A2(n_687),
.B(n_634),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1125),
.A2(n_851),
.B(n_850),
.Y(n_1222)
);

AOI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1087),
.A2(n_832),
.B(n_851),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1131),
.B(n_1090),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1138),
.B(n_1072),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1142),
.A2(n_1043),
.B(n_1063),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1149),
.B(n_1118),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1191),
.B(n_1119),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1222),
.A2(n_1091),
.B(n_1067),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1147),
.A2(n_1119),
.B(n_1090),
.C(n_1095),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1155),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1150),
.B(n_1095),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1141),
.A2(n_1074),
.B(n_1069),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1137),
.B(n_1065),
.Y(n_1234)
);

OA22x2_ASAP7_75t_L g1235 ( 
.A1(n_1159),
.A2(n_773),
.B1(n_464),
.B2(n_477),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1144),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1212),
.B(n_1045),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1174),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_1172),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1147),
.A2(n_1078),
.B(n_664),
.C(n_673),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1194),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1191),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1167),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_R g1244 ( 
.A(n_1146),
.B(n_1049),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1130),
.A2(n_687),
.B(n_1040),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1217),
.Y(n_1246)
);

CKINVDCx8_ASAP7_75t_R g1247 ( 
.A(n_1220),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1169),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1154),
.A2(n_698),
.B(n_703),
.C(n_694),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1132),
.A2(n_687),
.B(n_1040),
.Y(n_1250)
);

NOR3xp33_ASAP7_75t_L g1251 ( 
.A(n_1171),
.B(n_745),
.C(n_647),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1186),
.B(n_1040),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1201),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1135),
.B(n_1073),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1213),
.B(n_1061),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1218),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_SL g1257 ( 
.A1(n_1129),
.A2(n_718),
.B(n_722),
.C(n_705),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1198),
.A2(n_687),
.B(n_1040),
.Y(n_1258)
);

NOR2x1_ASAP7_75t_L g1259 ( 
.A(n_1134),
.B(n_725),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1189),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1157),
.A2(n_1041),
.B(n_739),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_R g1262 ( 
.A(n_1200),
.B(n_1061),
.Y(n_1262)
);

INVx6_ASAP7_75t_L g1263 ( 
.A(n_1211),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1175),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1152),
.B(n_1041),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1188),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1204),
.B(n_721),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1148),
.A2(n_726),
.B(n_855),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1172),
.B(n_855),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1172),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1201),
.B(n_1041),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1143),
.A2(n_1041),
.B(n_520),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_SL g1273 ( 
.A(n_1218),
.B(n_724),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1211),
.B(n_735),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1173),
.A2(n_752),
.B1(n_738),
.B2(n_1000),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1219),
.B(n_672),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_SL g1277 ( 
.A1(n_1153),
.A2(n_700),
.B(n_706),
.C(n_546),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1193),
.A2(n_430),
.B1(n_433),
.B2(n_428),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1158),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1151),
.B(n_727),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1164),
.B(n_730),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1170),
.B(n_1177),
.Y(n_1282)
);

BUFx2_ASAP7_75t_SL g1283 ( 
.A(n_1158),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_L g1284 ( 
.A(n_1165),
.B(n_511),
.C(n_506),
.Y(n_1284)
);

CKINVDCx8_ASAP7_75t_R g1285 ( 
.A(n_1158),
.Y(n_1285)
);

NOR3xp33_ASAP7_75t_L g1286 ( 
.A(n_1136),
.B(n_487),
.C(n_454),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1196),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1203),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1207),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1178),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1179),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1133),
.A2(n_535),
.B(n_524),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_R g1293 ( 
.A(n_1209),
.B(n_428),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1195),
.B(n_672),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1168),
.B(n_636),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1180),
.A2(n_540),
.B(n_537),
.Y(n_1296)
);

OAI21xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1181),
.A2(n_576),
.B(n_491),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1140),
.B(n_471),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1192),
.Y(n_1299)
);

NOR3xp33_ASAP7_75t_SL g1300 ( 
.A(n_1182),
.B(n_440),
.C(n_439),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1182),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_SL g1302 ( 
.A(n_1176),
.B(n_750),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1139),
.A2(n_457),
.B(n_458),
.C(n_452),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1160),
.A2(n_547),
.B(n_544),
.Y(n_1304)
);

BUFx12f_ASAP7_75t_L g1305 ( 
.A(n_1161),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1183),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1223),
.A2(n_1145),
.B(n_1163),
.Y(n_1307)
);

AOI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1166),
.A2(n_864),
.B(n_859),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1187),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1161),
.Y(n_1310)
);

OR2x6_ASAP7_75t_SL g1311 ( 
.A(n_1197),
.B(n_439),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_R g1312 ( 
.A(n_1215),
.B(n_430),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1156),
.A2(n_571),
.B(n_569),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1202),
.A2(n_585),
.B(n_573),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1190),
.A2(n_1000),
.B(n_864),
.Y(n_1315)
);

NOR2xp67_ASAP7_75t_L g1316 ( 
.A(n_1185),
.B(n_316),
.Y(n_1316)
);

AND2x6_ASAP7_75t_L g1317 ( 
.A(n_1184),
.B(n_491),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1205),
.B(n_433),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1205),
.B(n_437),
.Y(n_1319)
);

NAND2x1p5_ASAP7_75t_L g1320 ( 
.A(n_1239),
.B(n_1199),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1247),
.Y(n_1321)
);

CKINVDCx16_ASAP7_75t_R g1322 ( 
.A(n_1244),
.Y(n_1322)
);

OR2x6_ASAP7_75t_L g1323 ( 
.A(n_1230),
.B(n_1206),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1242),
.B(n_1162),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1246),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1260),
.Y(n_1326)
);

BUFx8_ASAP7_75t_L g1327 ( 
.A(n_1231),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1285),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1287),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1241),
.Y(n_1330)
);

INVxp33_ASAP7_75t_L g1331 ( 
.A(n_1225),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1266),
.Y(n_1332)
);

INVx5_ASAP7_75t_L g1333 ( 
.A(n_1239),
.Y(n_1333)
);

BUFx8_ASAP7_75t_L g1334 ( 
.A(n_1279),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1279),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1238),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1270),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1236),
.Y(n_1338)
);

INVx4_ASAP7_75t_L g1339 ( 
.A(n_1270),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1309),
.B(n_1208),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1279),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1263),
.Y(n_1342)
);

INVx5_ASAP7_75t_L g1343 ( 
.A(n_1287),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1262),
.Y(n_1344)
);

INVx1_ASAP7_75t_SL g1345 ( 
.A(n_1306),
.Y(n_1345)
);

INVx8_ASAP7_75t_L g1346 ( 
.A(n_1305),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1290),
.B(n_750),
.Y(n_1347)
);

BUFx4_ASAP7_75t_SL g1348 ( 
.A(n_1256),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1291),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1287),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1243),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1228),
.B(n_437),
.Y(n_1352)
);

INVx4_ASAP7_75t_L g1353 ( 
.A(n_1269),
.Y(n_1353)
);

INVx4_ASAP7_75t_L g1354 ( 
.A(n_1289),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1293),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1237),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1248),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1267),
.B(n_445),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1253),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1264),
.Y(n_1360)
);

AND2x6_ASAP7_75t_L g1361 ( 
.A(n_1289),
.B(n_1184),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1311),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1288),
.Y(n_1363)
);

BUFx12f_ASAP7_75t_L g1364 ( 
.A(n_1301),
.Y(n_1364)
);

INVxp67_ASAP7_75t_SL g1365 ( 
.A(n_1299),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1282),
.B(n_1000),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_SL g1367 ( 
.A(n_1317),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1310),
.Y(n_1368)
);

CKINVDCx16_ASAP7_75t_R g1369 ( 
.A(n_1273),
.Y(n_1369)
);

BUFx8_ASAP7_75t_L g1370 ( 
.A(n_1295),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1234),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1229),
.Y(n_1372)
);

BUFx2_ASAP7_75t_SL g1373 ( 
.A(n_1274),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_1227),
.Y(n_1374)
);

INVxp67_ASAP7_75t_SL g1375 ( 
.A(n_1224),
.Y(n_1375)
);

INVx4_ASAP7_75t_L g1376 ( 
.A(n_1283),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1232),
.B(n_1221),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1251),
.A2(n_516),
.B1(n_519),
.B2(n_513),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1255),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1275),
.A2(n_717),
.B1(n_636),
.B2(n_603),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1240),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1280),
.B(n_445),
.Y(n_1382)
);

INVx3_ASAP7_75t_SL g1383 ( 
.A(n_1235),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1317),
.Y(n_1384)
);

BUFx4f_ASAP7_75t_SL g1385 ( 
.A(n_1276),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1254),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1271),
.Y(n_1387)
);

INVx6_ASAP7_75t_SL g1388 ( 
.A(n_1286),
.Y(n_1388)
);

BUFx12f_ASAP7_75t_L g1389 ( 
.A(n_1317),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1312),
.Y(n_1390)
);

INVx6_ASAP7_75t_SL g1391 ( 
.A(n_1297),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1252),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1259),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1259),
.Y(n_1394)
);

BUFx4_ASAP7_75t_SL g1395 ( 
.A(n_1284),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1372),
.A2(n_1245),
.B(n_1261),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1358),
.A2(n_1294),
.B(n_1298),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1321),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1349),
.B(n_1281),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1380),
.A2(n_1275),
.B(n_1300),
.C(n_1297),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1325),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1326),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1332),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1372),
.A2(n_1307),
.B(n_1268),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1365),
.A2(n_1250),
.B(n_1258),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1331),
.B(n_1277),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1320),
.A2(n_1308),
.B(n_1226),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1323),
.A2(n_1272),
.B(n_1292),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1382),
.A2(n_1380),
.B(n_1378),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1365),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1320),
.A2(n_1233),
.B(n_1216),
.Y(n_1411)
);

NAND3xp33_ASAP7_75t_L g1412 ( 
.A(n_1378),
.B(n_1302),
.C(n_1249),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1366),
.A2(n_1214),
.B(n_1210),
.Y(n_1413)
);

O2A1O1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1383),
.A2(n_1265),
.B(n_1278),
.C(n_1303),
.Y(n_1414)
);

OR2x6_ASAP7_75t_L g1415 ( 
.A(n_1323),
.B(n_1316),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1381),
.A2(n_1315),
.B(n_1304),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1374),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1374),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1338),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1366),
.A2(n_1296),
.B(n_1318),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1349),
.B(n_1319),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1340),
.A2(n_1313),
.B(n_859),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1351),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1357),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1371),
.B(n_1314),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1371),
.B(n_755),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1360),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1327),
.Y(n_1428)
);

AOI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1345),
.A2(n_526),
.B1(n_531),
.B2(n_525),
.C(n_521),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1375),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1356),
.B(n_459),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1340),
.A2(n_870),
.B(n_1257),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1393),
.A2(n_1394),
.B(n_1375),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1368),
.A2(n_870),
.B(n_1184),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1368),
.A2(n_870),
.B(n_609),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1329),
.A2(n_609),
.B(n_576),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1330),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1385),
.A2(n_441),
.B1(n_448),
.B2(n_440),
.Y(n_1438)
);

AO21x2_ASAP7_75t_L g1439 ( 
.A1(n_1377),
.A2(n_467),
.B(n_460),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1329),
.A2(n_651),
.B(n_632),
.Y(n_1440)
);

CKINVDCx16_ASAP7_75t_R g1441 ( 
.A(n_1322),
.Y(n_1441)
);

OAI33xp33_ASAP7_75t_L g1442 ( 
.A1(n_1395),
.A2(n_451),
.A3(n_448),
.B1(n_461),
.B2(n_455),
.B3(n_441),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1356),
.B(n_438),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1387),
.Y(n_1444)
);

AOI22x1_ASAP7_75t_L g1445 ( 
.A1(n_1369),
.A2(n_743),
.B1(n_746),
.B2(n_464),
.Y(n_1445)
);

AO21x1_ASAP7_75t_L g1446 ( 
.A1(n_1377),
.A2(n_485),
.B(n_482),
.Y(n_1446)
);

BUFx2_ASAP7_75t_SL g1447 ( 
.A(n_1328),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1345),
.B(n_438),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1367),
.A2(n_651),
.B(n_632),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1367),
.A2(n_681),
.B(n_667),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1359),
.Y(n_1451)
);

INVx4_ASAP7_75t_L g1452 ( 
.A(n_1343),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1350),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1437),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1433),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1412),
.A2(n_1347),
.B(n_1352),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1401),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1402),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1451),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1433),
.Y(n_1460)
);

NAND2xp33_ASAP7_75t_SL g1461 ( 
.A(n_1398),
.B(n_1390),
.Y(n_1461)
);

AOI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1408),
.A2(n_1324),
.B(n_1355),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1419),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1410),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1419),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1399),
.B(n_1392),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1410),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1453),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1417),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1418),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1403),
.B(n_1361),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1418),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1424),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1444),
.Y(n_1474)
);

CKINVDCx8_ASAP7_75t_R g1475 ( 
.A(n_1447),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1415),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1453),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1424),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1423),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1430),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1427),
.Y(n_1481)
);

OAI222xp33_ASAP7_75t_L g1482 ( 
.A1(n_1425),
.A2(n_1385),
.B1(n_1336),
.B2(n_1354),
.C1(n_1386),
.C2(n_736),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1427),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1404),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1409),
.A2(n_1373),
.B1(n_1362),
.B2(n_1391),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1428),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1439),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1397),
.A2(n_1364),
.B1(n_1379),
.B2(n_1336),
.Y(n_1488)
);

INVxp67_ASAP7_75t_SL g1489 ( 
.A(n_1421),
.Y(n_1489)
);

AO21x1_ASAP7_75t_L g1490 ( 
.A1(n_1406),
.A2(n_495),
.B(n_486),
.Y(n_1490)
);

AO21x2_ASAP7_75t_L g1491 ( 
.A1(n_1432),
.A2(n_1324),
.B(n_1361),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1443),
.B(n_1387),
.Y(n_1492)
);

BUFx10_ASAP7_75t_L g1493 ( 
.A(n_1406),
.Y(n_1493)
);

AOI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1446),
.A2(n_1391),
.B(n_514),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1444),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1448),
.B(n_1361),
.Y(n_1496)
);

AOI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1415),
.A2(n_515),
.B(n_502),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1415),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1439),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1442),
.A2(n_1370),
.B1(n_1388),
.B2(n_1387),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1478),
.Y(n_1501)
);

BUFx2_ASAP7_75t_SL g1502 ( 
.A(n_1475),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1495),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1489),
.B(n_1441),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_R g1505 ( 
.A(n_1475),
.B(n_1398),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1476),
.B(n_1498),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1495),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1479),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1486),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1459),
.B(n_1431),
.Y(n_1510)
);

CKINVDCx16_ASAP7_75t_R g1511 ( 
.A(n_1486),
.Y(n_1511)
);

CKINVDCx16_ASAP7_75t_R g1512 ( 
.A(n_1461),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_SL g1513 ( 
.A(n_1462),
.B(n_1452),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1476),
.B(n_1449),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1485),
.A2(n_1400),
.B1(n_1388),
.B2(n_1363),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1478),
.Y(n_1516)
);

OA21x2_ASAP7_75t_L g1517 ( 
.A1(n_1484),
.A2(n_1499),
.B(n_1487),
.Y(n_1517)
);

NAND2xp33_ASAP7_75t_R g1518 ( 
.A(n_1466),
.B(n_1426),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1457),
.B(n_1400),
.Y(n_1519)
);

OR2x6_ASAP7_75t_L g1520 ( 
.A(n_1476),
.B(n_1449),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1458),
.Y(n_1521)
);

NAND2xp33_ASAP7_75t_R g1522 ( 
.A(n_1496),
.B(n_1450),
.Y(n_1522)
);

NOR3xp33_ASAP7_75t_SL g1523 ( 
.A(n_1482),
.B(n_455),
.C(n_451),
.Y(n_1523)
);

AO31x2_ASAP7_75t_L g1524 ( 
.A1(n_1487),
.A2(n_1452),
.A3(n_1353),
.B(n_681),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1488),
.B(n_1370),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1462),
.A2(n_1432),
.B(n_1411),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1454),
.B(n_1344),
.Y(n_1527)
);

NOR3xp33_ASAP7_75t_SL g1528 ( 
.A(n_1456),
.B(n_1488),
.C(n_465),
.Y(n_1528)
);

NAND2xp33_ASAP7_75t_R g1529 ( 
.A(n_1496),
.B(n_1450),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1500),
.A2(n_1414),
.B1(n_1354),
.B2(n_1353),
.Y(n_1530)
);

AO31x2_ASAP7_75t_L g1531 ( 
.A1(n_1499),
.A2(n_707),
.A3(n_736),
.B(n_667),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_R g1532 ( 
.A(n_1498),
.B(n_1416),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1474),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1474),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1474),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1463),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1465),
.Y(n_1537)
);

NOR3xp33_ASAP7_75t_SL g1538 ( 
.A(n_1492),
.B(n_465),
.C(n_461),
.Y(n_1538)
);

NAND2xp33_ASAP7_75t_R g1539 ( 
.A(n_1498),
.B(n_1416),
.Y(n_1539)
);

NAND2xp33_ASAP7_75t_R g1540 ( 
.A(n_1498),
.B(n_1416),
.Y(n_1540)
);

AO32x2_ASAP7_75t_L g1541 ( 
.A1(n_1493),
.A2(n_1438),
.A3(n_1339),
.B1(n_1337),
.B2(n_1342),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1480),
.B(n_1361),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1473),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1473),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1490),
.A2(n_442),
.B1(n_438),
.B2(n_1384),
.Y(n_1545)
);

NAND3xp33_ASAP7_75t_L g1546 ( 
.A(n_1519),
.B(n_1480),
.C(n_1469),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1506),
.B(n_1471),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1528),
.A2(n_1497),
.B1(n_1494),
.B2(n_1471),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1510),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1517),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1533),
.B(n_1460),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1501),
.Y(n_1552)
);

INVx5_ASAP7_75t_L g1553 ( 
.A(n_1514),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1543),
.B(n_1544),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1543),
.B(n_1470),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1507),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1517),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1501),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1504),
.B(n_1472),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1516),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1516),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1507),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1521),
.Y(n_1563)
);

INVxp67_ASAP7_75t_SL g1564 ( 
.A(n_1544),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1508),
.Y(n_1565)
);

NOR2x1_ASAP7_75t_L g1566 ( 
.A(n_1502),
.B(n_1472),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1534),
.B(n_1464),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1535),
.B(n_1460),
.Y(n_1568)
);

OR2x6_ASAP7_75t_L g1569 ( 
.A(n_1514),
.B(n_1497),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1503),
.B(n_1460),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1521),
.Y(n_1571)
);

AOI211x1_ASAP7_75t_L g1572 ( 
.A1(n_1546),
.A2(n_1490),
.B(n_1515),
.C(n_1527),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1552),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1550),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1550),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1569),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1558),
.Y(n_1577)
);

AO31x2_ASAP7_75t_L g1578 ( 
.A1(n_1557),
.A2(n_1513),
.A3(n_1484),
.B(n_1542),
.Y(n_1578)
);

AND4x1_ASAP7_75t_L g1579 ( 
.A(n_1566),
.B(n_1525),
.C(n_1523),
.D(n_1538),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1557),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1571),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1569),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1565),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1554),
.Y(n_1584)
);

NAND4xp25_ASAP7_75t_L g1585 ( 
.A(n_1548),
.B(n_1518),
.C(n_1429),
.D(n_1522),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1549),
.B(n_1537),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1553),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1560),
.A2(n_1526),
.B(n_1455),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1555),
.Y(n_1589)
);

A2O1A1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1553),
.A2(n_1545),
.B(n_1530),
.C(n_744),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1553),
.B(n_1512),
.Y(n_1591)
);

OAI21xp33_ASAP7_75t_L g1592 ( 
.A1(n_1569),
.A2(n_1505),
.B(n_476),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1554),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1555),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1553),
.Y(n_1595)
);

AOI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1559),
.A2(n_522),
.B(n_523),
.C(n_517),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1567),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1547),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1560),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1587),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1598),
.B(n_1547),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1583),
.B(n_1564),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1585),
.A2(n_1569),
.B1(n_744),
.B2(n_707),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1573),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1574),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1577),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1598),
.B(n_1553),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1594),
.B(n_1567),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1591),
.B(n_1551),
.Y(n_1609)
);

INVxp67_ASAP7_75t_SL g1610 ( 
.A(n_1574),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1581),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1575),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1589),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1587),
.B(n_1568),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1595),
.B(n_1570),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_L g1616 ( 
.A(n_1595),
.B(n_1509),
.Y(n_1616)
);

AO21x2_ASAP7_75t_L g1617 ( 
.A1(n_1575),
.A2(n_1570),
.B(n_1561),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1572),
.A2(n_552),
.B1(n_554),
.B2(n_545),
.C(n_533),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1576),
.B(n_1556),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1576),
.B(n_1556),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1588),
.A2(n_1563),
.B(n_1455),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1584),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1580),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1576),
.B(n_1556),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1592),
.A2(n_442),
.B1(n_438),
.B2(n_1445),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1576),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1580),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1619),
.B(n_1582),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1619),
.B(n_1582),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1604),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1600),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1603),
.A2(n_1596),
.B1(n_1590),
.B2(n_1529),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1620),
.B(n_1593),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1613),
.B(n_1597),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1624),
.B(n_1593),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1613),
.B(n_1599),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1624),
.B(n_1578),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1617),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1600),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1617),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1615),
.B(n_1578),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1615),
.B(n_1578),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1615),
.B(n_1578),
.Y(n_1643)
);

NOR4xp25_ASAP7_75t_SL g1644 ( 
.A(n_1618),
.B(n_1539),
.C(n_1540),
.D(n_1532),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1616),
.B(n_1599),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1600),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1609),
.B(n_1586),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1616),
.B(n_1588),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1609),
.B(n_1586),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1623),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1617),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1631),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1639),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1650),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1626),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1634),
.B(n_1608),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1628),
.B(n_1629),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1631),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1631),
.B(n_1626),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1646),
.B(n_1626),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1646),
.B(n_1606),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1646),
.B(n_1626),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1629),
.B(n_1614),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_SL g1664 ( 
.A(n_1645),
.Y(n_1664)
);

NAND2x1p5_ASAP7_75t_L g1665 ( 
.A(n_1645),
.B(n_1509),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1630),
.Y(n_1666)
);

NAND2x1p5_ASAP7_75t_L g1667 ( 
.A(n_1645),
.B(n_1579),
.Y(n_1667)
);

AOI32xp33_ASAP7_75t_L g1668 ( 
.A1(n_1647),
.A2(n_1618),
.A3(n_1607),
.B1(n_1601),
.B2(n_1625),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1634),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1636),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1636),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1647),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1633),
.B(n_1606),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1633),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1632),
.B(n_1511),
.Y(n_1675)
);

NOR2x1_ASAP7_75t_L g1676 ( 
.A(n_1645),
.B(n_1607),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1635),
.B(n_1611),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1649),
.B(n_1611),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1649),
.B(n_1622),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1638),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1653),
.Y(n_1681)
);

INVx4_ASAP7_75t_L g1682 ( 
.A(n_1660),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1660),
.B(n_1601),
.Y(n_1683)
);

NAND2x1p5_ASAP7_75t_L g1684 ( 
.A(n_1659),
.B(n_1632),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1657),
.B(n_1663),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_SL g1686 ( 
.A(n_1667),
.B(n_1590),
.Y(n_1686)
);

NAND2x1p5_ASAP7_75t_L g1687 ( 
.A(n_1662),
.B(n_1376),
.Y(n_1687)
);

AOI222xp33_ASAP7_75t_L g1688 ( 
.A1(n_1675),
.A2(n_1625),
.B1(n_717),
.B2(n_572),
.C1(n_563),
.C2(n_582),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1672),
.B(n_1608),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1654),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1656),
.B(n_1602),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1662),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1674),
.B(n_1637),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1655),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1669),
.B(n_1670),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1655),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1665),
.B(n_1637),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1652),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1671),
.B(n_1610),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1658),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1664),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1661),
.B(n_1648),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1661),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1666),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1668),
.B(n_1627),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1679),
.Y(n_1706)
);

AND2x2_ASAP7_75t_SL g1707 ( 
.A(n_1678),
.B(n_1648),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1679),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1678),
.B(n_1641),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1673),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1677),
.B(n_1641),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1680),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1653),
.B(n_1623),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1653),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1660),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1653),
.B(n_1627),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1653),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1664),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1653),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1676),
.A2(n_1612),
.B(n_1605),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1653),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_SL g1722 ( 
.A1(n_1667),
.A2(n_1642),
.B1(n_1643),
.B2(n_1648),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1653),
.Y(n_1723)
);

OAI21xp33_ASAP7_75t_L g1724 ( 
.A1(n_1675),
.A2(n_1643),
.B(n_1642),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1664),
.Y(n_1725)
);

BUFx12f_ASAP7_75t_L g1726 ( 
.A(n_1667),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1681),
.B(n_1605),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1713),
.Y(n_1728)
);

INVxp67_ASAP7_75t_L g1729 ( 
.A(n_1715),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1713),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1716),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1715),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_SL g1733 ( 
.A1(n_1684),
.A2(n_1644),
.B1(n_1638),
.B2(n_1640),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1701),
.B(n_1725),
.Y(n_1734)
);

AOI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1724),
.A2(n_1705),
.B1(n_1718),
.B2(n_1684),
.C(n_1717),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1682),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1716),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1686),
.B(n_1612),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1714),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1683),
.B(n_1640),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1719),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1683),
.B(n_1640),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1721),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1723),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1726),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1691),
.B(n_1651),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1712),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1703),
.B(n_1651),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1689),
.B(n_1706),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1690),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1708),
.B(n_1698),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1700),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1694),
.B(n_1621),
.Y(n_1753)
);

CKINVDCx16_ASAP7_75t_R g1754 ( 
.A(n_1697),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1724),
.B(n_1346),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1720),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1704),
.Y(n_1757)
);

O2A1O1Ixp33_ASAP7_75t_L g1758 ( 
.A1(n_1688),
.A2(n_570),
.B(n_584),
.C(n_557),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1699),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1693),
.B(n_1696),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1702),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1709),
.B(n_1562),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1695),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1722),
.B(n_1507),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1707),
.B(n_1563),
.Y(n_1765)
);

NOR3xp33_ASAP7_75t_L g1766 ( 
.A(n_1710),
.B(n_589),
.C(n_588),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1711),
.B(n_1621),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1687),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1722),
.B(n_1621),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1681),
.B(n_469),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1685),
.B(n_1541),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1685),
.B(n_1541),
.Y(n_1772)
);

AOI211xp5_ASAP7_75t_L g1773 ( 
.A1(n_1701),
.A2(n_477),
.B(n_478),
.C(n_476),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1692),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_SL g1775 ( 
.A(n_1681),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1732),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1735),
.A2(n_481),
.B1(n_732),
.B2(n_480),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1733),
.B(n_481),
.C(n_480),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1729),
.B(n_617),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1745),
.A2(n_1520),
.B1(n_733),
.B2(n_741),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1749),
.Y(n_1781)
);

AOI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1775),
.A2(n_637),
.B1(n_642),
.B2(n_627),
.C(n_625),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1736),
.B(n_644),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1758),
.A2(n_1755),
.B(n_1764),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1761),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1768),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1760),
.B(n_645),
.Y(n_1787)
);

OAI31xp33_ASAP7_75t_L g1788 ( 
.A1(n_1769),
.A2(n_653),
.A3(n_656),
.B(n_646),
.Y(n_1788)
);

AOI222xp33_ASAP7_75t_L g1789 ( 
.A1(n_1728),
.A2(n_1731),
.B1(n_1730),
.B2(n_1737),
.C1(n_1741),
.C2(n_1739),
.Y(n_1789)
);

INVxp67_ASAP7_75t_L g1790 ( 
.A(n_1752),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1751),
.Y(n_1791)
);

AOI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1743),
.A2(n_676),
.B1(n_682),
.B2(n_669),
.C(n_668),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1744),
.B(n_1531),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1751),
.B(n_1531),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1727),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1727),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1759),
.B(n_1346),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1740),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1748),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1773),
.B(n_685),
.Y(n_1800)
);

OAI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1756),
.A2(n_696),
.B(n_686),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1742),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1748),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1763),
.B(n_720),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1750),
.Y(n_1805)
);

OAI22xp33_ASAP7_75t_SL g1806 ( 
.A1(n_1746),
.A2(n_746),
.B1(n_748),
.B2(n_742),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1747),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1757),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1762),
.B(n_1773),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1770),
.B(n_753),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1766),
.B(n_754),
.Y(n_1811)
);

INVxp67_ASAP7_75t_L g1812 ( 
.A(n_1765),
.Y(n_1812)
);

AOI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1771),
.A2(n_538),
.B1(n_539),
.B2(n_532),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1772),
.B(n_543),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1767),
.B(n_1524),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1753),
.B(n_548),
.Y(n_1816)
);

AOI32xp33_ASAP7_75t_L g1817 ( 
.A1(n_1753),
.A2(n_560),
.A3(n_562),
.B1(n_555),
.B2(n_551),
.Y(n_1817)
);

OAI21xp33_ASAP7_75t_L g1818 ( 
.A1(n_1745),
.A2(n_1477),
.B(n_1468),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1774),
.B(n_566),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1774),
.B(n_574),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1774),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1774),
.B(n_575),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1774),
.Y(n_1823)
);

O2A1O1Ixp5_ASAP7_75t_SL g1824 ( 
.A1(n_1729),
.A2(n_578),
.B(n_579),
.C(n_577),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1774),
.Y(n_1825)
);

OAI21xp33_ASAP7_75t_SL g1826 ( 
.A1(n_1738),
.A2(n_1536),
.B(n_1348),
.Y(n_1826)
);

INVx3_ASAP7_75t_L g1827 ( 
.A(n_1732),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1774),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1734),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1754),
.B(n_1333),
.Y(n_1830)
);

OAI32xp33_ASAP7_75t_L g1831 ( 
.A1(n_1754),
.A2(n_597),
.A3(n_598),
.B1(n_596),
.B2(n_594),
.Y(n_1831)
);

AND3x1_ASAP7_75t_L g1832 ( 
.A(n_1735),
.B(n_1334),
.C(n_1455),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1734),
.B(n_0),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1774),
.B(n_599),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1754),
.B(n_1334),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1774),
.B(n_604),
.Y(n_1836)
);

AOI222xp33_ASAP7_75t_L g1837 ( 
.A1(n_1735),
.A2(n_611),
.B1(n_606),
.B2(n_612),
.C1(n_608),
.C2(n_605),
.Y(n_1837)
);

INVx1_ASAP7_75t_SL g1838 ( 
.A(n_1734),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1734),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1735),
.A2(n_615),
.B(n_613),
.Y(n_1840)
);

OAI221xp5_ASAP7_75t_SL g1841 ( 
.A1(n_1735),
.A2(n_1483),
.B1(n_1481),
.B2(n_1467),
.C(n_22),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1774),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1735),
.A2(n_623),
.B1(n_624),
.B2(n_622),
.C(n_621),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1735),
.A2(n_629),
.B(n_626),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1774),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1734),
.Y(n_1846)
);

AOI222xp33_ASAP7_75t_L g1847 ( 
.A1(n_1735),
.A2(n_641),
.B1(n_631),
.B2(n_648),
.C1(n_640),
.C2(n_630),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1734),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1734),
.B(n_2),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1774),
.B(n_654),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1735),
.A2(n_670),
.B1(n_671),
.B2(n_657),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1845),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1838),
.B(n_678),
.Y(n_1853)
);

INVx1_ASAP7_75t_SL g1854 ( 
.A(n_1839),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1835),
.B(n_680),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1829),
.B(n_683),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1846),
.B(n_1848),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1833),
.Y(n_1858)
);

INVx2_ASAP7_75t_SL g1859 ( 
.A(n_1827),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1781),
.B(n_690),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1786),
.B(n_691),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1849),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1821),
.B(n_693),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1812),
.B(n_695),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1823),
.B(n_697),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1809),
.B(n_1825),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1828),
.B(n_6),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1842),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_1832),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1777),
.A2(n_708),
.B1(n_711),
.B2(n_704),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1798),
.B(n_712),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1802),
.B(n_8),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1776),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1785),
.B(n_723),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1787),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1790),
.B(n_9),
.Y(n_1876)
);

NOR2xp67_ASAP7_75t_L g1877 ( 
.A(n_1826),
.B(n_1791),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1784),
.B(n_10),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1783),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1795),
.Y(n_1880)
);

NAND3xp33_ASAP7_75t_L g1881 ( 
.A(n_1837),
.B(n_1847),
.C(n_1843),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1796),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_SL g1883 ( 
.A(n_1841),
.B(n_1341),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1779),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1789),
.B(n_11),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1810),
.B(n_11),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1778),
.A2(n_1780),
.B1(n_1813),
.B2(n_1851),
.Y(n_1887)
);

INVx2_ASAP7_75t_SL g1888 ( 
.A(n_1830),
.Y(n_1888)
);

INVxp67_ASAP7_75t_L g1889 ( 
.A(n_1797),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1799),
.Y(n_1890)
);

NAND2x1_ASAP7_75t_L g1891 ( 
.A(n_1808),
.B(n_1341),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1818),
.B(n_16),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1803),
.B(n_16),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1793),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1794),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1814),
.B(n_1819),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1805),
.B(n_17),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1807),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1820),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1822),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1834),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1831),
.B(n_19),
.Y(n_1902)
);

NAND2xp33_ASAP7_75t_SL g1903 ( 
.A(n_1836),
.B(n_1335),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1788),
.B(n_21),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_R g1905 ( 
.A(n_1850),
.B(n_22),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1844),
.B(n_23),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1800),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1817),
.B(n_24),
.Y(n_1908)
);

NAND3xp33_ASAP7_75t_SL g1909 ( 
.A(n_1840),
.B(n_453),
.C(n_450),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1804),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1816),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1854),
.B(n_1806),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1859),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1857),
.B(n_1811),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1867),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1872),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1897),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1893),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1876),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1878),
.B(n_1801),
.Y(n_1920)
);

INVxp67_ASAP7_75t_L g1921 ( 
.A(n_1883),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1875),
.B(n_1782),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1858),
.B(n_1815),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1862),
.B(n_1792),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1869),
.B(n_1824),
.Y(n_1925)
);

CKINVDCx14_ASAP7_75t_R g1926 ( 
.A(n_1905),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1868),
.Y(n_1927)
);

NAND2xp33_ASAP7_75t_SL g1928 ( 
.A(n_1891),
.B(n_1335),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1877),
.B(n_28),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1873),
.B(n_1888),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1853),
.B(n_30),
.Y(n_1931)
);

AOI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1881),
.A2(n_692),
.B1(n_674),
.B2(n_442),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1856),
.B(n_30),
.Y(n_1933)
);

NOR3xp33_ASAP7_75t_L g1934 ( 
.A(n_1887),
.B(n_453),
.C(n_450),
.Y(n_1934)
);

NAND2xp33_ASAP7_75t_SL g1935 ( 
.A(n_1861),
.B(n_1335),
.Y(n_1935)
);

OAI21xp33_ASAP7_75t_L g1936 ( 
.A1(n_1889),
.A2(n_692),
.B(n_674),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1892),
.A2(n_692),
.B1(n_674),
.B2(n_442),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1900),
.B(n_31),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1911),
.B(n_32),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1886),
.B(n_32),
.Y(n_1940)
);

OAI21xp33_ASAP7_75t_L g1941 ( 
.A1(n_1910),
.A2(n_1483),
.B(n_692),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1860),
.B(n_33),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1908),
.B(n_35),
.Y(n_1943)
);

INVxp33_ASAP7_75t_L g1944 ( 
.A(n_1902),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1907),
.B(n_35),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1896),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1879),
.B(n_1884),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1904),
.B(n_37),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1899),
.B(n_37),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1890),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1906),
.B(n_38),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1880),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1882),
.Y(n_1953)
);

AOI221xp5_ASAP7_75t_L g1954 ( 
.A1(n_1903),
.A2(n_475),
.B1(n_479),
.B2(n_474),
.C(n_463),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1898),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1901),
.B(n_40),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1855),
.B(n_40),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1864),
.B(n_42),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1863),
.B(n_42),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1870),
.B(n_1895),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1870),
.B(n_1350),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1909),
.A2(n_1420),
.B(n_479),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1871),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1865),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1894),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1874),
.B(n_43),
.Y(n_1966)
);

OR2x2_ASAP7_75t_L g1967 ( 
.A(n_1854),
.B(n_45),
.Y(n_1967)
);

NOR2xp67_ASAP7_75t_L g1968 ( 
.A(n_1852),
.B(n_46),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1852),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1859),
.B(n_48),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1859),
.B(n_52),
.Y(n_1971)
);

OAI21xp5_ASAP7_75t_SL g1972 ( 
.A1(n_1854),
.A2(n_52),
.B(n_53),
.Y(n_1972)
);

AOI221xp5_ASAP7_75t_L g1973 ( 
.A1(n_1885),
.A2(n_729),
.B1(n_740),
.B2(n_728),
.C(n_475),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1859),
.B(n_53),
.Y(n_1974)
);

INVx2_ASAP7_75t_SL g1975 ( 
.A(n_1859),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1859),
.B(n_54),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1866),
.B(n_55),
.Y(n_1977)
);

AOI22xp33_ASAP7_75t_SL g1978 ( 
.A1(n_1854),
.A2(n_442),
.B1(n_438),
.B2(n_1389),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1852),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1852),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1859),
.B(n_57),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1859),
.B(n_59),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1852),
.Y(n_1983)
);

NAND2xp33_ASAP7_75t_L g1984 ( 
.A(n_1852),
.B(n_438),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1852),
.Y(n_1985)
);

INVxp67_ASAP7_75t_L g1986 ( 
.A(n_1852),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1917),
.B(n_60),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1968),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1926),
.B(n_61),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_L g1990 ( 
.A(n_1986),
.B(n_62),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1975),
.B(n_1981),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1981),
.B(n_63),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1944),
.B(n_64),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1968),
.Y(n_1994)
);

XNOR2xp5_ASAP7_75t_L g1995 ( 
.A(n_1912),
.B(n_64),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1969),
.B(n_67),
.Y(n_1996)
);

AOI32xp33_ASAP7_75t_L g1997 ( 
.A1(n_1913),
.A2(n_1440),
.A3(n_1436),
.B1(n_69),
.B2(n_67),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1977),
.Y(n_1998)
);

NOR3x1_ASAP7_75t_L g1999 ( 
.A(n_1972),
.B(n_69),
.C(n_70),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1930),
.B(n_1918),
.Y(n_2000)
);

AO21x1_ASAP7_75t_L g2001 ( 
.A1(n_1929),
.A2(n_74),
.B(n_76),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1967),
.Y(n_2002)
);

NOR2x1_ASAP7_75t_L g2003 ( 
.A(n_1979),
.B(n_77),
.Y(n_2003)
);

OAI21xp33_ASAP7_75t_L g2004 ( 
.A1(n_1921),
.A2(n_1467),
.B(n_618),
.Y(n_2004)
);

NOR2x1_ASAP7_75t_L g2005 ( 
.A(n_1980),
.B(n_79),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1983),
.B(n_80),
.Y(n_2006)
);

AOI211xp5_ASAP7_75t_L g2007 ( 
.A1(n_1985),
.A2(n_85),
.B(n_82),
.C(n_83),
.Y(n_2007)
);

INVx1_ASAP7_75t_SL g2008 ( 
.A(n_1939),
.Y(n_2008)
);

AOI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1984),
.A2(n_639),
.B(n_633),
.Y(n_2009)
);

NAND4xp75_ASAP7_75t_L g2010 ( 
.A(n_1925),
.B(n_92),
.C(n_87),
.D(n_88),
.Y(n_2010)
);

NOR2x1_ASAP7_75t_L g2011 ( 
.A(n_1915),
.B(n_93),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1946),
.B(n_442),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1916),
.B(n_94),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1970),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1927),
.B(n_649),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1951),
.A2(n_97),
.B(n_95),
.C(n_96),
.Y(n_2016)
);

NAND3xp33_ASAP7_75t_L g2017 ( 
.A(n_1973),
.B(n_659),
.C(n_655),
.Y(n_2017)
);

NOR2xp67_ASAP7_75t_SL g2018 ( 
.A(n_1919),
.B(n_660),
.Y(n_2018)
);

NOR3xp33_ASAP7_75t_L g2019 ( 
.A(n_1914),
.B(n_675),
.C(n_666),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1971),
.Y(n_2020)
);

NAND4xp25_ASAP7_75t_L g2021 ( 
.A(n_1922),
.B(n_102),
.C(n_99),
.D(n_100),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1974),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1976),
.B(n_103),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1982),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1949),
.Y(n_2025)
);

NAND4xp25_ASAP7_75t_L g2026 ( 
.A(n_1924),
.B(n_110),
.C(n_108),
.D(n_109),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_1965),
.Y(n_2027)
);

NAND3xp33_ASAP7_75t_SL g2028 ( 
.A(n_1960),
.B(n_1923),
.C(n_1920),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1956),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1948),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1988),
.B(n_1945),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1994),
.B(n_1938),
.Y(n_2032)
);

AOI221xp5_ASAP7_75t_L g2033 ( 
.A1(n_2028),
.A2(n_1935),
.B1(n_1952),
.B2(n_1953),
.C(n_1950),
.Y(n_2033)
);

AOI222xp33_ASAP7_75t_L g2034 ( 
.A1(n_1995),
.A2(n_1955),
.B1(n_2027),
.B2(n_2000),
.C1(n_1991),
.C2(n_2008),
.Y(n_2034)
);

BUFx6f_ASAP7_75t_L g2035 ( 
.A(n_2027),
.Y(n_2035)
);

A2O1A1Ixp33_ASAP7_75t_L g2036 ( 
.A1(n_1996),
.A2(n_1928),
.B(n_1932),
.C(n_1940),
.Y(n_2036)
);

AOI321xp33_ASAP7_75t_L g2037 ( 
.A1(n_1998),
.A2(n_1947),
.A3(n_1964),
.B1(n_1963),
.B2(n_1934),
.C(n_1961),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_2001),
.B(n_1978),
.Y(n_2038)
);

AOI221xp5_ASAP7_75t_L g2039 ( 
.A1(n_1990),
.A2(n_1941),
.B1(n_1936),
.B2(n_1962),
.C(n_1954),
.Y(n_2039)
);

OAI221xp5_ASAP7_75t_L g2040 ( 
.A1(n_2006),
.A2(n_1937),
.B1(n_1943),
.B2(n_1936),
.C(n_1931),
.Y(n_2040)
);

AND4x1_ASAP7_75t_L g2041 ( 
.A(n_1989),
.B(n_1942),
.C(n_1933),
.D(n_1966),
.Y(n_2041)
);

AOI221xp5_ASAP7_75t_L g2042 ( 
.A1(n_2004),
.A2(n_1932),
.B1(n_1958),
.B2(n_1957),
.C(n_1959),
.Y(n_2042)
);

AOI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1993),
.A2(n_1491),
.B1(n_1396),
.B2(n_1405),
.Y(n_2043)
);

AOI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_2002),
.A2(n_1491),
.B1(n_1405),
.B2(n_1422),
.Y(n_2044)
);

AOI221xp5_ASAP7_75t_L g2045 ( 
.A1(n_2025),
.A2(n_116),
.B1(n_113),
.B2(n_115),
.C(n_117),
.Y(n_2045)
);

NAND3xp33_ASAP7_75t_L g2046 ( 
.A(n_2011),
.B(n_2005),
.C(n_2003),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_2029),
.A2(n_1411),
.B1(n_1434),
.B2(n_1413),
.Y(n_2047)
);

OAI211xp5_ASAP7_75t_L g2048 ( 
.A1(n_1987),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_2048)
);

NAND4xp25_ASAP7_75t_L g2049 ( 
.A(n_1999),
.B(n_125),
.C(n_123),
.D(n_124),
.Y(n_2049)
);

AOI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_2030),
.A2(n_1434),
.B1(n_1413),
.B2(n_1407),
.Y(n_2050)
);

AOI221xp5_ASAP7_75t_L g2051 ( 
.A1(n_2014),
.A2(n_131),
.B1(n_127),
.B2(n_129),
.C(n_132),
.Y(n_2051)
);

AOI211xp5_ASAP7_75t_L g2052 ( 
.A1(n_2020),
.A2(n_131),
.B(n_127),
.C(n_129),
.Y(n_2052)
);

AOI221xp5_ASAP7_75t_L g2053 ( 
.A1(n_2022),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.C(n_136),
.Y(n_2053)
);

AOI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_2012),
.A2(n_134),
.B(n_138),
.Y(n_2054)
);

AOI221xp5_ASAP7_75t_L g2055 ( 
.A1(n_2024),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.C(n_144),
.Y(n_2055)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2056 ( 
.A1(n_2016),
.A2(n_149),
.B(n_147),
.C(n_148),
.D(n_150),
.Y(n_2056)
);

NAND4xp25_ASAP7_75t_SL g2057 ( 
.A(n_2007),
.B(n_150),
.C(n_148),
.D(n_149),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2013),
.B(n_153),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2010),
.Y(n_2059)
);

OAI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_2023),
.A2(n_1435),
.B(n_154),
.Y(n_2060)
);

NAND2xp33_ASAP7_75t_SL g2061 ( 
.A(n_2018),
.B(n_155),
.Y(n_2061)
);

NOR4xp75_ASAP7_75t_SL g2062 ( 
.A(n_1992),
.B(n_158),
.C(n_155),
.D(n_157),
.Y(n_2062)
);

AOI221xp5_ASAP7_75t_L g2063 ( 
.A1(n_2019),
.A2(n_165),
.B1(n_162),
.B2(n_163),
.C(n_166),
.Y(n_2063)
);

O2A1O1Ixp33_ASAP7_75t_L g2064 ( 
.A1(n_2056),
.A2(n_2015),
.B(n_2021),
.C(n_2026),
.Y(n_2064)
);

BUFx6f_ASAP7_75t_L g2065 ( 
.A(n_2035),
.Y(n_2065)
);

BUFx3_ASAP7_75t_L g2066 ( 
.A(n_2035),
.Y(n_2066)
);

NOR3xp33_ASAP7_75t_L g2067 ( 
.A(n_2031),
.B(n_2032),
.C(n_2046),
.Y(n_2067)
);

OAI211xp5_ASAP7_75t_L g2068 ( 
.A1(n_2034),
.A2(n_2017),
.B(n_2009),
.C(n_1997),
.Y(n_2068)
);

AOI211xp5_ASAP7_75t_L g2069 ( 
.A1(n_2033),
.A2(n_167),
.B(n_163),
.C(n_165),
.Y(n_2069)
);

OA211x2_ASAP7_75t_L g2070 ( 
.A1(n_2057),
.A2(n_2038),
.B(n_2055),
.C(n_2045),
.Y(n_2070)
);

AOI221xp5_ASAP7_75t_SL g2071 ( 
.A1(n_2036),
.A2(n_2040),
.B1(n_2059),
.B2(n_2042),
.C(n_2049),
.Y(n_2071)
);

OAI221xp5_ASAP7_75t_SL g2072 ( 
.A1(n_2037),
.A2(n_179),
.B1(n_174),
.B2(n_178),
.C(n_180),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2052),
.B(n_182),
.Y(n_2073)
);

INVx1_ASAP7_75t_SL g2074 ( 
.A(n_2061),
.Y(n_2074)
);

OA22x2_ASAP7_75t_L g2075 ( 
.A1(n_2048),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_SL g2076 ( 
.A1(n_2058),
.A2(n_187),
.B1(n_184),
.B2(n_185),
.Y(n_2076)
);

AOI211x1_ASAP7_75t_SL g2077 ( 
.A1(n_2054),
.A2(n_191),
.B(n_187),
.C(n_190),
.Y(n_2077)
);

OAI221xp5_ASAP7_75t_L g2078 ( 
.A1(n_2039),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.C(n_194),
.Y(n_2078)
);

NOR2x1_ASAP7_75t_L g2079 ( 
.A(n_2066),
.B(n_2062),
.Y(n_2079)
);

AOI221xp5_ASAP7_75t_L g2080 ( 
.A1(n_2072),
.A2(n_2063),
.B1(n_2053),
.B2(n_2051),
.C(n_2060),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2065),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2074),
.B(n_2041),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2076),
.B(n_2065),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_2064),
.A2(n_2043),
.B(n_2044),
.Y(n_2084)
);

NAND4xp75_ASAP7_75t_L g2085 ( 
.A(n_2071),
.B(n_196),
.C(n_194),
.D(n_195),
.Y(n_2085)
);

NOR3xp33_ASAP7_75t_SL g2086 ( 
.A(n_2068),
.B(n_196),
.C(n_197),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2077),
.B(n_2047),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2075),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_2067),
.A2(n_2050),
.B1(n_200),
.B2(n_198),
.Y(n_2089)
);

NAND4xp75_ASAP7_75t_L g2090 ( 
.A(n_2070),
.B(n_201),
.C(n_199),
.D(n_200),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2069),
.B(n_202),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2081),
.B(n_2088),
.Y(n_2092)
);

NOR2x1_ASAP7_75t_L g2093 ( 
.A(n_2090),
.B(n_2073),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_2085),
.B(n_2078),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2083),
.Y(n_2095)
);

BUFx12f_ASAP7_75t_L g2096 ( 
.A(n_2082),
.Y(n_2096)
);

OAI211xp5_ASAP7_75t_L g2097 ( 
.A1(n_2089),
.A2(n_2091),
.B(n_2084),
.C(n_2080),
.Y(n_2097)
);

OAI211xp5_ASAP7_75t_L g2098 ( 
.A1(n_2087),
.A2(n_207),
.B(n_204),
.C(n_206),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2079),
.B(n_208),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2086),
.B(n_210),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_2096),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2100),
.Y(n_2102)
);

NOR2x1p5_ASAP7_75t_L g2103 ( 
.A(n_2092),
.B(n_211),
.Y(n_2103)
);

BUFx2_ASAP7_75t_L g2104 ( 
.A(n_2093),
.Y(n_2104)
);

HB1xp67_ASAP7_75t_L g2105 ( 
.A(n_2099),
.Y(n_2105)
);

NOR2xp67_ASAP7_75t_L g2106 ( 
.A(n_2098),
.B(n_2097),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2094),
.B(n_211),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2095),
.B(n_215),
.Y(n_2108)
);

AOI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_2096),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2108),
.Y(n_2110)
);

AOI21xp5_ASAP7_75t_L g2111 ( 
.A1(n_2107),
.A2(n_217),
.B(n_218),
.Y(n_2111)
);

OR2x6_ASAP7_75t_L g2112 ( 
.A(n_2104),
.B(n_2106),
.Y(n_2112)
);

AOI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_2101),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2103),
.Y(n_2114)
);

OAI22x1_ASAP7_75t_L g2115 ( 
.A1(n_2109),
.A2(n_227),
.B1(n_223),
.B2(n_225),
.Y(n_2115)
);

OAI21xp5_ASAP7_75t_L g2116 ( 
.A1(n_2105),
.A2(n_228),
.B(n_230),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2102),
.B(n_231),
.Y(n_2117)
);

OAI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_2101),
.A2(n_235),
.B1(n_231),
.B2(n_232),
.Y(n_2118)
);

OAI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_2106),
.A2(n_232),
.B(n_235),
.Y(n_2119)
);

OAI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_2101),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2117),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_2115),
.Y(n_2122)
);

BUFx2_ASAP7_75t_L g2123 ( 
.A(n_2116),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2112),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2119),
.Y(n_2125)
);

INVx1_ASAP7_75t_SL g2126 ( 
.A(n_2114),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2121),
.Y(n_2127)
);

HB1xp67_ASAP7_75t_L g2128 ( 
.A(n_2122),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2123),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2125),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2126),
.Y(n_2131)
);

AOI22x1_ASAP7_75t_L g2132 ( 
.A1(n_2128),
.A2(n_2111),
.B1(n_2110),
.B2(n_2124),
.Y(n_2132)
);

AOI22xp33_ASAP7_75t_L g2133 ( 
.A1(n_2131),
.A2(n_2118),
.B1(n_2120),
.B2(n_2113),
.Y(n_2133)
);

OAI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_2129),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2127),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_2135)
);

NOR3xp33_ASAP7_75t_L g2136 ( 
.A(n_2130),
.B(n_252),
.C(n_254),
.Y(n_2136)
);

OAI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_2131),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2131),
.Y(n_2138)
);

AOI22xp5_ASAP7_75t_L g2139 ( 
.A1(n_2131),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2131),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_2138),
.Y(n_2141)
);

OAI22xp33_ASAP7_75t_L g2142 ( 
.A1(n_2140),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_2142)
);

OAI21x1_ASAP7_75t_L g2143 ( 
.A1(n_2132),
.A2(n_2133),
.B(n_2137),
.Y(n_2143)
);

OAI211xp5_ASAP7_75t_L g2144 ( 
.A1(n_2139),
.A2(n_266),
.B(n_267),
.C(n_268),
.Y(n_2144)
);

AO21x2_ASAP7_75t_L g2145 ( 
.A1(n_2136),
.A2(n_2134),
.B(n_2135),
.Y(n_2145)
);

BUFx2_ASAP7_75t_SL g2146 ( 
.A(n_2141),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2143),
.Y(n_2147)
);

AOI331xp33_ASAP7_75t_L g2148 ( 
.A1(n_2145),
.A2(n_281),
.A3(n_282),
.B1(n_283),
.B2(n_284),
.B3(n_285),
.C1(n_287),
.Y(n_2148)
);

OAI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_2147),
.A2(n_2144),
.B(n_2142),
.Y(n_2149)
);

OR2x6_ASAP7_75t_L g2150 ( 
.A(n_2148),
.B(n_853),
.Y(n_2150)
);

AOI22xp33_ASAP7_75t_SL g2151 ( 
.A1(n_2146),
.A2(n_288),
.B1(n_291),
.B2(n_293),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_L g2152 ( 
.A1(n_2146),
.A2(n_288),
.B1(n_293),
.B2(n_294),
.Y(n_2152)
);

AOI22xp33_ASAP7_75t_SL g2153 ( 
.A1(n_2146),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_2153)
);

AOI22xp33_ASAP7_75t_L g2154 ( 
.A1(n_2150),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_2150),
.A2(n_298),
.B1(n_300),
.B2(n_302),
.Y(n_2155)
);

AOI22xp33_ASAP7_75t_L g2156 ( 
.A1(n_2149),
.A2(n_300),
.B1(n_303),
.B2(n_304),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2154),
.B(n_2155),
.Y(n_2157)
);

AOI221xp5_ASAP7_75t_L g2158 ( 
.A1(n_2157),
.A2(n_2156),
.B1(n_2152),
.B2(n_2153),
.C(n_2151),
.Y(n_2158)
);

AOI211xp5_ASAP7_75t_L g2159 ( 
.A1(n_2158),
.A2(n_306),
.B(n_307),
.C(n_308),
.Y(n_2159)
);


endmodule