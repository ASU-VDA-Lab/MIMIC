module fake_netlist_6_3994_n_1829 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1829);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1829;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g183 ( 
.A(n_56),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_7),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_163),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_4),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_142),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_126),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_87),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_177),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_80),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_77),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_48),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_46),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_29),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_72),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_78),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_10),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_13),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_53),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_26),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_169),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_64),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_83),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_145),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_125),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_103),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_82),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_140),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_84),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_86),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_136),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_91),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_92),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_51),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_101),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_85),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_21),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_143),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_173),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_7),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_11),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_100),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_141),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_18),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_105),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_154),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_99),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_38),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_146),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_41),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_139),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_114),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_68),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_120),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_108),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_97),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_129),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_96),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_98),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_2),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_2),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_47),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_55),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_5),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_46),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_66),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_111),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_8),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_180),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_14),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_149),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_74),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_53),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_135),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_17),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_34),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_75),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_168),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_144),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_79),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_164),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_57),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_48),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_104),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_102),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_131),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_134),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_153),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_88),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_37),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_112),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_171),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_47),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_17),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_69),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_71),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_132),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_6),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_179),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_109),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_32),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_57),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_113),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_63),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_50),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_41),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_124),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_12),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_56),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_8),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_36),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_121),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_32),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_178),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_62),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_152),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_58),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_20),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_58),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_22),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_165),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_42),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_34),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_138),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_6),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_127),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_26),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_106),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_49),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_44),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_28),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_30),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_29),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_70),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_94),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_73),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_43),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_40),
.Y(n_327)
);

BUFx10_ASAP7_75t_L g328 ( 
.A(n_160),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_1),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_37),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_24),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_60),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_155),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_59),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_170),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_30),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_174),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_18),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_23),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_95),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_49),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_61),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_130),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_172),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_12),
.Y(n_345)
);

BUFx5_ASAP7_75t_L g346 ( 
.A(n_4),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_54),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_89),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_0),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_0),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_156),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_19),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_44),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_33),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_122),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_151),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_176),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_93),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_25),
.Y(n_359)
);

BUFx10_ASAP7_75t_L g360 ( 
.A(n_76),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_43),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_90),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_54),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_118),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_19),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_346),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g367 ( 
.A(n_203),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_346),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_199),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_208),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_346),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_194),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_352),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_346),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_240),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_346),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_255),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_346),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_243),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_346),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_251),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_251),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_333),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_185),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_222),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_251),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_251),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_194),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_274),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_185),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_198),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_251),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_233),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_225),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_233),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_259),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_259),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_297),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_195),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_294),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_290),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_187),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_294),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_297),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_183),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_198),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_218),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_229),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_209),
.Y(n_412)
);

INVxp33_ASAP7_75t_SL g413 ( 
.A(n_187),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_239),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_252),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_260),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_253),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_257),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_206),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_230),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_290),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_262),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_270),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_237),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_290),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_249),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_276),
.Y(n_427)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_254),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_196),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_324),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_209),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_271),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_264),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_287),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_265),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_272),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_303),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_291),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_223),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_224),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_279),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_298),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_228),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_299),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_308),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_228),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_282),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_314),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_319),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_210),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_320),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_295),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_327),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_329),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_331),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_336),
.Y(n_456)
);

OAI22x1_ASAP7_75t_R g457 ( 
.A1(n_369),
.A2(n_250),
.B1(n_361),
.B2(n_283),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_378),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_382),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_372),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_378),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_385),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_372),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_431),
.B(n_186),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_372),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_387),
.B(n_210),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_372),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_439),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_382),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_392),
.B(n_364),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_381),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_381),
.Y(n_472)
);

CKINVDCx8_ASAP7_75t_R g473 ( 
.A(n_443),
.Y(n_473)
);

BUFx2_ASAP7_75t_SL g474 ( 
.A(n_440),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_370),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_375),
.B(n_196),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_387),
.B(n_364),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_372),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_383),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_377),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_409),
.B(n_245),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_383),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_389),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_431),
.B(n_186),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_450),
.B(n_307),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

AO22x1_ASAP7_75t_SL g491 ( 
.A1(n_420),
.A2(n_307),
.B1(n_362),
.B2(n_266),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_386),
.Y(n_492)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_412),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_368),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_390),
.B(n_227),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_366),
.A2(n_245),
.B(n_190),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_431),
.B(n_188),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_373),
.A2(n_350),
.B1(n_354),
.B2(n_197),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_388),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_393),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_374),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_384),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_412),
.B(n_228),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_366),
.B(n_194),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_376),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_387),
.B(n_188),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_394),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_371),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_371),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_379),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_379),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_394),
.B(n_184),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_367),
.A2(n_363),
.B1(n_332),
.B2(n_359),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_386),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_399),
.B(n_200),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_399),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_410),
.A2(n_363),
.B1(n_359),
.B2(n_197),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_407),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_419),
.Y(n_521)
);

AND2x2_ASAP7_75t_SL g522 ( 
.A(n_430),
.B(n_194),
.Y(n_522)
);

INVxp33_ASAP7_75t_SL g523 ( 
.A(n_395),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_400),
.B(n_189),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_413),
.B(n_278),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_437),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_401),
.B(n_305),
.Y(n_527)
);

INVxp33_ASAP7_75t_L g528 ( 
.A(n_391),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_416),
.A2(n_342),
.B1(n_332),
.B2(n_334),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_423),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_395),
.B(n_325),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_420),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_405),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_458),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_510),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_460),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_460),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_483),
.B(n_411),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_483),
.B(n_411),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_458),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_458),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_461),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_510),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g545 ( 
.A(n_463),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_504),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_460),
.Y(n_547)
);

NAND3xp33_ASAP7_75t_L g548 ( 
.A(n_495),
.B(n_415),
.C(n_414),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_532),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_498),
.A2(n_529),
.B1(n_491),
.B2(n_483),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_470),
.B(n_414),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_510),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_460),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_461),
.Y(n_554)
);

INVx8_ASAP7_75t_L g555 ( 
.A(n_505),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_461),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_525),
.B(n_415),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_511),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_470),
.B(n_417),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_522),
.B(n_446),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_522),
.B(n_417),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_460),
.Y(n_562)
);

AND3x1_ASAP7_75t_L g563 ( 
.A(n_514),
.B(n_429),
.C(n_403),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_511),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_471),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_468),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_470),
.B(n_418),
.Y(n_567)
);

AOI21x1_ASAP7_75t_L g568 ( 
.A1(n_494),
.A2(n_216),
.B(n_213),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_471),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_514),
.A2(n_202),
.B1(n_205),
.B2(n_201),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_511),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_522),
.B(n_418),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_471),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_462),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_460),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_512),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_472),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_460),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_466),
.B(n_422),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_472),
.Y(n_580)
);

AOI21x1_ASAP7_75t_L g581 ( 
.A1(n_494),
.A2(n_219),
.B(n_217),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_472),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_465),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_517),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_512),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_517),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_466),
.B(n_422),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_518),
.B(n_427),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_517),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_465),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_512),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_509),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_517),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_517),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_517),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_494),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_474),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_502),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_491),
.B(n_474),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_465),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_463),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_502),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_502),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_498),
.A2(n_341),
.B1(n_342),
.B2(n_339),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_515),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_506),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_506),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_506),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_459),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_459),
.Y(n_611)
);

OAI21xp33_ASAP7_75t_SL g612 ( 
.A1(n_489),
.A2(n_406),
.B(n_402),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_469),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_469),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_SL g615 ( 
.A(n_528),
.B(n_433),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_481),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_481),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_505),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_484),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_523),
.B(n_433),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_484),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_490),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_493),
.B(n_435),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_504),
.B(n_435),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_490),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_493),
.B(n_436),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_465),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_499),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_493),
.B(n_436),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_466),
.B(n_477),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_499),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_500),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_509),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_466),
.B(n_441),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_529),
.B(n_421),
.C(n_404),
.Y(n_635)
);

NOR2x1p5_ASAP7_75t_L g636 ( 
.A(n_524),
.B(n_201),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_500),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_493),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_465),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_501),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_493),
.B(n_441),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_501),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_464),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_464),
.B(n_447),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_465),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_509),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_477),
.B(n_447),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_509),
.Y(n_648)
);

INVxp33_ASAP7_75t_L g649 ( 
.A(n_476),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_521),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_476),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_521),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_462),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_477),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_L g655 ( 
.A1(n_534),
.A2(n_524),
.B1(n_497),
.B2(n_488),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_509),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_530),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_465),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_477),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_488),
.B(n_452),
.C(n_425),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_492),
.B(n_380),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_475),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_513),
.B(n_194),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_521),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_492),
.B(n_380),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_521),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_SL g667 ( 
.A(n_534),
.B(n_202),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_507),
.B(n_231),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_L g669 ( 
.A(n_507),
.B(n_204),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_509),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_505),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_505),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_473),
.B(n_380),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_526),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_521),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_521),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_509),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_513),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_516),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_516),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_527),
.B(n_396),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_516),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_516),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_463),
.B(n_232),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_654),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_572),
.B(n_473),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_611),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_678),
.A2(n_496),
.B1(n_263),
.B2(n_204),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_574),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_630),
.A2(n_480),
.B(n_467),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_643),
.B(n_527),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_566),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_643),
.A2(n_480),
.B(n_467),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_551),
.B(n_559),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_655),
.B(n_546),
.Y(n_695)
);

INVxp67_ASAP7_75t_SL g696 ( 
.A(n_638),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_611),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_546),
.B(n_473),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_613),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_567),
.B(n_518),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_600),
.B(n_432),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_539),
.B(n_428),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_561),
.A2(n_280),
.B1(n_234),
.B2(n_235),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_678),
.B(n_521),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_574),
.B(n_448),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_653),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_668),
.B(n_463),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_540),
.B(n_453),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_654),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_613),
.Y(n_710)
);

AO221x1_ASAP7_75t_L g711 ( 
.A1(n_550),
.A2(n_204),
.B1(n_263),
.B2(n_340),
.C(n_226),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_600),
.B(n_457),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_550),
.A2(n_679),
.B1(n_683),
.B2(n_682),
.Y(n_713)
);

INVx8_ASAP7_75t_L g714 ( 
.A(n_598),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_557),
.B(n_549),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_659),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_659),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_549),
.B(n_533),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_679),
.B(n_478),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_548),
.B(n_189),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_549),
.B(n_533),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_680),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_682),
.B(n_478),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_615),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_616),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_683),
.B(n_478),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_681),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_680),
.B(n_479),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_644),
.A2(n_275),
.B1(n_241),
.B2(n_242),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_610),
.B(n_479),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_616),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_612),
.B(n_204),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_579),
.B(n_191),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_662),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_550),
.A2(n_496),
.B1(n_204),
.B2(n_263),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_560),
.A2(n_281),
.B1(n_246),
.B2(n_247),
.Y(n_736)
);

OAI221xp5_ASAP7_75t_L g737 ( 
.A1(n_612),
.A2(n_408),
.B1(n_442),
.B2(n_444),
.C(n_445),
.Y(n_737)
);

AO221x1_ASAP7_75t_L g738 ( 
.A1(n_550),
.A2(n_263),
.B1(n_313),
.B2(n_220),
.C(n_221),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_588),
.B(n_263),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_663),
.A2(n_496),
.B1(n_236),
.B2(n_238),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_610),
.B(n_479),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_621),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_614),
.B(n_485),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_621),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_614),
.B(n_617),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_638),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_R g747 ( 
.A(n_657),
.B(n_482),
.Y(n_747)
);

OR2x6_ASAP7_75t_SL g748 ( 
.A(n_598),
.B(n_657),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_634),
.B(n_424),
.Y(n_749)
);

AO221x1_ASAP7_75t_L g750 ( 
.A1(n_563),
.A2(n_277),
.B1(n_248),
.B2(n_256),
.C(n_258),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_555),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_617),
.B(n_485),
.Y(n_752)
);

O2A1O1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_647),
.A2(n_438),
.B(n_424),
.C(n_426),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_660),
.B(n_191),
.Y(n_754)
);

AOI221xp5_ASAP7_75t_L g755 ( 
.A1(n_570),
.A2(n_334),
.B1(n_205),
.B2(n_338),
.C(n_339),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_624),
.B(n_192),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_625),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_623),
.B(n_192),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_626),
.B(n_193),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_619),
.B(n_485),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_625),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_SL g762 ( 
.A(n_606),
.B(n_503),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_636),
.A2(n_641),
.B1(n_629),
.B2(n_681),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_619),
.B(n_486),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_622),
.B(n_486),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_622),
.B(n_193),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_628),
.B(n_486),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_628),
.B(n_207),
.Y(n_768)
);

NAND2xp33_ASAP7_75t_L g769 ( 
.A(n_663),
.B(n_268),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_646),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_631),
.B(n_640),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_663),
.A2(n_267),
.B1(n_323),
.B2(n_261),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_631),
.B(n_487),
.Y(n_773)
);

BUFx12f_ASAP7_75t_L g774 ( 
.A(n_606),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_667),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_640),
.Y(n_776)
);

INVx8_ASAP7_75t_L g777 ( 
.A(n_600),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_642),
.B(n_207),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_632),
.Y(n_779)
);

BUFx12f_ASAP7_75t_SL g780 ( 
.A(n_600),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_632),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_SL g782 ( 
.A(n_606),
.B(n_305),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_661),
.B(n_434),
.C(n_426),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_637),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_545),
.B(n_487),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_620),
.B(n_665),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_673),
.B(n_434),
.C(n_438),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_637),
.B(n_570),
.Y(n_788)
);

AO22x1_ASAP7_75t_L g789 ( 
.A1(n_635),
.A2(n_349),
.B1(n_338),
.B2(n_341),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_602),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_597),
.Y(n_791)
);

INVxp33_ASAP7_75t_L g792 ( 
.A(n_651),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_618),
.B(n_244),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_537),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_684),
.B(n_211),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_646),
.B(n_505),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_599),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_603),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_636),
.B(n_449),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_606),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_L g801 ( 
.A(n_674),
.B(n_605),
.C(n_454),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_648),
.B(n_505),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_648),
.B(n_505),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_618),
.B(n_212),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_656),
.B(n_505),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_656),
.B(n_505),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_L g807 ( 
.A(n_663),
.B(n_269),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_670),
.B(n_520),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_674),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_670),
.B(n_677),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_603),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_589),
.B(n_451),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_618),
.B(n_214),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_618),
.B(n_215),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_535),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_541),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_536),
.B(n_520),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_663),
.A2(n_284),
.B1(n_273),
.B2(n_304),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_589),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_541),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_669),
.A2(n_285),
.B1(n_286),
.B2(n_288),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_542),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_542),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_649),
.B(n_451),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_663),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_604),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_543),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_555),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_SL g829 ( 
.A(n_555),
.B(n_305),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_608),
.B(n_454),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_618),
.B(n_215),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_536),
.B(n_335),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_604),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_663),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_671),
.B(n_335),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_543),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_607),
.Y(n_837)
);

NAND2xp33_ASAP7_75t_SL g838 ( 
.A(n_538),
.B(n_345),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_607),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_544),
.B(n_337),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_544),
.B(n_337),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_554),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_687),
.Y(n_843)
);

BUFx8_ASAP7_75t_L g844 ( 
.A(n_734),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_687),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_694),
.A2(n_700),
.B1(n_763),
.B2(n_759),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_716),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_704),
.A2(n_555),
.B(n_593),
.Y(n_848)
);

INVx5_ASAP7_75t_L g849 ( 
.A(n_751),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_694),
.B(n_552),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_716),
.Y(n_851)
);

NOR2x2_ASAP7_75t_L g852 ( 
.A(n_712),
.B(n_457),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_697),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_735),
.B(n_558),
.Y(n_854)
);

INVx5_ASAP7_75t_L g855 ( 
.A(n_751),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_697),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_711),
.A2(n_738),
.B1(n_788),
.B2(n_735),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_745),
.B(n_558),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_689),
.B(n_455),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_771),
.B(n_564),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_699),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_824),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_702),
.B(n_564),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_692),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_702),
.B(n_571),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_788),
.A2(n_609),
.B1(n_576),
.B2(n_592),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_751),
.B(n_671),
.Y(n_867)
);

NOR3xp33_ASAP7_75t_SL g868 ( 
.A(n_755),
.B(n_349),
.C(n_347),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_699),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_716),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_710),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_774),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_688),
.A2(n_555),
.B(n_593),
.Y(n_873)
);

AND2x2_ASAP7_75t_SL g874 ( 
.A(n_782),
.B(n_455),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_716),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_747),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_747),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_710),
.Y(n_878)
);

O2A1O1Ixp5_ASAP7_75t_L g879 ( 
.A1(n_695),
.A2(n_568),
.B(n_581),
.C(n_608),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_715),
.B(n_593),
.Y(n_880)
);

NAND2x1p5_ASAP7_75t_L g881 ( 
.A(n_751),
.B(n_671),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_746),
.Y(n_882)
);

NOR2xp67_ASAP7_75t_L g883 ( 
.A(n_800),
.B(n_774),
.Y(n_883)
);

INVx5_ASAP7_75t_L g884 ( 
.A(n_828),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_725),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_727),
.B(n_671),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_725),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_731),
.Y(n_888)
);

OR2x6_ASAP7_75t_L g889 ( 
.A(n_777),
.B(n_456),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_706),
.B(n_708),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_731),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_742),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_776),
.B(n_571),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_722),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_742),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_691),
.B(n_576),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_722),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_828),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_691),
.B(n_586),
.Y(n_899)
);

OR2x6_ASAP7_75t_SL g900 ( 
.A(n_749),
.B(n_353),
.Y(n_900)
);

O2A1O1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_695),
.A2(n_732),
.B(n_737),
.C(n_713),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_718),
.B(n_671),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_705),
.B(n_456),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_744),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_799),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_746),
.B(n_531),
.Y(n_906)
);

OAI22xp33_ASAP7_75t_L g907 ( 
.A1(n_829),
.A2(n_343),
.B1(n_351),
.B2(n_344),
.Y(n_907)
);

AND2x2_ASAP7_75t_SL g908 ( 
.A(n_762),
.B(n_397),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_790),
.B(n_586),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_721),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_757),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_713),
.A2(n_609),
.B1(n_592),
.B2(n_556),
.Y(n_912)
);

INVx5_ASAP7_75t_L g913 ( 
.A(n_794),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_795),
.A2(n_676),
.B1(n_675),
.B2(n_650),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_757),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_799),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_812),
.B(n_397),
.Y(n_917)
);

AO22x1_ASAP7_75t_L g918 ( 
.A1(n_754),
.A2(n_353),
.B1(n_300),
.B2(n_302),
.Y(n_918)
);

NOR2x2_ASAP7_75t_L g919 ( 
.A(n_712),
.B(n_310),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_714),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_688),
.B(n_554),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_761),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_685),
.B(n_650),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_786),
.B(n_672),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_792),
.B(n_633),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_830),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_756),
.B(n_398),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_761),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_781),
.B(n_556),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_781),
.B(n_565),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_756),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_779),
.Y(n_932)
);

AND2x6_ASAP7_75t_L g933 ( 
.A(n_709),
.B(n_652),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_794),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_754),
.B(n_306),
.Y(n_935)
);

INVx5_ASAP7_75t_L g936 ( 
.A(n_777),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_784),
.B(n_565),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_795),
.B(n_672),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_717),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_740),
.A2(n_775),
.B1(n_724),
.B2(n_701),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_801),
.B(n_686),
.Y(n_941)
);

AND2x6_ASAP7_75t_L g942 ( 
.A(n_796),
.B(n_652),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_766),
.B(n_672),
.Y(n_943)
);

AO22x1_ASAP7_75t_L g944 ( 
.A1(n_787),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_791),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_766),
.B(n_672),
.Y(n_946)
);

AND3x1_ASAP7_75t_SL g947 ( 
.A(n_789),
.B(n_326),
.C(n_316),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_714),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_780),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_732),
.A2(n_580),
.B(n_582),
.C(n_577),
.Y(n_950)
);

CKINVDCx8_ASAP7_75t_R g951 ( 
.A(n_714),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_797),
.B(n_569),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_739),
.A2(n_676),
.B1(n_675),
.B2(n_666),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_798),
.B(n_569),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_811),
.B(n_573),
.Y(n_955)
);

AND3x1_ASAP7_75t_L g956 ( 
.A(n_783),
.B(n_519),
.C(n_508),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_826),
.B(n_573),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_698),
.B(n_318),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_750),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_809),
.B(n_321),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_833),
.B(n_837),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_777),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_839),
.B(n_577),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_730),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_701),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_741),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_SL g967 ( 
.A(n_720),
.B(n_348),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_L g968 ( 
.A(n_740),
.B(n_672),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_815),
.B(n_580),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_R g970 ( 
.A(n_838),
.B(n_348),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_733),
.B(n_633),
.Y(n_971)
);

BUFx4f_ASAP7_75t_L g972 ( 
.A(n_701),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_816),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_819),
.B(n_322),
.Y(n_974)
);

INVx6_ASAP7_75t_L g975 ( 
.A(n_712),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_748),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_758),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_SL g978 ( 
.A1(n_729),
.A2(n_330),
.B1(n_355),
.B2(n_351),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_768),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_696),
.B(n_664),
.Y(n_980)
);

BUFx5_ASAP7_75t_L g981 ( 
.A(n_802),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_739),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_SL g983 ( 
.A1(n_768),
.A2(n_310),
.B1(n_360),
.B2(n_328),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_820),
.Y(n_984)
);

XNOR2xp5_ASAP7_75t_L g985 ( 
.A(n_736),
.B(n_355),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_778),
.B(n_672),
.Y(n_986)
);

OR2x6_ASAP7_75t_L g987 ( 
.A(n_753),
.B(n_825),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_719),
.A2(n_582),
.B1(n_666),
.B2(n_664),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_822),
.B(n_583),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_778),
.B(n_633),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_832),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_772),
.A2(n_358),
.B1(n_357),
.B2(n_356),
.Y(n_992)
);

CKINVDCx16_ASAP7_75t_R g993 ( 
.A(n_703),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_832),
.B(n_310),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_728),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_743),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_840),
.B(n_841),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_841),
.B(n_357),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_810),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_752),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_760),
.Y(n_1001)
);

CKINVDCx6p67_ASAP7_75t_R g1002 ( 
.A(n_804),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_822),
.B(n_583),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_823),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_723),
.A2(n_585),
.B1(n_587),
.B2(n_590),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_770),
.B(n_585),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_823),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_764),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_834),
.B(n_726),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_707),
.B(n_358),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_SL g1011 ( 
.A1(n_769),
.A2(n_360),
.B1(n_328),
.B2(n_293),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_765),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_803),
.A2(n_587),
.B(n_590),
.C(n_594),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_827),
.B(n_594),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_767),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_827),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_773),
.B(n_595),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_836),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_931),
.B(n_785),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_846),
.B(n_821),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_997),
.B(n_836),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_897),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_979),
.B(n_693),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_864),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_R g1025 ( 
.A(n_876),
.B(n_807),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_991),
.B(n_842),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_996),
.B(n_842),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_873),
.A2(n_690),
.B(n_805),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_SL g1029 ( 
.A1(n_874),
.A2(n_328),
.B1(n_360),
.B2(n_301),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_SL g1030 ( 
.A1(n_998),
.A2(n_595),
.B(n_596),
.C(n_772),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_850),
.B(n_817),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_850),
.B(n_808),
.Y(n_1032)
);

NAND2x1p5_ASAP7_75t_L g1033 ( 
.A(n_936),
.B(n_793),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_SL g1034 ( 
.A1(n_908),
.A2(n_296),
.B1(n_292),
.B2(n_289),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_945),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_862),
.B(n_903),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_910),
.B(n_818),
.Y(n_1037)
);

CKINVDCx6p67_ASAP7_75t_R g1038 ( 
.A(n_872),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_854),
.A2(n_818),
.B1(n_806),
.B2(n_793),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_854),
.A2(n_835),
.B1(n_831),
.B2(n_814),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_901),
.A2(n_813),
.B(n_596),
.C(n_562),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_996),
.B(n_537),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_926),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_847),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1001),
.B(n_537),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_873),
.A2(n_968),
.B(n_855),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_890),
.B(n_547),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_845),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_941),
.B(n_315),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_853),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_857),
.A2(n_901),
.B1(n_993),
.B2(n_983),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1008),
.B(n_547),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_844),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_847),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_844),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_849),
.A2(n_855),
.B(n_848),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_935),
.A2(n_658),
.B(n_553),
.C(n_639),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_879),
.A2(n_1013),
.B(n_921),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_977),
.B(n_317),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_973),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_849),
.A2(n_538),
.B(n_645),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_SL g1062 ( 
.A(n_983),
.B(n_1),
.C(n_3),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_856),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_949),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_962),
.B(n_553),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_917),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_859),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_847),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_861),
.Y(n_1069)
);

AO22x1_ASAP7_75t_L g1070 ( 
.A1(n_994),
.A2(n_3),
.B1(n_5),
.B2(n_9),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_918),
.B(n_581),
.C(n_658),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_940),
.B(n_645),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_863),
.B(n_578),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_974),
.B(n_584),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_984),
.Y(n_1075)
);

AO32x2_ASAP7_75t_L g1076 ( 
.A1(n_940),
.A2(n_9),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_897),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_SL g1078 ( 
.A1(n_961),
.A2(n_115),
.B(n_181),
.Y(n_1078)
);

BUFx4f_ASAP7_75t_L g1079 ( 
.A(n_962),
.Y(n_1079)
);

AO32x2_ASAP7_75t_L g1080 ( 
.A1(n_959),
.A2(n_15),
.A3(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_927),
.B(n_578),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_985),
.B(n_575),
.Y(n_1082)
);

AOI33xp33_ASAP7_75t_L g1083 ( 
.A1(n_958),
.A2(n_22),
.A3(n_23),
.B1(n_24),
.B2(n_27),
.B3(n_28),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_SL g1084 ( 
.A1(n_990),
.A2(n_645),
.B(n_627),
.C(n_601),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_863),
.A2(n_645),
.B1(n_627),
.B2(n_601),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_865),
.B(n_645),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_960),
.B(n_27),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_849),
.A2(n_627),
.B(n_601),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_869),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_851),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_877),
.B(n_627),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_905),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_849),
.A2(n_627),
.B(n_601),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_865),
.B(n_591),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_851),
.Y(n_1095)
);

BUFx8_ASAP7_75t_SL g1096 ( 
.A(n_965),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_885),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_851),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_855),
.A2(n_591),
.B(n_538),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_925),
.B(n_880),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_879),
.A2(n_591),
.B(n_538),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_907),
.A2(n_31),
.B(n_33),
.C(n_35),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_R g1103 ( 
.A(n_951),
.B(n_119),
.Y(n_1103)
);

BUFx12f_ASAP7_75t_L g1104 ( 
.A(n_975),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_962),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_889),
.Y(n_1106)
);

INVx3_ASAP7_75t_SL g1107 ( 
.A(n_852),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_992),
.A2(n_31),
.B(n_35),
.C(n_36),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_SL g1109 ( 
.A(n_970),
.B(n_38),
.C(n_39),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_999),
.B(n_39),
.Y(n_1110)
);

OAI21xp33_ASAP7_75t_SL g1111 ( 
.A1(n_921),
.A2(n_40),
.B(n_42),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_964),
.B(n_45),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_950),
.A2(n_137),
.B(n_175),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1010),
.A2(n_480),
.B(n_467),
.C(n_51),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_SL g1115 ( 
.A1(n_972),
.A2(n_975),
.B1(n_978),
.B2(n_916),
.Y(n_1115)
);

AO32x2_ASAP7_75t_L g1116 ( 
.A1(n_982),
.A2(n_45),
.A3(n_50),
.B1(n_52),
.B2(n_59),
.Y(n_1116)
);

NOR3xp33_ASAP7_75t_L g1117 ( 
.A(n_967),
.B(n_52),
.C(n_60),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_906),
.B(n_889),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_975),
.Y(n_1119)
);

BUFx12f_ASAP7_75t_L g1120 ( 
.A(n_948),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_887),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_950),
.A2(n_148),
.B(n_65),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_868),
.B(n_61),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_SL g1124 ( 
.A(n_1011),
.B(n_67),
.C(n_81),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_920),
.B(n_900),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1004),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_966),
.B(n_107),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1012),
.B(n_116),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1015),
.B(n_128),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_888),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_992),
.A2(n_133),
.B(n_147),
.C(n_150),
.Y(n_1131)
);

INVx4_ASAP7_75t_L g1132 ( 
.A(n_936),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_936),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_939),
.B(n_157),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_896),
.B(n_161),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_939),
.B(n_162),
.Y(n_1136)
);

NOR3xp33_ASAP7_75t_SL g1137 ( 
.A(n_919),
.B(n_166),
.C(n_467),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_947),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_936),
.B(n_882),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_889),
.B(n_467),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_882),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_848),
.A2(n_480),
.B(n_858),
.Y(n_1142)
);

BUFx4f_ASAP7_75t_L g1143 ( 
.A(n_1002),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_870),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_891),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_961),
.A2(n_480),
.B(n_899),
.C(n_932),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_989),
.A2(n_1014),
.B(n_1003),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_972),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_898),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_944),
.B(n_899),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_938),
.A2(n_943),
.B(n_986),
.C(n_946),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_860),
.B(n_995),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_883),
.B(n_875),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_989),
.A2(n_1014),
.B(n_1003),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_971),
.A2(n_1009),
.B(n_893),
.C(n_909),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_SL g1156 ( 
.A1(n_870),
.A2(n_875),
.B(n_866),
.C(n_934),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_898),
.B(n_884),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1035),
.Y(n_1158)
);

NOR4xp25_ASAP7_75t_L g1159 ( 
.A(n_1062),
.B(n_893),
.C(n_909),
.D(n_924),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1046),
.A2(n_884),
.B(n_867),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1119),
.B(n_1009),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1067),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_1024),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1048),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1066),
.B(n_1067),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1096),
.Y(n_1166)
);

NAND3xp33_ASAP7_75t_SL g1167 ( 
.A(n_1029),
.B(n_914),
.C(n_902),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1079),
.Y(n_1168)
);

NAND2xp33_ASAP7_75t_R g1169 ( 
.A(n_1025),
.B(n_987),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1050),
.Y(n_1170)
);

BUFx24_ASAP7_75t_L g1171 ( 
.A(n_1157),
.Y(n_1171)
);

AOI211x1_ASAP7_75t_L g1172 ( 
.A1(n_1051),
.A2(n_1070),
.B(n_1123),
.C(n_1112),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1152),
.B(n_1000),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1021),
.B(n_1019),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_SL g1175 ( 
.A1(n_1078),
.A2(n_963),
.B(n_957),
.Y(n_1175)
);

BUFx10_ASAP7_75t_L g1176 ( 
.A(n_1125),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_1036),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1104),
.Y(n_1178)
);

INVx4_ASAP7_75t_L g1179 ( 
.A(n_1079),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1051),
.A2(n_894),
.B(n_995),
.C(n_1000),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1063),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1069),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1066),
.A2(n_912),
.B1(n_1006),
.B2(n_987),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1100),
.B(n_995),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1027),
.B(n_1006),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1142),
.A2(n_954),
.A3(n_963),
.B(n_957),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1101),
.A2(n_930),
.B(n_929),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1026),
.B(n_904),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1031),
.B(n_922),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_1105),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1028),
.A2(n_867),
.B(n_881),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1082),
.B(n_913),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1043),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1020),
.A2(n_1058),
.B(n_1041),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1057),
.A2(n_955),
.A3(n_954),
.B(n_952),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1147),
.A2(n_929),
.B(n_930),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1032),
.A2(n_913),
.B(n_955),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1064),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1118),
.B(n_976),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1132),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1150),
.B(n_843),
.Y(n_1201)
);

NOR2x1_ASAP7_75t_L g1202 ( 
.A(n_1149),
.B(n_987),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1032),
.A2(n_913),
.B1(n_952),
.B2(n_956),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_L g1204 ( 
.A(n_1117),
.B(n_923),
.C(n_1005),
.Y(n_1204)
);

BUFx10_ASAP7_75t_L g1205 ( 
.A(n_1153),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1047),
.B(n_871),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1056),
.A2(n_969),
.B(n_937),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1074),
.B(n_878),
.Y(n_1208)
);

OA22x2_ASAP7_75t_L g1209 ( 
.A1(n_1113),
.A2(n_980),
.B1(n_1018),
.B2(n_953),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_L g1210 ( 
.A(n_1102),
.B(n_988),
.C(n_892),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1154),
.A2(n_928),
.B(n_895),
.Y(n_1211)
);

AO32x2_ASAP7_75t_L g1212 ( 
.A1(n_1040),
.A2(n_1085),
.A3(n_1039),
.B1(n_1076),
.B2(n_1116),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1122),
.A2(n_980),
.B1(n_911),
.B2(n_915),
.Y(n_1213)
);

INVxp33_ASAP7_75t_L g1214 ( 
.A(n_1087),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1148),
.B(n_1007),
.Y(n_1215)
);

AOI221xp5_ASAP7_75t_L g1216 ( 
.A1(n_1108),
.A2(n_1017),
.B1(n_1016),
.B2(n_886),
.C(n_981),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1154),
.A2(n_1151),
.B(n_1085),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1122),
.A2(n_1017),
.B(n_933),
.C(n_942),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1061),
.A2(n_1093),
.B(n_1088),
.Y(n_1219)
);

AO21x1_ASAP7_75t_L g1220 ( 
.A1(n_1072),
.A2(n_933),
.B(n_942),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1099),
.A2(n_981),
.B(n_942),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1094),
.A2(n_942),
.B(n_981),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1106),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1110),
.B(n_981),
.Y(n_1224)
);

O2A1O1Ixp5_ASAP7_75t_L g1225 ( 
.A1(n_1049),
.A2(n_933),
.B(n_981),
.C(n_1023),
.Y(n_1225)
);

AOI221xp5_ASAP7_75t_L g1226 ( 
.A1(n_1109),
.A2(n_933),
.B1(n_1111),
.B2(n_1124),
.C(n_1114),
.Y(n_1226)
);

NOR2xp67_ASAP7_75t_SL g1227 ( 
.A(n_1120),
.B(n_1132),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1133),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1040),
.A2(n_1039),
.A3(n_1094),
.B(n_1086),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1105),
.Y(n_1230)
);

CKINVDCx8_ASAP7_75t_R g1231 ( 
.A(n_1053),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1073),
.B(n_1081),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1135),
.A2(n_1146),
.B(n_1071),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1089),
.B(n_1097),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1127),
.A2(n_1129),
.B(n_1128),
.C(n_1131),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1121),
.B(n_1130),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1059),
.B(n_1092),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1145),
.Y(n_1238)
);

AO21x1_ASAP7_75t_L g1239 ( 
.A1(n_1134),
.A2(n_1136),
.B(n_1037),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1042),
.B(n_1052),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1084),
.A2(n_1156),
.B(n_1030),
.Y(n_1241)
);

NAND2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1133),
.B(n_1157),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1022),
.A2(n_1077),
.B(n_1139),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1060),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1045),
.B(n_1075),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1033),
.A2(n_1022),
.B(n_1077),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1044),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1126),
.A2(n_1091),
.A3(n_1076),
.B(n_1116),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1034),
.B(n_1083),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1115),
.B(n_1141),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1141),
.B(n_1149),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1138),
.A2(n_1107),
.B1(n_1143),
.B2(n_1153),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1090),
.B(n_1105),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1065),
.B(n_1144),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1140),
.A2(n_1144),
.B(n_1044),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1038),
.Y(n_1256)
);

CKINVDCx11_ASAP7_75t_R g1257 ( 
.A(n_1055),
.Y(n_1257)
);

NOR3xp33_ASAP7_75t_L g1258 ( 
.A(n_1137),
.B(n_1143),
.C(n_1103),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1044),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1140),
.A2(n_1076),
.B(n_1116),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1098),
.B(n_1054),
.Y(n_1261)
);

NAND2x1p5_ASAP7_75t_L g1262 ( 
.A(n_1054),
.B(n_1068),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1054),
.Y(n_1263)
);

INVx3_ASAP7_75t_SL g1264 ( 
.A(n_1068),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1095),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1095),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1098),
.A2(n_846),
.B1(n_997),
.B2(n_735),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1098),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1080),
.A2(n_1046),
.B(n_873),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1080),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1080),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_SL g1272 ( 
.A1(n_1078),
.A2(n_901),
.B(n_1113),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1051),
.A2(n_997),
.B(n_846),
.C(n_998),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1155),
.A2(n_997),
.B(n_846),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1019),
.B(n_997),
.Y(n_1275)
);

OA21x2_ASAP7_75t_L g1276 ( 
.A1(n_1058),
.A2(n_1122),
.B(n_1113),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1066),
.B(n_931),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1051),
.A2(n_997),
.B(n_846),
.C(n_998),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_1067),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_1043),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1051),
.A2(n_997),
.B1(n_369),
.B2(n_375),
.Y(n_1281)
);

AOI221xp5_ASAP7_75t_L g1282 ( 
.A1(n_1051),
.A2(n_700),
.B1(n_557),
.B2(n_755),
.C(n_997),
.Y(n_1282)
);

INVxp67_ASAP7_75t_SL g1283 ( 
.A(n_1152),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1024),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1019),
.B(n_997),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1119),
.B(n_962),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1132),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1043),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1051),
.A2(n_997),
.B1(n_369),
.B2(n_375),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1051),
.A2(n_997),
.B1(n_369),
.B2(n_375),
.Y(n_1290)
);

CKINVDCx16_ASAP7_75t_R g1291 ( 
.A(n_1024),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_1024),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1101),
.A2(n_1028),
.B(n_1147),
.Y(n_1293)
);

OAI22x1_ASAP7_75t_L g1294 ( 
.A1(n_1049),
.A2(n_846),
.B1(n_985),
.B2(n_589),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1024),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1036),
.B(n_1066),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1273),
.A2(n_1278),
.B(n_1282),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1274),
.A2(n_1285),
.B1(n_1275),
.B2(n_1290),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1296),
.B(n_1177),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1284),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1241),
.A2(n_1269),
.A3(n_1239),
.B(n_1218),
.Y(n_1301)
);

INVx3_ASAP7_75t_L g1302 ( 
.A(n_1179),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1293),
.A2(n_1207),
.B(n_1191),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1292),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1179),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1198),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1221),
.A2(n_1219),
.B(n_1196),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1257),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1166),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1281),
.B(n_1289),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1274),
.A2(n_1235),
.B(n_1225),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1249),
.A2(n_1294),
.B1(n_1276),
.B2(n_1194),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1233),
.A2(n_1194),
.B(n_1217),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1158),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1187),
.A2(n_1211),
.B(n_1160),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1276),
.A2(n_1267),
.B1(n_1174),
.B2(n_1209),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1258),
.A2(n_1169),
.B1(n_1237),
.B2(n_1252),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1174),
.A2(n_1209),
.B1(n_1226),
.B2(n_1167),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1173),
.B(n_1202),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1177),
.B(n_1215),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1162),
.B(n_1279),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1197),
.A2(n_1175),
.B(n_1246),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1220),
.A2(n_1203),
.A3(n_1213),
.B(n_1271),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1203),
.A2(n_1213),
.A3(n_1270),
.B(n_1180),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1247),
.B(n_1200),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1283),
.B(n_1184),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1173),
.B(n_1254),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1232),
.A2(n_1192),
.B(n_1222),
.Y(n_1328)
);

OAI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1260),
.A2(n_1214),
.B1(n_1279),
.B2(n_1162),
.Y(n_1329)
);

OR2x6_ASAP7_75t_L g1330 ( 
.A(n_1172),
.B(n_1224),
.Y(n_1330)
);

OAI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1250),
.A2(n_1201),
.B1(n_1183),
.B2(n_1234),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1243),
.A2(n_1232),
.B(n_1240),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1183),
.A2(n_1189),
.B(n_1204),
.C(n_1210),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1165),
.A2(n_1204),
.B1(n_1210),
.B2(n_1277),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1199),
.A2(n_1223),
.B(n_1161),
.Y(n_1335)
);

AOI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1206),
.A2(n_1208),
.B(n_1245),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1185),
.B(n_1188),
.Y(n_1337)
);

INVx3_ASAP7_75t_SL g1338 ( 
.A(n_1295),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1234),
.B(n_1236),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1236),
.Y(n_1340)
);

AOI221xp5_ASAP7_75t_L g1341 ( 
.A1(n_1159),
.A2(n_1280),
.B1(n_1193),
.B2(n_1288),
.C(n_1170),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1245),
.B(n_1244),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1255),
.A2(n_1216),
.B(n_1287),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1164),
.A2(n_1238),
.B1(n_1182),
.B2(n_1181),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1263),
.Y(n_1345)
);

NAND2x1p5_ASAP7_75t_L g1346 ( 
.A(n_1247),
.B(n_1228),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1264),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1291),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1251),
.B(n_1287),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1186),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1265),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1242),
.A2(n_1261),
.B(n_1262),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1163),
.B(n_1253),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_SL g1354 ( 
.A(n_1231),
.B(n_1178),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1286),
.A2(n_1227),
.B(n_1259),
.Y(n_1355)
);

NAND2x1p5_ASAP7_75t_L g1356 ( 
.A(n_1247),
.B(n_1190),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1186),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1176),
.B(n_1268),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1266),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1186),
.Y(n_1360)
);

AO31x2_ASAP7_75t_L g1361 ( 
.A1(n_1212),
.A2(n_1229),
.A3(n_1195),
.B(n_1248),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1256),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1286),
.A2(n_1171),
.B1(n_1190),
.B2(n_1230),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1205),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1195),
.A2(n_1229),
.B(n_1212),
.Y(n_1365)
);

INVx8_ASAP7_75t_L g1366 ( 
.A(n_1230),
.Y(n_1366)
);

NOR2xp67_ASAP7_75t_L g1367 ( 
.A(n_1280),
.B(n_692),
.Y(n_1367)
);

AO21x1_ASAP7_75t_L g1368 ( 
.A1(n_1274),
.A2(n_1051),
.B(n_997),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1233),
.A2(n_1241),
.B(n_1272),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1211),
.Y(n_1370)
);

INVx6_ASAP7_75t_L g1371 ( 
.A(n_1168),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1173),
.B(n_1202),
.Y(n_1372)
);

AO21x2_ASAP7_75t_L g1373 ( 
.A1(n_1233),
.A2(n_1241),
.B(n_1272),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_1193),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1193),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1282),
.A2(n_1273),
.B(n_1278),
.C(n_997),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1275),
.B(n_1285),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1162),
.Y(n_1378)
);

AND2x6_ASAP7_75t_L g1379 ( 
.A(n_1202),
.B(n_1224),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1198),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1211),
.Y(n_1381)
);

A2O1A1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1282),
.A2(n_1273),
.B(n_1278),
.C(n_997),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1168),
.Y(n_1383)
);

AO31x2_ASAP7_75t_L g1384 ( 
.A1(n_1241),
.A2(n_1269),
.A3(n_1239),
.B(n_1218),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_SL g1385 ( 
.A1(n_1233),
.A2(n_997),
.B(n_1274),
.C(n_998),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1282),
.A2(n_1289),
.B1(n_1290),
.B2(n_1281),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1179),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1284),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1273),
.A2(n_997),
.B(n_1278),
.Y(n_1389)
);

AO32x2_ASAP7_75t_L g1390 ( 
.A1(n_1267),
.A2(n_1051),
.A3(n_1212),
.B1(n_1203),
.B2(n_1183),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1198),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1292),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1233),
.A2(n_1269),
.B(n_1241),
.Y(n_1393)
);

NAND2x1p5_ASAP7_75t_L g1394 ( 
.A(n_1202),
.B(n_1132),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1202),
.B(n_1132),
.Y(n_1395)
);

O2A1O1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1273),
.A2(n_1278),
.B(n_1282),
.C(n_1051),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1173),
.B(n_1202),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1282),
.A2(n_1062),
.B1(n_983),
.B2(n_997),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1282),
.A2(n_1275),
.B1(n_1285),
.B2(n_1278),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1211),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1158),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1198),
.Y(n_1402)
);

INVx3_ASAP7_75t_SL g1403 ( 
.A(n_1284),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1233),
.A2(n_1241),
.B(n_1272),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1158),
.Y(n_1405)
);

AO21x2_ASAP7_75t_L g1406 ( 
.A1(n_1233),
.A2(n_1241),
.B(n_1272),
.Y(n_1406)
);

NOR2xp67_ASAP7_75t_L g1407 ( 
.A(n_1280),
.B(n_692),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1179),
.Y(n_1408)
);

A2O1A1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1282),
.A2(n_1273),
.B(n_1278),
.C(n_997),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1162),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1233),
.A2(n_1269),
.B(n_1241),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1211),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_SL g1413 ( 
.A1(n_1220),
.A2(n_1078),
.B(n_1175),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1158),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1233),
.A2(n_1269),
.B(n_1241),
.Y(n_1415)
);

OR2x6_ASAP7_75t_L g1416 ( 
.A(n_1202),
.B(n_1046),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1385),
.A2(n_1389),
.B(n_1382),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1321),
.Y(n_1418)
);

O2A1O1Ixp5_ASAP7_75t_L g1419 ( 
.A1(n_1297),
.A2(n_1368),
.B(n_1385),
.C(n_1382),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1376),
.A2(n_1409),
.B(n_1311),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1299),
.B(n_1326),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1309),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1376),
.A2(n_1409),
.B(n_1396),
.Y(n_1423)
);

AOI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1398),
.A2(n_1396),
.B1(n_1399),
.B2(n_1310),
.C(n_1386),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1298),
.B(n_1377),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1327),
.B(n_1378),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1298),
.B(n_1339),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1319),
.B(n_1372),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1337),
.B(n_1340),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1310),
.B(n_1410),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1309),
.Y(n_1431)
);

CKINVDCx16_ASAP7_75t_R g1432 ( 
.A(n_1308),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1330),
.B(n_1312),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1374),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1374),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1342),
.B(n_1398),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1330),
.B(n_1312),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1308),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1334),
.B(n_1375),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1338),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1334),
.B(n_1375),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1347),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1347),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1317),
.A2(n_1318),
.B1(n_1335),
.B2(n_1364),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1314),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_1380),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1318),
.A2(n_1364),
.B1(n_1358),
.B2(n_1407),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1333),
.A2(n_1331),
.B(n_1341),
.C(n_1329),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1331),
.A2(n_1329),
.B(n_1353),
.C(n_1413),
.Y(n_1449)
);

O2A1O1Ixp5_ASAP7_75t_L g1450 ( 
.A1(n_1328),
.A2(n_1360),
.B(n_1357),
.C(n_1350),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1397),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1345),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1358),
.A2(n_1367),
.B1(n_1344),
.B2(n_1391),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1316),
.A2(n_1343),
.B(n_1355),
.C(n_1332),
.Y(n_1454)
);

NAND2x1_ASAP7_75t_L g1455 ( 
.A(n_1416),
.B(n_1379),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1401),
.B(n_1405),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1351),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1414),
.B(n_1344),
.Y(n_1458)
);

AOI211xp5_ASAP7_75t_L g1459 ( 
.A1(n_1338),
.A2(n_1403),
.B(n_1363),
.C(n_1348),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1306),
.B(n_1352),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1349),
.A2(n_1406),
.B(n_1404),
.C(n_1373),
.Y(n_1461)
);

O2A1O1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1349),
.A2(n_1404),
.B(n_1369),
.C(n_1373),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1402),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1316),
.A2(n_1305),
.B1(n_1408),
.B2(n_1302),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1403),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1336),
.B(n_1379),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1304),
.B(n_1392),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1302),
.A2(n_1408),
.B1(n_1387),
.B2(n_1305),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1304),
.B(n_1392),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1387),
.A2(n_1371),
.B1(n_1362),
.B2(n_1394),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1371),
.A2(n_1395),
.B1(n_1394),
.B2(n_1300),
.Y(n_1471)
);

INVx3_ASAP7_75t_SL g1472 ( 
.A(n_1371),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1395),
.A2(n_1388),
.B1(n_1346),
.B2(n_1325),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1324),
.B(n_1323),
.Y(n_1474)
);

CKINVDCx16_ASAP7_75t_R g1475 ( 
.A(n_1354),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_SL g1476 ( 
.A1(n_1346),
.A2(n_1356),
.B(n_1383),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1359),
.B(n_1390),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1393),
.A2(n_1415),
.B(n_1411),
.C(n_1360),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1359),
.B(n_1356),
.Y(n_1479)
);

AOI31xp33_ASAP7_75t_L g1480 ( 
.A1(n_1370),
.A2(n_1400),
.A3(n_1412),
.B(n_1381),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1393),
.B(n_1415),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1324),
.B(n_1323),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1307),
.A2(n_1315),
.B(n_1303),
.Y(n_1483)
);

OA22x2_ASAP7_75t_L g1484 ( 
.A1(n_1365),
.A2(n_1322),
.B1(n_1412),
.B2(n_1381),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1393),
.A2(n_1411),
.B(n_1313),
.C(n_1301),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1379),
.B(n_1301),
.Y(n_1486)
);

AND2x2_ASAP7_75t_SL g1487 ( 
.A(n_1313),
.B(n_1379),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1366),
.Y(n_1488)
);

O2A1O1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1313),
.A2(n_1384),
.B(n_1324),
.C(n_1379),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1324),
.B(n_1323),
.Y(n_1490)
);

O2A1O1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1361),
.A2(n_1273),
.B(n_1278),
.C(n_1376),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1361),
.B(n_1299),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1361),
.B(n_1299),
.Y(n_1493)
);

NOR4xp25_ASAP7_75t_L g1494 ( 
.A(n_1398),
.B(n_1282),
.C(n_1062),
.D(n_1376),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1386),
.A2(n_1398),
.B1(n_1282),
.B2(n_1310),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1386),
.A2(n_1398),
.B1(n_1282),
.B2(n_1310),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1386),
.A2(n_1398),
.B1(n_1282),
.B2(n_1310),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1326),
.B(n_1399),
.Y(n_1498)
);

O2A1O1Ixp33_ASAP7_75t_L g1499 ( 
.A1(n_1376),
.A2(n_1273),
.B(n_1278),
.C(n_1382),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1299),
.B(n_1320),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1310),
.A2(n_1282),
.B(n_997),
.C(n_1386),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1299),
.B(n_1320),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1321),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1309),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1386),
.A2(n_1398),
.B1(n_1282),
.B2(n_1310),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1385),
.A2(n_1278),
.B(n_1273),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1492),
.B(n_1493),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1477),
.B(n_1433),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_1418),
.Y(n_1509)
);

OAI21xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1423),
.A2(n_1424),
.B(n_1494),
.Y(n_1510)
);

NAND3xp33_ASAP7_75t_L g1511 ( 
.A(n_1501),
.B(n_1496),
.C(n_1495),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1497),
.B(n_1505),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1503),
.B(n_1498),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1421),
.B(n_1429),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1417),
.A2(n_1506),
.B(n_1420),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1484),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1460),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1455),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1451),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1474),
.B(n_1482),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1466),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1481),
.Y(n_1522)
);

AO21x2_ASAP7_75t_L g1523 ( 
.A1(n_1454),
.A2(n_1485),
.B(n_1478),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1457),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1490),
.B(n_1486),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1427),
.B(n_1425),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1480),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1450),
.Y(n_1528)
);

OR2x6_ASAP7_75t_L g1529 ( 
.A(n_1461),
.B(n_1462),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1487),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1428),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1483),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1434),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1419),
.A2(n_1437),
.B(n_1458),
.Y(n_1534)
);

AO21x2_ASAP7_75t_L g1535 ( 
.A1(n_1461),
.A2(n_1489),
.B(n_1491),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1489),
.A2(n_1491),
.B(n_1448),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1428),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1445),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1426),
.B(n_1439),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_1448),
.B(n_1499),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1430),
.B(n_1441),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1452),
.B(n_1435),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1499),
.B(n_1449),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1444),
.B(n_1447),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1463),
.B(n_1456),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1419),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1446),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1464),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1449),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1500),
.B(n_1502),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1453),
.B(n_1467),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1471),
.B(n_1436),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1470),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1468),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1473),
.Y(n_1555)
);

INVxp67_ASAP7_75t_SL g1556 ( 
.A(n_1528),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1522),
.B(n_1516),
.Y(n_1557)
);

NOR2xp67_ASAP7_75t_L g1558 ( 
.A(n_1517),
.B(n_1442),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1520),
.B(n_1525),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1521),
.B(n_1469),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1518),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1538),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1521),
.B(n_1459),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1520),
.B(n_1465),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_SL g1565 ( 
.A1(n_1511),
.A2(n_1475),
.B1(n_1432),
.B2(n_1438),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1518),
.Y(n_1566)
);

AND2x4_ASAP7_75t_SL g1567 ( 
.A(n_1530),
.B(n_1443),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1538),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1511),
.A2(n_1443),
.B1(n_1440),
.B2(n_1488),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1512),
.A2(n_1540),
.B1(n_1544),
.B2(n_1510),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1538),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1524),
.Y(n_1572)
);

OR2x6_ASAP7_75t_SL g1573 ( 
.A(n_1552),
.B(n_1422),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1530),
.B(n_1476),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1525),
.B(n_1443),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1519),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1510),
.A2(n_1479),
.B1(n_1504),
.B2(n_1431),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1532),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1507),
.B(n_1508),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1507),
.B(n_1508),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1570),
.A2(n_1540),
.B1(n_1573),
.B2(n_1543),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1562),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1562),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1559),
.B(n_1546),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_SL g1585 ( 
.A1(n_1574),
.A2(n_1515),
.B(n_1540),
.Y(n_1585)
);

AOI21xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1565),
.A2(n_1515),
.B(n_1540),
.Y(n_1586)
);

OAI31xp33_ASAP7_75t_L g1587 ( 
.A1(n_1570),
.A2(n_1549),
.A3(n_1548),
.B(n_1555),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1579),
.B(n_1530),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1573),
.B(n_1541),
.Y(n_1589)
);

OAI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1565),
.A2(n_1540),
.B1(n_1577),
.B2(n_1543),
.C(n_1569),
.Y(n_1590)
);

AOI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1569),
.A2(n_1549),
.B1(n_1526),
.B2(n_1536),
.C(n_1513),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1559),
.B(n_1534),
.Y(n_1592)
);

OAI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1573),
.A2(n_1543),
.B1(n_1552),
.B2(n_1551),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1577),
.A2(n_1543),
.B1(n_1536),
.B2(n_1555),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1561),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1564),
.A2(n_1543),
.B1(n_1536),
.B2(n_1534),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1579),
.B(n_1530),
.Y(n_1597)
);

NAND2xp33_ASAP7_75t_R g1598 ( 
.A(n_1563),
.B(n_1534),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1568),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1564),
.A2(n_1536),
.B1(n_1534),
.B2(n_1535),
.Y(n_1600)
);

OAI31xp33_ASAP7_75t_L g1601 ( 
.A1(n_1563),
.A2(n_1551),
.A3(n_1553),
.B(n_1527),
.Y(n_1601)
);

CKINVDCx16_ASAP7_75t_R g1602 ( 
.A(n_1564),
.Y(n_1602)
);

NAND3xp33_ASAP7_75t_L g1603 ( 
.A(n_1572),
.B(n_1529),
.C(n_1533),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1574),
.A2(n_1539),
.B1(n_1535),
.B2(n_1537),
.Y(n_1604)
);

NAND2xp33_ASAP7_75t_SL g1605 ( 
.A(n_1572),
.B(n_1550),
.Y(n_1605)
);

OAI31xp33_ASAP7_75t_L g1606 ( 
.A1(n_1567),
.A2(n_1554),
.A3(n_1547),
.B(n_1539),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1574),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1561),
.Y(n_1608)
);

INVx4_ASAP7_75t_L g1609 ( 
.A(n_1574),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1579),
.B(n_1535),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1574),
.A2(n_1535),
.B1(n_1537),
.B2(n_1531),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1556),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1561),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1580),
.B(n_1523),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1580),
.B(n_1523),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1578),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1571),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1559),
.B(n_1509),
.Y(n_1618)
);

OAI31xp33_ASAP7_75t_L g1619 ( 
.A1(n_1567),
.A2(n_1554),
.A3(n_1545),
.B(n_1514),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1580),
.B(n_1523),
.Y(n_1620)
);

NAND3xp33_ASAP7_75t_SL g1621 ( 
.A(n_1576),
.B(n_1542),
.C(n_1545),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1566),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1599),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1585),
.B(n_1574),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1599),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1601),
.B(n_1560),
.Y(n_1626)
);

AO21x1_ASAP7_75t_L g1627 ( 
.A1(n_1598),
.A2(n_1560),
.B(n_1556),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1589),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1584),
.B(n_1576),
.Y(n_1629)
);

INVx4_ASAP7_75t_SL g1630 ( 
.A(n_1607),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1608),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1616),
.Y(n_1632)
);

BUFx8_ASAP7_75t_L g1633 ( 
.A(n_1607),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1617),
.Y(n_1634)
);

AND2x4_ASAP7_75t_SL g1635 ( 
.A(n_1588),
.B(n_1597),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1610),
.B(n_1557),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1608),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_SL g1638 ( 
.A1(n_1591),
.A2(n_1529),
.B(n_1566),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1602),
.Y(n_1639)
);

BUFx8_ASAP7_75t_L g1640 ( 
.A(n_1607),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1608),
.Y(n_1641)
);

CKINVDCx14_ASAP7_75t_R g1642 ( 
.A(n_1581),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1613),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1593),
.B(n_1558),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1582),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1582),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1583),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1601),
.B(n_1575),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1591),
.A2(n_1529),
.B(n_1523),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1583),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1613),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1613),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1618),
.B(n_1575),
.Y(n_1653)
);

OA21x2_ASAP7_75t_L g1654 ( 
.A1(n_1600),
.A2(n_1592),
.B(n_1596),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1610),
.B(n_1557),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1623),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1630),
.B(n_1614),
.Y(n_1657)
);

NOR2x1_ASAP7_75t_L g1658 ( 
.A(n_1638),
.B(n_1621),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1630),
.B(n_1614),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1630),
.B(n_1610),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1627),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1630),
.B(n_1614),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1645),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1633),
.Y(n_1664)
);

NAND2x1_ASAP7_75t_L g1665 ( 
.A(n_1638),
.B(n_1595),
.Y(n_1665)
);

AND4x1_ASAP7_75t_L g1666 ( 
.A(n_1649),
.B(n_1587),
.C(n_1594),
.D(n_1596),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1635),
.B(n_1609),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1629),
.B(n_1584),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1623),
.Y(n_1669)
);

BUFx2_ASAP7_75t_SL g1670 ( 
.A(n_1627),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1624),
.B(n_1609),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1632),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1625),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1632),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1625),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1634),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1626),
.B(n_1592),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1648),
.B(n_1615),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1634),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1639),
.B(n_1615),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1642),
.B(n_1620),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1633),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1628),
.B(n_1602),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1636),
.B(n_1622),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1645),
.B(n_1646),
.Y(n_1685)
);

INVx4_ASAP7_75t_L g1686 ( 
.A(n_1637),
.Y(n_1686)
);

OAI222xp33_ASAP7_75t_L g1687 ( 
.A1(n_1624),
.A2(n_1590),
.B1(n_1581),
.B2(n_1593),
.C1(n_1604),
.C2(n_1611),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1633),
.Y(n_1688)
);

OAI31xp33_ASAP7_75t_L g1689 ( 
.A1(n_1644),
.A2(n_1590),
.A3(n_1587),
.B(n_1603),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1643),
.B(n_1588),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1646),
.B(n_1612),
.Y(n_1691)
);

OAI21xp33_ASAP7_75t_L g1692 ( 
.A1(n_1624),
.A2(n_1586),
.B(n_1603),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1655),
.B(n_1622),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1681),
.B(n_1631),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1681),
.B(n_1631),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1662),
.B(n_1631),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1663),
.Y(n_1697)
);

NOR2xp67_ASAP7_75t_SL g1698 ( 
.A(n_1670),
.B(n_1607),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1663),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1668),
.B(n_1629),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1656),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1693),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1683),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1662),
.B(n_1657),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1667),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1677),
.B(n_1654),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1677),
.B(n_1654),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1664),
.B(n_1654),
.Y(n_1708)
);

AOI211xp5_ASAP7_75t_L g1709 ( 
.A1(n_1687),
.A2(n_1586),
.B(n_1607),
.C(n_1621),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1664),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1667),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1656),
.Y(n_1712)
);

OAI21xp33_ASAP7_75t_L g1713 ( 
.A1(n_1666),
.A2(n_1624),
.B(n_1653),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1668),
.B(n_1647),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1664),
.B(n_1654),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1669),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1657),
.B(n_1643),
.Y(n_1717)
);

OAI31xp33_ASAP7_75t_L g1718 ( 
.A1(n_1692),
.A2(n_1605),
.A3(n_1619),
.B(n_1606),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1691),
.B(n_1647),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1667),
.B(n_1637),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1689),
.B(n_1640),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1669),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1684),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1682),
.B(n_1641),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1691),
.B(n_1650),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1657),
.B(n_1641),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1659),
.B(n_1651),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1659),
.B(n_1651),
.Y(n_1728)
);

OAI31xp33_ASAP7_75t_L g1729 ( 
.A1(n_1692),
.A2(n_1619),
.A3(n_1606),
.B(n_1652),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1717),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1720),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1697),
.Y(n_1732)
);

NAND2xp33_ASAP7_75t_SL g1733 ( 
.A(n_1721),
.B(n_1665),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1700),
.B(n_1714),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1717),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1726),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1704),
.B(n_1658),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1702),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1697),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1702),
.Y(n_1740)
);

INVx1_ASAP7_75t_SL g1741 ( 
.A(n_1726),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1709),
.A2(n_1670),
.B1(n_1661),
.B2(n_1666),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1700),
.B(n_1685),
.Y(n_1743)
);

CKINVDCx16_ASAP7_75t_R g1744 ( 
.A(n_1710),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1724),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1727),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1699),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1699),
.Y(n_1748)
);

INVx3_ASAP7_75t_SL g1749 ( 
.A(n_1720),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1723),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1704),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1701),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1723),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1727),
.B(n_1658),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1705),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1742),
.A2(n_1713),
.B(n_1661),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1751),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1734),
.Y(n_1758)
);

OAI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1733),
.A2(n_1689),
.B1(n_1718),
.B2(n_1729),
.C(n_1665),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1744),
.B(n_1703),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1744),
.B(n_1728),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1745),
.B(n_1682),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1749),
.A2(n_1688),
.B1(n_1682),
.B2(n_1678),
.Y(n_1763)
);

NOR2x1p5_ASAP7_75t_SL g1764 ( 
.A(n_1730),
.B(n_1701),
.Y(n_1764)
);

AOI31xp33_ASAP7_75t_L g1765 ( 
.A1(n_1736),
.A2(n_1688),
.A3(n_1711),
.B(n_1705),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1754),
.B(n_1728),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1737),
.A2(n_1707),
.B1(n_1706),
.B2(n_1671),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1741),
.B(n_1746),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_SL g1769 ( 
.A1(n_1754),
.A2(n_1698),
.B(n_1715),
.C(n_1708),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1755),
.Y(n_1770)
);

AOI222xp33_ASAP7_75t_L g1771 ( 
.A1(n_1737),
.A2(n_1687),
.B1(n_1698),
.B2(n_1678),
.C1(n_1695),
.C2(n_1694),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1731),
.A2(n_1711),
.B(n_1720),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_L g1773 ( 
.A(n_1731),
.B(n_1686),
.C(n_1719),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1734),
.A2(n_1695),
.B(n_1694),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1730),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1730),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1757),
.B(n_1735),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1766),
.B(n_1749),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1757),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1760),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1774),
.B(n_1749),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1761),
.B(n_1735),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1770),
.B(n_1735),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1768),
.B(n_1743),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1770),
.B(n_1732),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1762),
.B(n_1688),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1758),
.B(n_1732),
.Y(n_1787)
);

OAI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1780),
.A2(n_1756),
.B1(n_1759),
.B2(n_1771),
.C(n_1769),
.Y(n_1788)
);

AOI21xp33_ASAP7_75t_L g1789 ( 
.A1(n_1784),
.A2(n_1765),
.B(n_1773),
.Y(n_1789)
);

OAI32xp33_ASAP7_75t_L g1790 ( 
.A1(n_1785),
.A2(n_1763),
.A3(n_1772),
.B1(n_1767),
.B2(n_1775),
.Y(n_1790)
);

AOI21xp33_ASAP7_75t_SL g1791 ( 
.A1(n_1786),
.A2(n_1776),
.B(n_1747),
.Y(n_1791)
);

AOI221x1_ASAP7_75t_L g1792 ( 
.A1(n_1779),
.A2(n_1748),
.B1(n_1747),
.B2(n_1739),
.C(n_1750),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1785),
.A2(n_1748),
.B(n_1739),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1777),
.A2(n_1740),
.B(n_1738),
.Y(n_1794)
);

AOI211xp5_ASAP7_75t_L g1795 ( 
.A1(n_1778),
.A2(n_1752),
.B(n_1753),
.C(n_1740),
.Y(n_1795)
);

AOI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1783),
.A2(n_1752),
.B1(n_1743),
.B2(n_1738),
.C(n_1750),
.Y(n_1796)
);

NOR3x1_ASAP7_75t_L g1797 ( 
.A(n_1777),
.B(n_1725),
.C(n_1719),
.Y(n_1797)
);

OAI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1788),
.A2(n_1686),
.B1(n_1787),
.B2(n_1740),
.Y(n_1798)
);

OAI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1789),
.A2(n_1781),
.B1(n_1795),
.B2(n_1796),
.C(n_1793),
.Y(n_1799)
);

O2A1O1Ixp33_ASAP7_75t_L g1800 ( 
.A1(n_1790),
.A2(n_1782),
.B(n_1764),
.C(n_1738),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1794),
.A2(n_1753),
.B(n_1750),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1792),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1800),
.B(n_1791),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1802),
.B(n_1797),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1799),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1801),
.B(n_1696),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1798),
.B(n_1725),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1800),
.B(n_1753),
.Y(n_1808)
);

AOI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1803),
.A2(n_1722),
.B1(n_1716),
.B2(n_1712),
.C(n_1686),
.Y(n_1809)
);

XNOR2xp5_ASAP7_75t_L g1810 ( 
.A(n_1805),
.B(n_1696),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1804),
.A2(n_1686),
.B1(n_1671),
.B2(n_1659),
.Y(n_1811)
);

OAI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1806),
.A2(n_1716),
.B(n_1712),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1807),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1813),
.B(n_1808),
.Y(n_1814)
);

NAND4xp25_ASAP7_75t_SL g1815 ( 
.A(n_1811),
.B(n_1722),
.C(n_1660),
.D(n_1714),
.Y(n_1815)
);

NOR2x1_ASAP7_75t_L g1816 ( 
.A(n_1810),
.B(n_1685),
.Y(n_1816)
);

NAND4xp75_ASAP7_75t_L g1817 ( 
.A(n_1814),
.B(n_1809),
.C(n_1812),
.D(n_1680),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1817),
.B(n_1816),
.Y(n_1818)
);

XOR2x2_ASAP7_75t_L g1819 ( 
.A(n_1818),
.B(n_1815),
.Y(n_1819)
);

OR4x1_ASAP7_75t_L g1820 ( 
.A(n_1818),
.B(n_1676),
.C(n_1679),
.D(n_1673),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1819),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1820),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1822),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_1821),
.B1(n_1672),
.B2(n_1674),
.Y(n_1824)
);

AOI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1824),
.A2(n_1671),
.B1(n_1667),
.B2(n_1680),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1825),
.B(n_1690),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1826),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1827),
.A2(n_1671),
.B1(n_1690),
.B2(n_1675),
.Y(n_1828)
);

AOI211xp5_ASAP7_75t_L g1829 ( 
.A1(n_1828),
.A2(n_1472),
.B(n_1679),
.C(n_1676),
.Y(n_1829)
);


endmodule