module real_jpeg_31612_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_553;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g168 ( 
.A(n_0),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_0),
.Y(n_294)
);

BUFx12f_ASAP7_75t_L g339 ( 
.A(n_0),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_0),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_0),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_1),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_1),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_1),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_1),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_1),
.B(n_39),
.Y(n_337)
);

AND2x2_ASAP7_75t_SL g468 ( 
.A(n_1),
.B(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_1),
.B(n_495),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_2),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_2),
.B(n_333),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_2),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_2),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_2),
.B(n_504),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_2),
.B(n_509),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_2),
.B(n_514),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_22),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_3),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_6),
.Y(n_301)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_7),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_7),
.Y(n_199)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_7),
.Y(n_280)
);

AND2x4_ASAP7_75t_L g33 ( 
.A(n_8),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_8),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_8),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_8),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_8),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_8),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_8),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_9),
.B(n_44),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_9),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_9),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_9),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_9),
.B(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_9),
.B(n_491),
.Y(n_490)
);

AND2x2_ASAP7_75t_SL g501 ( 
.A(n_9),
.B(n_254),
.Y(n_501)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_10),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_10),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_10),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_11),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_12),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_12),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g270 ( 
.A(n_12),
.B(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_12),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_12),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_12),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_12),
.B(n_443),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_12),
.B(n_472),
.Y(n_471)
);

AND2x6_ASAP7_75t_SL g66 ( 
.A(n_13),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_13),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_13),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_13),
.B(n_156),
.Y(n_155)
);

NAND2x1_ASAP7_75t_L g205 ( 
.A(n_13),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_13),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_13),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_13),
.B(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_14),
.Y(n_106)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_14),
.Y(n_145)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_14),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_15),
.Y(n_92)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_15),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_30),
.Y(n_29)
);

NAND2x1_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_16),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_16),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_16),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_16),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_17),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_17),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_17),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_17),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_17),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_17),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_17),
.B(n_339),
.Y(n_338)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_114),
.A3(n_115),
.B1(n_538),
.B2(n_544),
.C(n_550),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI322xp5_ASAP7_75t_L g550 ( 
.A1(n_20),
.A2(n_538),
.A3(n_545),
.B1(n_548),
.B2(n_551),
.C1(n_552),
.C2(n_553),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_21),
.B(n_546),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_21),
.Y(n_553)
);

INVxp33_ASAP7_75t_L g546 ( 
.A(n_23),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_113),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_76),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_25),
.B(n_76),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_51),
.Y(n_25)
);

BUFx24_ASAP7_75t_SL g554 ( 
.A(n_26),
.Y(n_554)
);

FAx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_41),
.CI(n_46),
.CON(n_26),
.SN(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.C(n_37),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_28),
.A2(n_29),
.B1(n_71),
.B2(n_72),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_28),
.B(n_136),
.C(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_28),
.A2(n_29),
.B1(n_238),
.B2(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_29),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_32),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_32),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_32),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_37),
.B1(n_38),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_33),
.B(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_33),
.B(n_129),
.C(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_36),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_36),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_38),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_37),
.B(n_246),
.C(n_252),
.Y(n_245)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2x1_ASAP7_75t_L g385 ( 
.A(n_38),
.B(n_253),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_R g83 ( 
.A(n_41),
.B(n_84),
.C(n_88),
.Y(n_83)
);

XOR2x2_ASAP7_75t_L g121 ( 
.A(n_41),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_45),
.Y(n_195)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_47),
.B(n_160),
.C(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_47),
.B(n_161),
.Y(n_202)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.C(n_64),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_65),
.C(n_71),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_59),
.B1(n_64),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_70),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_70),
.Y(n_211)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_70),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_103),
.C(n_107),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_R g177 ( 
.A1(n_71),
.A2(n_72),
.B1(n_103),
.B2(n_154),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_71),
.B(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_71),
.B(n_142),
.C(n_343),
.Y(n_369)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_73),
.Y(n_313)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.C(n_96),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_77),
.A2(n_78),
.B1(n_81),
.B2(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g542 ( 
.A(n_81),
.Y(n_542)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_90),
.C(n_93),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_83),
.B1(n_98),
.B2(n_100),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_84),
.A2(n_88),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_88),
.B(n_205),
.C(n_208),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_88),
.A2(n_124),
.B1(n_208),
.B2(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_165),
.C(n_169),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_90),
.B(n_204),
.C(n_210),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_90),
.A2(n_91),
.B1(n_169),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_90),
.A2(n_91),
.B1(n_210),
.B2(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_92),
.Y(n_320)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_96),
.B(n_541),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.C(n_111),
.Y(n_96)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_97),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2x1_ASAP7_75t_L g173 ( 
.A(n_102),
.B(n_111),
.Y(n_173)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_103),
.B(n_155),
.C(n_160),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_103),
.B(n_297),
.C(n_303),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_103),
.B(n_297),
.Y(n_309)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_106),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_177),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21x1_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_262),
.B(n_533),
.Y(n_115)
);

NAND2x1_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_222),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_118),
.A2(n_535),
.B(n_536),
.Y(n_534)
);

AOI21x1_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_180),
.B(n_183),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_171),
.Y(n_119)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_120),
.A2(n_171),
.B1(n_181),
.B2(n_182),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_120),
.B(n_172),
.C(n_175),
.Y(n_543)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.C(n_164),
.Y(n_120)
);

XNOR2x1_ASAP7_75t_SL g221 ( 
.A(n_121),
.B(n_164),
.Y(n_221)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_126),
.B(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_138),
.C(n_151),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_127),
.B(n_138),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_132),
.B1(n_136),
.B2(n_137),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_129),
.A2(n_136),
.B1(n_371),
.B2(n_373),
.Y(n_370)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_130),
.Y(n_505)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_146),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_139),
.A2(n_146),
.B1(n_147),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_143),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_142),
.A2(n_143),
.B1(n_343),
.B2(n_346),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_145),
.Y(n_440)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_151),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_160),
.B2(n_161),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_158),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_159),
.Y(n_364)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_161),
.B(n_250),
.Y(n_436)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_163),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_165),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_197),
.Y(n_200)
);

XOR2x2_ASAP7_75t_SL g201 ( 
.A(n_166),
.B(n_202),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g242 ( 
.A(n_166),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_166),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_166),
.A2(n_442),
.B1(n_444),
.B2(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_168),
.Y(n_251)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_179),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_179),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_183),
.B(n_537),
.Y(n_536)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_216),
.C(n_219),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_185),
.B(n_261),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_203),
.C(n_212),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_192),
.C(n_201),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_188),
.B(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_192),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_196),
.B(n_200),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_193),
.A2(n_194),
.B1(n_197),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_197),
.B(n_290),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_197),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_198),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_199),
.Y(n_470)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_199),
.Y(n_493)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_200),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_200),
.A2(n_327),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_201),
.B(n_411),
.Y(n_410)
);

XNOR2x1_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_213),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_204),
.B(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_207),
.Y(n_305)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_209),
.Y(n_334)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_220),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_260),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_223),
.B(n_260),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.C(n_231),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_225),
.B(n_228),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_231),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_245),
.C(n_256),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_232),
.A2(n_233),
.B1(n_406),
.B2(n_407),
.Y(n_405)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_242),
.Y(n_233)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_234),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_237),
.B(n_242),
.Y(n_390)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_238),
.Y(n_372)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_245),
.A2(n_256),
.B1(n_257),
.B2(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_245),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_246),
.B(n_385),
.Y(n_384)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.C(n_250),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_247),
.B(n_249),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_250),
.B(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_425),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_394),
.B1(n_419),
.B2(n_424),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_374),
.B(n_391),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_347),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_266),
.B(n_347),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_307),
.C(n_324),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_267),
.B(n_325),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_287),
.B2(n_306),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_268),
.B(n_288),
.C(n_296),
.Y(n_356)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g354 ( 
.A(n_270),
.B(n_276),
.C(n_281),
.Y(n_354)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_281),
.B2(n_282),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_295),
.B2(n_296),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_290),
.A2(n_291),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_294),
.Y(n_472)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_302),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_302),
.B(n_465),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_303),
.B(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_307),
.B(n_431),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.C(n_321),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_308),
.B(n_434),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_310),
.B(n_321),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.C(n_317),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_311),
.B(n_480),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_315),
.B(n_318),
.Y(n_480)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_316),
.Y(n_462)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_335),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_326),
.B(n_336),
.C(n_341),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.C(n_331),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_328),
.A2(n_329),
.B1(n_331),
.B2(n_332),
.Y(n_446)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_341),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B(n_340),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_338),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_354),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_351),
.C(n_354),
.Y(n_382)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_355),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

MAJx2_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_350),
.C(n_355),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_358),
.C(n_370),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_370),
.Y(n_357)
);

XNOR2x2_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_368),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_365),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_365),
.C(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_369),
.Y(n_387)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_371),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

AOI21x1_ASAP7_75t_L g391 ( 
.A1(n_375),
.A2(n_392),
.B(n_393),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_379),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_397),
.C(n_398),
.Y(n_396)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_380),
.Y(n_392)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_388),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_381),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_384),
.C(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_386),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_388),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_391),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_414),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_400),
.Y(n_395)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_396),
.Y(n_422)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_400),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_405),
.C(n_409),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_409),
.B1(n_410),
.B2(n_413),
.Y(n_404)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_405),
.Y(n_413)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_414),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_415),
.Y(n_421)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_416),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_426),
.C(n_428),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_422),
.B2(n_423),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_448),
.B(n_532),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_432),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_430),
.B(n_432),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.C(n_445),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_433),
.B(n_530),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_435),
.B(n_445),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.C(n_441),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_436),
.A2(n_437),
.B1(n_438),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_436),
.Y(n_485)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_440),
.Y(n_466)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_440),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_441),
.B(n_484),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.Y(n_441)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_442),
.Y(n_475)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_446),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_526),
.B(n_531),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_450),
.A2(n_486),
.B(n_525),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_476),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_451),
.B(n_476),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_467),
.C(n_473),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_452),
.A2(n_453),
.B1(n_521),
.B2(n_523),
.Y(n_520)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_464),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_456),
.B1(n_460),
.B2(n_463),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_463),
.C(n_464),
.Y(n_478)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_460),
.Y(n_463)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_467),
.A2(n_473),
.B1(n_474),
.B2(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_467),
.Y(n_522)
);

NAND2x1_ASAP7_75t_SL g467 ( 
.A(n_468),
.B(n_471),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_468),
.B(n_471),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_483),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_481),
.B2(n_482),
.Y(n_477)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_478),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_479),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_479),
.B(n_481),
.C(n_528),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_483),
.Y(n_528)
);

AOI21x1_ASAP7_75t_SL g486 ( 
.A1(n_487),
.A2(n_518),
.B(n_524),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_488),
.A2(n_506),
.B(n_517),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_497),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_489),
.B(n_497),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_494),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_490),
.B(n_494),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_490),
.B(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

BUFx4f_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_501),
.C(n_502),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_500),
.A2(n_501),
.B1(n_502),
.B2(n_503),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_507),
.A2(n_512),
.B(n_516),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_511),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_508),
.B(n_511),
.Y(n_516)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_520),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_SL g524 ( 
.A(n_519),
.B(n_520),
.Y(n_524)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_521),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_529),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_529),
.Y(n_531)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_539),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_543),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_540),
.B(n_543),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_547),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_549),
.Y(n_551)
);


endmodule