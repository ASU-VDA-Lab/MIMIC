module fake_jpeg_9073_n_45 (n_3, n_2, n_1, n_0, n_4, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_3),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx2_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

NOR3xp33_ASAP7_75t_SL g23 ( 
.A(n_14),
.B(n_15),
.C(n_16),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_0),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_3),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_2),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_19),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_6),
.A2(n_3),
.B1(n_5),
.B2(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

NOR2x1_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_16),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

AO221x1_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_16),
.B1(n_18),
.B2(n_23),
.C(n_20),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_37),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_33),
.C(n_32),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_20),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_23),
.A3(n_18),
.B1(n_13),
.B2(n_9),
.C1(n_7),
.C2(n_11),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_7),
.B(n_11),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_41),
.B(n_7),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_9),
.B1(n_11),
.B2(n_38),
.Y(n_45)
);


endmodule