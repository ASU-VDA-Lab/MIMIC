module real_jpeg_24669_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_215;
wire n_221;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_4),
.A2(n_7),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_4),
.A2(n_33),
.B1(n_47),
.B2(n_48),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_4),
.A2(n_33),
.B1(n_52),
.B2(n_53),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_4),
.B(n_22),
.C(n_24),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_21),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_4),
.B(n_48),
.C(n_59),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_4),
.B(n_49),
.C(n_52),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_4),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_4),
.B(n_72),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_4),
.B(n_77),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_30),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_6),
.A2(n_30),
.B1(n_47),
.B2(n_48),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_6),
.A2(n_30),
.B1(n_52),
.B2(n_53),
.Y(n_173)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_55),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_62),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_11),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_109),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_108),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_15),
.B(n_93),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_68),
.C(n_78),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_16),
.A2(n_17),
.B1(n_68),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_38),
.B2(n_39),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_18),
.B(n_41),
.C(n_56),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_18),
.A2(n_19),
.B1(n_98),
.B2(n_107),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_18),
.B(n_125),
.C(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_18),
.A2(n_19),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_18),
.A2(n_19),
.B1(n_147),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_19),
.B(n_139),
.C(n_147),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_27),
.B(n_31),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_36),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_21),
.A2(n_32),
.B1(n_36),
.B2(n_104),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_26),
.B1(n_28),
.B2(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_23),
.A2(n_24),
.B1(n_58),
.B2(n_59),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_24),
.B(n_203),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_35),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_56),
.B2(n_67),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_40),
.A2(n_41),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_54),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_43),
.B(n_88),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_51),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_45),
.A2(n_72),
.B1(n_88),
.B2(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

OA22x2_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_48),
.B(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_71),
.B(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_51),
.A2(n_87),
.B(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_52),
.B(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_63),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_57),
.A2(n_63),
.B(n_76),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_57),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_61),
.A2(n_64),
.B1(n_77),
.B2(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_66),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_64),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_68),
.A2(n_69),
.B(n_74),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_68),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_74),
.A2(n_103),
.B1(n_106),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_74),
.B(n_187),
.C(n_189),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_74),
.A2(n_177),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_74),
.B(n_103),
.C(n_166),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_128),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_85),
.B(n_89),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_89),
.B1(n_90),
.B2(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_79),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_79),
.A2(n_86),
.B1(n_115),
.B2(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_81),
.B(n_175),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_84),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_83),
.A2(n_120),
.B(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_83),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_86),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_103),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_118),
.C(n_125),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_106),
.B1(n_125),
.B2(n_126),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_130),
.B(n_271),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_127),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_112),
.B(n_127),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_117),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_116),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_119),
.A2(n_122),
.B1(n_123),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_119),
.Y(n_262)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_122),
.A2(n_123),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_122),
.A2(n_123),
.B1(n_200),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_194),
.C(n_200),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_123),
.B(n_171),
.C(n_233),
.Y(n_237)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_125),
.A2(n_126),
.B1(n_162),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_125),
.A2(n_126),
.B1(n_145),
.B2(n_159),
.Y(n_239)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_126),
.B(n_145),
.C(n_240),
.Y(n_243)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_152),
.B(n_270),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_150),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_133),
.B(n_150),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.C(n_138),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_134),
.B(n_136),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_138),
.B(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_139),
.A2(n_140),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_145),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_141),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_143),
.A2(n_173),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_145),
.A2(n_159),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_145),
.B(n_217),
.Y(n_229)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_147),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_265),
.B(n_269),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_190),
.B(n_251),
.C(n_264),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_179),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_155),
.B(n_179),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_165),
.B2(n_178),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_158),
.B(n_164),
.C(n_178),
.Y(n_252)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_176),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_170),
.A2(n_171),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_171),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_225),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.C(n_186),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_181),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_186),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_189),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_187),
.B(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_250),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_209),
.B(n_249),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_206),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_193),
.B(n_206),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_195),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_199),
.B(n_214),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_242),
.B(n_248),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_236),
.B(n_241),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_228),
.B(n_235),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_218),
.B(n_227),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_215),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_224),
.B(n_226),
.Y(n_218)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_229),
.B(n_230),
.Y(n_235)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_253),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_263),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_260),
.B2(n_261),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_261),
.C(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_267),
.Y(n_269)
);


endmodule