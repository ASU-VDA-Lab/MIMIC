module fake_jpeg_13788_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_23),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_0),
.B(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_27),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_16),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NAND2x1p5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_51),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_72),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_74),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_1),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_84),
.B(n_78),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_62),
.B(n_50),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_38),
.C(n_29),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_92),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_91),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_43),
.B1(n_42),
.B2(n_46),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_50),
.B1(n_47),
.B2(n_42),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_2),
.Y(n_94)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_98),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_78),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_97),
.C(n_101),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_20),
.B(n_37),
.C(n_35),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_12),
.C(n_34),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_105),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_4),
.Y(n_101)
);

NOR4xp25_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_18),
.C(n_32),
.D(n_30),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_28),
.C(n_26),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_5),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_107),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_112),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_114),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_21),
.C(n_91),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_118),
.B(n_100),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_106),
.C(n_8),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_6),
.C(n_7),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_120),
.C(n_115),
.Y(n_124)
);

AOI322xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_96),
.A3(n_100),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_8),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_113),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_123),
.A2(n_113),
.B(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

OAI21x1_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_121),
.B(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_127),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_110),
.C(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_120),
.Y(n_133)
);


endmodule