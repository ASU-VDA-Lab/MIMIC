module fake_jpeg_31063_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

AND2x2_ASAP7_75t_SL g7 ( 
.A(n_4),
.B(n_2),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx24_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_4),
.B(n_6),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_5),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_20),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_10),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_7),
.B1(n_9),
.B2(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_13),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_14),
.B(n_7),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_7),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_7),
.B1(n_21),
.B2(n_9),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_16),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_7),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_23),
.C(n_24),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_26),
.B1(n_21),
.B2(n_19),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_25),
.C(n_29),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_34),
.C(n_32),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_13),
.C(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_31),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_38),
.B(n_9),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_33),
.B(n_18),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_8),
.B(n_3),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_22),
.C(n_10),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_10),
.C(n_13),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_47),
.C(n_48),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_9),
.B(n_8),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_44),
.C(n_5),
.Y(n_51)
);

AOI31xp33_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_1),
.A3(n_6),
.B(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_55),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_51),
.B(n_6),
.Y(n_55)
);


endmodule