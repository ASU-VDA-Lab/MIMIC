module fake_jpeg_845_n_28 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_28);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_28;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_10),
.B(n_9),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_1),
.C(n_2),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_10),
.A2(n_8),
.B1(n_7),
.B2(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_4),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_16),
.A2(n_3),
.B(n_4),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_21),
.C(n_16),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_24),
.C(n_18),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_24)
);

AOI322xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_5),
.A3(n_6),
.B1(n_17),
.B2(n_18),
.C1(n_21),
.C2(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_26),
.Y(n_27)
);

MAJx2_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_22),
.C(n_17),
.Y(n_28)
);


endmodule