module real_aes_9966_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_0), .A2(n_194), .B1(n_958), .B2(n_960), .Y(n_957) );
AOI22xp33_ASAP7_75t_SL g997 ( .A1(n_0), .A2(n_4), .B1(n_384), .B2(n_998), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_1), .A2(n_403), .B1(n_653), .B2(n_655), .C(n_661), .Y(n_652) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_1), .A2(n_698), .B(n_699), .Y(n_697) );
AOI21xp33_ASAP7_75t_L g1029 ( .A1(n_2), .A2(n_461), .B(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1050 ( .A(n_2), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_3), .A2(n_62), .B1(n_1129), .B2(n_1145), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g955 ( .A1(n_4), .A2(n_162), .B1(n_454), .B2(n_908), .C(n_956), .Y(n_955) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_5), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_5), .B(n_182), .Y(n_353) );
AND2x2_ASAP7_75t_L g369 ( .A(n_5), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g441 ( .A(n_5), .Y(n_441) );
INVx1_ASAP7_75t_L g520 ( .A(n_6), .Y(n_520) );
INVxp67_ASAP7_75t_L g1405 ( .A(n_7), .Y(n_1405) );
OAI222xp33_ASAP7_75t_L g1419 ( .A1(n_7), .A2(n_41), .B1(n_241), .B2(n_470), .C1(n_574), .C2(n_646), .Y(n_1419) );
OAI221xp5_ASAP7_75t_L g731 ( .A1(n_8), .A2(n_545), .B1(n_732), .B2(n_738), .C(n_743), .Y(n_731) );
INVx1_ASAP7_75t_L g757 ( .A(n_8), .Y(n_757) );
INVx1_ASAP7_75t_L g526 ( .A(n_9), .Y(n_526) );
XNOR2x2_ASAP7_75t_L g876 ( .A(n_10), .B(n_877), .Y(n_876) );
AOI221xp5_ASAP7_75t_L g838 ( .A1(n_11), .A2(n_164), .B1(n_302), .B2(n_839), .C(n_840), .Y(n_838) );
INVx1_ASAP7_75t_L g861 ( .A(n_11), .Y(n_861) );
OAI221xp5_ASAP7_75t_L g666 ( .A1(n_12), .A2(n_21), .B1(n_391), .B2(n_397), .C(n_401), .Y(n_666) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_12), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_13), .A2(n_52), .B1(n_373), .B2(n_531), .C(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g762 ( .A(n_13), .Y(n_762) );
INVx1_ASAP7_75t_L g720 ( .A(n_14), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_14), .A2(n_54), .B1(n_303), .B2(n_593), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_15), .A2(n_77), .B1(n_848), .B2(n_1069), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_15), .A2(n_30), .B1(n_495), .B2(n_537), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_16), .A2(n_222), .B1(n_848), .B2(n_850), .Y(n_847) );
INVx1_ASAP7_75t_L g869 ( .A(n_16), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_17), .A2(n_37), .B1(n_302), .B2(n_946), .Y(n_945) );
INVxp33_ASAP7_75t_SL g987 ( .A(n_17), .Y(n_987) );
AOI22xp5_ASAP7_75t_L g1136 ( .A1(n_18), .A2(n_68), .B1(n_1125), .B2(n_1129), .Y(n_1136) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_19), .A2(n_233), .B1(n_282), .B2(n_289), .C(n_293), .Y(n_281) );
INVx1_ASAP7_75t_L g377 ( .A(n_19), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g1013 ( .A1(n_20), .A2(n_681), .B1(n_1014), .B2(n_1018), .C(n_1021), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_20), .A2(n_165), .B1(n_1038), .B2(n_1047), .Y(n_1046) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_21), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g739 ( .A(n_22), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g1091 ( .A1(n_23), .A2(n_138), .B1(n_531), .B2(n_1038), .C(n_1092), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_23), .A2(n_209), .B1(n_563), .B2(n_641), .Y(n_1100) );
INVx2_ASAP7_75t_L g296 ( .A(n_24), .Y(n_296) );
OR2x2_ASAP7_75t_L g308 ( .A(n_24), .B(n_309), .Y(n_308) );
AO22x1_ASAP7_75t_L g715 ( .A1(n_25), .A2(n_716), .B1(n_764), .B2(n_765), .Y(n_715) );
INVx1_ASAP7_75t_L g765 ( .A(n_25), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g1135 ( .A1(n_26), .A2(n_117), .B1(n_1113), .B2(n_1121), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_27), .A2(n_61), .B1(n_1065), .B2(n_1066), .Y(n_1064) );
INVx1_ASAP7_75t_L g1087 ( .A(n_27), .Y(n_1087) );
OAI221xp5_ASAP7_75t_L g782 ( .A1(n_28), .A2(n_96), .B1(n_396), .B2(n_783), .C(n_785), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_28), .A2(n_96), .B1(n_319), .B2(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g1406 ( .A(n_29), .Y(n_1406) );
OAI222xp33_ASAP7_75t_L g1099 ( .A1(n_30), .A2(n_138), .B1(n_143), .B2(n_354), .C1(n_643), .C2(n_645), .Y(n_1099) );
BUFx2_ASAP7_75t_L g278 ( .A(n_31), .Y(n_278) );
OR2x2_ASAP7_75t_L g352 ( .A(n_31), .B(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g356 ( .A(n_31), .Y(n_356) );
INVx1_ASAP7_75t_L g368 ( .A(n_31), .Y(n_368) );
INVx1_ASAP7_75t_L g1161 ( .A(n_32), .Y(n_1161) );
INVx1_ASAP7_75t_L g1429 ( .A(n_33), .Y(n_1429) );
OAI221xp5_ASAP7_75t_L g1435 ( .A1(n_33), .A2(n_73), .B1(n_1436), .B2(n_1437), .C(n_1439), .Y(n_1435) );
AOI22xp33_ASAP7_75t_SL g660 ( .A1(n_34), .A2(n_147), .B1(n_539), .B2(n_611), .Y(n_660) );
INVx1_ASAP7_75t_L g688 ( .A(n_34), .Y(n_688) );
INVx1_ASAP7_75t_L g580 ( .A(n_35), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_36), .A2(n_127), .B1(n_303), .B2(n_593), .Y(n_1028) );
INVx1_ASAP7_75t_L g1052 ( .A(n_36), .Y(n_1052) );
INVxp33_ASAP7_75t_SL g982 ( .A(n_37), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_38), .A2(n_79), .B1(n_385), .B2(n_663), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_38), .A2(n_79), .B1(n_347), .B2(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g1394 ( .A(n_39), .Y(n_1394) );
INVx1_ASAP7_75t_L g1227 ( .A(n_40), .Y(n_1227) );
INVxp67_ASAP7_75t_L g1403 ( .A(n_41), .Y(n_1403) );
INVx1_ASAP7_75t_L g737 ( .A(n_42), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_42), .A2(n_133), .B1(n_303), .B2(n_455), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_43), .A2(n_144), .B1(n_619), .B2(n_729), .Y(n_728) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_43), .A2(n_144), .B1(n_477), .B2(n_482), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_44), .A2(n_47), .B1(n_605), .B2(n_882), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_44), .A2(n_64), .B1(n_563), .B2(n_641), .Y(n_932) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_45), .Y(n_480) );
INVx1_ASAP7_75t_L g1076 ( .A(n_46), .Y(n_1076) );
OAI221xp5_ASAP7_75t_L g1094 ( .A1(n_46), .A2(n_78), .B1(n_619), .B2(n_729), .C(n_1095), .Y(n_1094) );
INVxp67_ASAP7_75t_SL g930 ( .A(n_47), .Y(n_930) );
AOI221xp5_ASAP7_75t_L g1352 ( .A1(n_48), .A2(n_67), .B1(n_404), .B2(n_673), .C(n_727), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_48), .A2(n_67), .B1(n_1069), .B2(n_1359), .Y(n_1358) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_49), .A2(n_90), .B1(n_1113), .B2(n_1121), .Y(n_1131) );
INVx1_ASAP7_75t_L g657 ( .A(n_50), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g685 ( .A1(n_50), .A2(n_326), .B(n_686), .Y(n_685) );
OAI22xp33_ASAP7_75t_L g1031 ( .A1(n_51), .A2(n_165), .B1(n_341), .B2(n_347), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_51), .A2(n_243), .B1(n_1040), .B2(n_1044), .Y(n_1043) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_52), .A2(n_100), .B1(n_557), .B2(n_563), .Y(n_763) );
INVx1_ASAP7_75t_L g899 ( .A(n_53), .Y(n_899) );
INVx1_ASAP7_75t_L g721 ( .A(n_54), .Y(n_721) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_55), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_56), .A2(n_177), .B1(n_582), .B2(n_583), .Y(n_581) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_56), .Y(n_630) );
INVx1_ASAP7_75t_L g802 ( .A(n_57), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_58), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_59), .A2(n_180), .B1(n_468), .B2(n_469), .Y(n_467) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_59), .A2(n_246), .B1(n_492), .B2(n_498), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g1382 ( .A1(n_60), .A2(n_1383), .B1(n_1384), .B2(n_1440), .Y(n_1382) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_60), .Y(n_1383) );
INVx1_ASAP7_75t_L g1086 ( .A(n_61), .Y(n_1086) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_63), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g884 ( .A1(n_64), .A2(n_173), .B1(n_531), .B2(n_885), .C(n_887), .Y(n_884) );
INVxp33_ASAP7_75t_SL g790 ( .A(n_65), .Y(n_790) );
AOI221xp5_ASAP7_75t_L g817 ( .A1(n_65), .A2(n_88), .B1(n_325), .B2(n_818), .C(n_820), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_66), .A2(n_102), .B1(n_1113), .B2(n_1121), .Y(n_1176) );
INVxp33_ASAP7_75t_SL g969 ( .A(n_69), .Y(n_969) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_69), .A2(n_105), .B1(n_995), .B2(n_1002), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_70), .A2(n_214), .B1(n_299), .B2(n_302), .Y(n_298) );
INVx1_ASAP7_75t_L g382 ( .A(n_70), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_71), .Y(n_659) );
INVxp33_ASAP7_75t_L g775 ( .A(n_72), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g812 ( .A1(n_72), .A2(n_248), .B1(n_302), .B2(n_813), .C(n_814), .Y(n_812) );
AOI221xp5_ASAP7_75t_L g1430 ( .A1(n_73), .A2(n_135), .B1(n_282), .B2(n_293), .C(n_1431), .Y(n_1430) );
AOI221xp5_ASAP7_75t_L g1342 ( .A1(n_74), .A2(n_92), .B1(n_531), .B2(n_1092), .C(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1364 ( .A(n_74), .Y(n_1364) );
INVx1_ASAP7_75t_L g297 ( .A(n_75), .Y(n_297) );
INVx1_ASAP7_75t_L g309 ( .A(n_75), .Y(n_309) );
INVxp33_ASAP7_75t_L g970 ( .A(n_76), .Y(n_970) );
AOI22xp33_ASAP7_75t_SL g999 ( .A1(n_76), .A2(n_188), .B1(n_384), .B2(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1093 ( .A(n_77), .Y(n_1093) );
INVx1_ASAP7_75t_L g1075 ( .A(n_78), .Y(n_1075) );
INVx1_ASAP7_75t_L g1019 ( .A(n_80), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_80), .A2(n_142), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_81), .A2(n_122), .B1(n_302), .B2(n_592), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_81), .A2(n_122), .B1(n_492), .B2(n_548), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g674 ( .A1(n_82), .A2(n_139), .B1(n_351), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_82), .A2(n_191), .B1(n_300), .B2(n_692), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_83), .A2(n_224), .B1(n_950), .B2(n_952), .Y(n_949) );
INVxp67_ASAP7_75t_SL g974 ( .A(n_83), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_84), .A2(n_191), .B1(n_669), .B2(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g694 ( .A(n_84), .Y(n_694) );
INVx1_ASAP7_75t_L g901 ( .A(n_85), .Y(n_901) );
AOI221xp5_ASAP7_75t_L g907 ( .A1(n_85), .A2(n_239), .B1(n_908), .B2(n_910), .C(n_912), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_86), .A2(n_187), .B1(n_1113), .B2(n_1121), .Y(n_1112) );
AOI22xp5_ASAP7_75t_L g1151 ( .A1(n_87), .A2(n_108), .B1(n_1113), .B2(n_1121), .Y(n_1151) );
INVxp67_ASAP7_75t_SL g793 ( .A(n_88), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_89), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_90), .A2(n_1010), .B1(n_1054), .B2(n_1055), .Y(n_1009) );
INVxp67_ASAP7_75t_SL g1054 ( .A(n_90), .Y(n_1054) );
AOI22xp5_ASAP7_75t_L g1132 ( .A1(n_91), .A2(n_119), .B1(n_1125), .B2(n_1129), .Y(n_1132) );
INVx1_ASAP7_75t_L g1366 ( .A(n_92), .Y(n_1366) );
INVx1_ASAP7_75t_L g1146 ( .A(n_93), .Y(n_1146) );
INVxp67_ASAP7_75t_L g1392 ( .A(n_94), .Y(n_1392) );
AOI221xp5_ASAP7_75t_L g1421 ( .A1(n_94), .A2(n_157), .B1(n_686), .B2(n_1422), .C(n_1423), .Y(n_1421) );
AOI22xp33_ASAP7_75t_SL g1067 ( .A1(n_95), .A2(n_148), .B1(n_282), .B2(n_917), .Y(n_1067) );
AOI21xp33_ASAP7_75t_L g1084 ( .A1(n_95), .A2(n_404), .B(n_539), .Y(n_1084) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_97), .A2(n_204), .B1(n_289), .B2(n_325), .C(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g422 ( .A(n_97), .Y(n_422) );
INVx1_ASAP7_75t_L g1348 ( .A(n_98), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g1361 ( .A1(n_98), .A2(n_217), .B1(n_303), .B2(n_593), .Y(n_1361) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_99), .A2(n_201), .B1(n_663), .B2(n_1090), .Y(n_1353) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_99), .A2(n_201), .B1(n_457), .B2(n_593), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_100), .A2(n_114), .B1(n_724), .B2(n_725), .Y(n_723) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_101), .A2(n_216), .B1(n_477), .B2(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g617 ( .A(n_101), .Y(n_617) );
INVx1_ASAP7_75t_L g255 ( .A(n_103), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_104), .Y(n_852) );
INVxp67_ASAP7_75t_SL g964 ( .A(n_105), .Y(n_964) );
AO22x1_ASAP7_75t_SL g1142 ( .A1(n_106), .A2(n_195), .B1(n_1113), .B2(n_1121), .Y(n_1142) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_107), .Y(n_348) );
XOR2x2_ASAP7_75t_L g568 ( .A(n_109), .B(n_569), .Y(n_568) );
OA22x2_ASAP7_75t_L g273 ( .A1(n_110), .A2(n_274), .B1(n_442), .B2(n_443), .Y(n_273) );
INVx1_ASAP7_75t_L g443 ( .A(n_110), .Y(n_443) );
INVx1_ASAP7_75t_L g588 ( .A(n_111), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g620 ( .A1(n_111), .A2(n_545), .B1(n_621), .B2(n_627), .C(n_632), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_112), .Y(n_938) );
AO221x2_ASAP7_75t_L g1156 ( .A1(n_113), .A2(n_235), .B1(n_1145), .B2(n_1157), .C(n_1158), .Y(n_1156) );
INVx1_ASAP7_75t_L g761 ( .A(n_114), .Y(n_761) );
INVx1_ASAP7_75t_L g1225 ( .A(n_115), .Y(n_1225) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_116), .A2(n_206), .B1(n_1090), .B2(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1367 ( .A(n_116), .Y(n_1367) );
XOR2xp5_ASAP7_75t_L g649 ( .A(n_117), .B(n_650), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_118), .A2(n_174), .B1(n_609), .B2(n_610), .C(n_612), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_118), .A2(n_159), .B1(n_563), .B2(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g805 ( .A(n_120), .Y(n_805) );
INVx1_ASAP7_75t_L g905 ( .A(n_121), .Y(n_905) );
OAI222xp33_ASAP7_75t_L g1387 ( .A1(n_123), .A2(n_151), .B1(n_240), .B2(n_351), .C1(n_1388), .C2(n_1389), .Y(n_1387) );
INVx1_ASAP7_75t_L g1414 ( .A(n_123), .Y(n_1414) );
INVx1_ASAP7_75t_L g603 ( .A(n_124), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_124), .A2(n_174), .B1(n_643), .B2(n_645), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_125), .A2(n_198), .B1(n_619), .B2(n_729), .Y(n_1346) );
INVx1_ASAP7_75t_L g1370 ( .A(n_125), .Y(n_1370) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_126), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_127), .A2(n_230), .B1(n_671), .B2(n_675), .Y(n_1053) );
CKINVDCx5p33_ASAP7_75t_R g1025 ( .A(n_128), .Y(n_1025) );
XNOR2xp5_ASAP7_75t_L g1059 ( .A(n_129), .B(n_1060), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_130), .A2(n_228), .B1(n_454), .B2(n_456), .Y(n_453) );
INVx1_ASAP7_75t_L g507 ( .A(n_130), .Y(n_507) );
INVx1_ASAP7_75t_L g797 ( .A(n_131), .Y(n_797) );
AOI221xp5_ASAP7_75t_L g845 ( .A1(n_132), .A2(n_242), .B1(n_686), .B2(n_820), .C(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g868 ( .A(n_132), .Y(n_868) );
INVx1_ASAP7_75t_L g735 ( .A(n_133), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g1124 ( .A1(n_134), .A2(n_231), .B1(n_1125), .B2(n_1129), .Y(n_1124) );
INVx1_ASAP7_75t_L g1371 ( .A(n_134), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_134), .A2(n_1377), .B1(n_1381), .B2(n_1441), .Y(n_1376) );
OAI332xp33_ASAP7_75t_L g1390 ( .A1(n_135), .A2(n_403), .A3(n_1391), .B1(n_1395), .B2(n_1398), .B3(n_1404), .C1(n_1407), .C2(n_1408), .Y(n_1390) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_136), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_137), .A2(n_160), .B1(n_619), .B2(n_729), .Y(n_889) );
OAI221xp5_ASAP7_75t_L g924 ( .A1(n_137), .A2(n_160), .B1(n_925), .B2(n_927), .C(n_928), .Y(n_924) );
INVx1_ASAP7_75t_L g701 ( .A(n_139), .Y(n_701) );
XNOR2xp5_ASAP7_75t_L g830 ( .A(n_140), .B(n_831), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_141), .Y(n_529) );
INVx1_ASAP7_75t_L g1015 ( .A(n_142), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_143), .A2(n_209), .B1(n_725), .B2(n_1090), .Y(n_1089) );
AOI22xp33_ASAP7_75t_SL g1070 ( .A1(n_145), .A2(n_156), .B1(n_457), .B2(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1079 ( .A(n_145), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_146), .A2(n_246), .B1(n_460), .B2(n_463), .Y(n_466) );
OAI22xp33_ASAP7_75t_L g544 ( .A1(n_146), .A2(n_180), .B1(n_545), .B2(n_548), .Y(n_544) );
INVx1_ASAP7_75t_L g684 ( .A(n_147), .Y(n_684) );
INVx1_ASAP7_75t_L g1083 ( .A(n_148), .Y(n_1083) );
AOI21xp33_ASAP7_75t_L g1020 ( .A1(n_149), .A2(n_326), .B(n_455), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_149), .A2(n_229), .B1(n_1040), .B2(n_1042), .Y(n_1039) );
INVxp33_ASAP7_75t_L g788 ( .A(n_150), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_150), .A2(n_178), .B1(n_823), .B2(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g1427 ( .A(n_151), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_152), .A2(n_215), .B1(n_1129), .B2(n_1145), .Y(n_1177) );
INVx1_ASAP7_75t_L g827 ( .A(n_153), .Y(n_827) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_154), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_154), .B(n_255), .Y(n_1120) );
AND3x2_ASAP7_75t_L g1126 ( .A(n_154), .B(n_255), .C(n_1117), .Y(n_1126) );
OAI22xp33_ASAP7_75t_SL g836 ( .A1(n_155), .A2(n_169), .B1(n_811), .B2(n_837), .Y(n_836) );
OAI221xp5_ASAP7_75t_L g862 ( .A1(n_155), .A2(n_169), .B1(n_396), .B2(n_783), .C(n_785), .Y(n_862) );
INVx1_ASAP7_75t_L g1080 ( .A(n_156), .Y(n_1080) );
INVx1_ASAP7_75t_L g1396 ( .A(n_157), .Y(n_1396) );
AOI221xp5_ASAP7_75t_L g941 ( .A1(n_158), .A2(n_221), .B1(n_463), .B2(n_942), .C(n_943), .Y(n_941) );
INVxp33_ASAP7_75t_SL g984 ( .A(n_158), .Y(n_984) );
INVx1_ASAP7_75t_L g607 ( .A(n_159), .Y(n_607) );
INVx2_ASAP7_75t_L g268 ( .A(n_161), .Y(n_268) );
AOI22xp33_ASAP7_75t_SL g992 ( .A1(n_162), .A2(n_194), .B1(n_993), .B2(n_995), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_163), .A2(n_223), .B1(n_282), .B2(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g410 ( .A(n_163), .Y(n_410) );
INVx1_ASAP7_75t_L g858 ( .A(n_164), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_166), .Y(n_335) );
OAI211xp5_ASAP7_75t_L g718 ( .A1(n_167), .A2(n_498), .B(n_719), .C(n_722), .Y(n_718) );
INVx1_ASAP7_75t_L g758 ( .A(n_167), .Y(n_758) );
INVx1_ASAP7_75t_L g1148 ( .A(n_168), .Y(n_1148) );
CKINVDCx5p33_ASAP7_75t_R g1024 ( .A(n_170), .Y(n_1024) );
INVx1_ASAP7_75t_L g897 ( .A(n_171), .Y(n_897) );
INVx1_ASAP7_75t_L g1117 ( .A(n_172), .Y(n_1117) );
INVxp67_ASAP7_75t_SL g931 ( .A(n_173), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_175), .A2(n_238), .B1(n_539), .B2(n_611), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_175), .A2(n_238), .B1(n_341), .B2(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_176), .A2(n_219), .B1(n_460), .B2(n_463), .Y(n_459) );
INVx1_ASAP7_75t_L g514 ( .A(n_176), .Y(n_514) );
INVxp67_ASAP7_75t_SL g628 ( .A(n_177), .Y(n_628) );
INVxp67_ASAP7_75t_SL g794 ( .A(n_178), .Y(n_794) );
OAI211xp5_ASAP7_75t_L g879 ( .A1(n_179), .A2(n_498), .B(n_880), .C(n_890), .Y(n_879) );
AOI221xp5_ASAP7_75t_L g914 ( .A1(n_179), .A2(n_185), .B1(n_460), .B2(n_915), .C(n_918), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g934 ( .A(n_181), .Y(n_934) );
INVx1_ASAP7_75t_L g270 ( .A(n_182), .Y(n_270) );
INVx2_ASAP7_75t_L g370 ( .A(n_182), .Y(n_370) );
INVx1_ASAP7_75t_L g891 ( .A(n_183), .Y(n_891) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_184), .B(n_350), .Y(n_1011) );
OAI221xp5_ASAP7_75t_L g893 ( .A1(n_185), .A2(n_545), .B1(n_632), .B2(n_894), .C(n_900), .Y(n_893) );
INVx1_ASAP7_75t_L g746 ( .A(n_186), .Y(n_746) );
INVxp67_ASAP7_75t_SL g948 ( .A(n_188), .Y(n_948) );
INVx1_ASAP7_75t_L g800 ( .A(n_189), .Y(n_800) );
AOI221xp5_ASAP7_75t_L g1221 ( .A1(n_190), .A2(n_192), .B1(n_1222), .B2(n_1223), .C(n_1224), .Y(n_1221) );
NOR2xp33_ASAP7_75t_L g1336 ( .A(n_193), .B(n_1337), .Y(n_1336) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_196), .Y(n_844) );
INVx1_ASAP7_75t_L g779 ( .A(n_197), .Y(n_779) );
INVx1_ASAP7_75t_L g1369 ( .A(n_198), .Y(n_1369) );
INVx1_ASAP7_75t_L g576 ( .A(n_199), .Y(n_576) );
INVx1_ASAP7_75t_L g540 ( .A(n_200), .Y(n_540) );
INVx1_ASAP7_75t_L g770 ( .A(n_202), .Y(n_770) );
XOR2xp5_ASAP7_75t_L g446 ( .A(n_203), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g416 ( .A(n_204), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_205), .Y(n_310) );
INVx1_ASAP7_75t_L g1363 ( .A(n_206), .Y(n_1363) );
INVx1_ASAP7_75t_L g524 ( .A(n_207), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_208), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_210), .A2(n_213), .B1(n_312), .B2(n_319), .Y(n_311) );
OAI221xp5_ASAP7_75t_L g389 ( .A1(n_210), .A2(n_213), .B1(n_390), .B2(n_396), .C(n_400), .Y(n_389) );
INVx1_ASAP7_75t_L g1118 ( .A(n_211), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_211), .B(n_1116), .Y(n_1123) );
INVx1_ASAP7_75t_L g1416 ( .A(n_212), .Y(n_1416) );
INVx1_ASAP7_75t_L g361 ( .A(n_214), .Y(n_361) );
INVx1_ASAP7_75t_L g614 ( .A(n_216), .Y(n_614) );
INVx1_ASAP7_75t_L g1349 ( .A(n_217), .Y(n_1349) );
INVx1_ASAP7_75t_L g1397 ( .A(n_218), .Y(n_1397) );
INVx1_ASAP7_75t_L g512 ( .A(n_219), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_220), .Y(n_841) );
INVxp33_ASAP7_75t_L g986 ( .A(n_221), .Y(n_986) );
INVx1_ASAP7_75t_L g865 ( .A(n_222), .Y(n_865) );
INVx1_ASAP7_75t_L g425 ( .A(n_223), .Y(n_425) );
INVxp67_ASAP7_75t_SL g978 ( .A(n_224), .Y(n_978) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_225), .Y(n_742) );
INVx2_ASAP7_75t_L g267 ( .A(n_226), .Y(n_267) );
INVx1_ASAP7_75t_L g590 ( .A(n_227), .Y(n_590) );
OAI211xp5_ASAP7_75t_SL g598 ( .A1(n_227), .A2(n_498), .B(n_599), .C(n_613), .Y(n_598) );
INVx1_ASAP7_75t_L g503 ( .A(n_228), .Y(n_503) );
INVx1_ASAP7_75t_L g1017 ( .A(n_229), .Y(n_1017) );
INVx1_ASAP7_75t_L g1027 ( .A(n_230), .Y(n_1027) );
INVx1_ASAP7_75t_L g892 ( .A(n_232), .Y(n_892) );
INVx1_ASAP7_75t_L g371 ( .A(n_233), .Y(n_371) );
INVx1_ASAP7_75t_L g777 ( .A(n_234), .Y(n_777) );
INVx1_ASAP7_75t_L g854 ( .A(n_236), .Y(n_854) );
INVx1_ASAP7_75t_L g1345 ( .A(n_237), .Y(n_1345) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_237), .A2(n_247), .B1(n_461), .B2(n_917), .Y(n_1360) );
AOI21xp33_ASAP7_75t_L g902 ( .A1(n_239), .A2(n_404), .B(n_885), .Y(n_902) );
INVx1_ASAP7_75t_L g1417 ( .A(n_240), .Y(n_1417) );
INVxp67_ASAP7_75t_L g1399 ( .A(n_241), .Y(n_1399) );
INVx1_ASAP7_75t_L g866 ( .A(n_242), .Y(n_866) );
OAI211xp5_ASAP7_75t_SL g1022 ( .A1(n_243), .A2(n_679), .B(n_1023), .C(n_1026), .Y(n_1022) );
BUFx3_ASAP7_75t_L g286 ( .A(n_244), .Y(n_286) );
INVx1_ASAP7_75t_L g305 ( .A(n_244), .Y(n_305) );
BUFx3_ASAP7_75t_L g288 ( .A(n_245), .Y(n_288) );
INVx1_ASAP7_75t_L g301 ( .A(n_245), .Y(n_301) );
INVx1_ASAP7_75t_L g1351 ( .A(n_247), .Y(n_1351) );
INVxp33_ASAP7_75t_L g780 ( .A(n_248), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_271), .B(n_1105), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_258), .Y(n_252) );
AND2x4_ASAP7_75t_L g1375 ( .A(n_253), .B(n_259), .Y(n_1375) );
NOR2xp33_ASAP7_75t_SL g253 ( .A(n_254), .B(n_256), .Y(n_253) );
INVx1_ASAP7_75t_SL g1380 ( .A(n_254), .Y(n_1380) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_254), .B(n_256), .Y(n_1446) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_256), .B(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_264), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g517 ( .A(n_262), .B(n_270), .Y(n_517) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g404 ( .A(n_263), .B(n_405), .Y(n_404) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .Y(n_264) );
OR2x2_ASAP7_75t_L g351 ( .A(n_265), .B(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g409 ( .A(n_265), .Y(n_409) );
INVx1_ASAP7_75t_L g528 ( .A(n_265), .Y(n_528) );
INVx2_ASAP7_75t_SL g625 ( .A(n_265), .Y(n_625) );
INVx2_ASAP7_75t_SL g741 ( .A(n_265), .Y(n_741) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_265), .Y(n_874) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
AND2x4_ASAP7_75t_L g365 ( .A(n_267), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g375 ( .A(n_267), .Y(n_375) );
AND2x2_ASAP7_75t_L g381 ( .A(n_267), .B(n_268), .Y(n_381) );
INVx2_ASAP7_75t_L g386 ( .A(n_267), .Y(n_386) );
INVx1_ASAP7_75t_L g415 ( .A(n_267), .Y(n_415) );
INVx2_ASAP7_75t_L g366 ( .A(n_268), .Y(n_366) );
INVx1_ASAP7_75t_L g388 ( .A(n_268), .Y(n_388) );
INVx1_ASAP7_75t_L g394 ( .A(n_268), .Y(n_394) );
INVx1_ASAP7_75t_L g414 ( .A(n_268), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_268), .B(n_386), .Y(n_421) );
INVx2_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
XNOR2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_711), .Y(n_271) );
OAI22xp33_ASAP7_75t_SL g272 ( .A1(n_273), .A2(n_444), .B1(n_709), .B2(n_710), .Y(n_272) );
INVx3_ASAP7_75t_L g709 ( .A(n_273), .Y(n_709) );
INVx1_ASAP7_75t_L g442 ( .A(n_274), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_358), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_279), .B1(n_348), .B2(n_349), .Y(n_275) );
INVx2_ASAP7_75t_L g634 ( .A(n_276), .Y(n_634) );
NOR2xp67_ASAP7_75t_L g638 ( .A(n_276), .B(n_535), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g832 ( .A1(n_276), .A2(n_828), .B1(n_833), .B2(n_854), .Y(n_832) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x6_ASAP7_75t_L g451 ( .A(n_277), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g665 ( .A(n_277), .B(n_532), .Y(n_665) );
OR2x2_ASAP7_75t_L g750 ( .A(n_277), .B(n_751), .Y(n_750) );
BUFx2_ASAP7_75t_L g903 ( .A(n_277), .Y(n_903) );
AND2x4_ASAP7_75t_L g991 ( .A(n_277), .B(n_517), .Y(n_991) );
AND2x4_ASAP7_75t_L g1035 ( .A(n_277), .B(n_517), .Y(n_1035) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x6_ASAP7_75t_L g403 ( .A(n_278), .B(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g551 ( .A(n_278), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_323), .C(n_338), .Y(n_279) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_298), .B1(n_306), .B2(n_310), .C(n_311), .Y(n_280) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g698 ( .A(n_283), .Y(n_698) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_283), .Y(n_849) );
INVx2_ASAP7_75t_L g911 ( .A(n_283), .Y(n_911) );
INVx6_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g357 ( .A(n_284), .B(n_314), .Y(n_357) );
INVx2_ASAP7_75t_L g462 ( .A(n_284), .Y(n_462) );
BUFx2_ASAP7_75t_L g1359 ( .A(n_284), .Y(n_1359) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_L g322 ( .A(n_285), .Y(n_322) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g292 ( .A(n_286), .B(n_288), .Y(n_292) );
AND2x4_ASAP7_75t_L g300 ( .A(n_286), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g318 ( .A(n_287), .Y(n_318) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g304 ( .A(n_288), .B(n_305), .Y(n_304) );
INVx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g1069 ( .A(n_290), .Y(n_1069) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_291), .Y(n_465) );
INVx1_ASAP7_75t_L g488 ( .A(n_291), .Y(n_488) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_292), .Y(n_334) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g474 ( .A(n_294), .B(n_356), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g699 ( .A(n_294), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g814 ( .A1(n_294), .A2(n_644), .B1(n_703), .B2(n_777), .C(n_779), .Y(n_814) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_294), .A2(n_644), .B1(n_703), .B2(n_841), .C(n_842), .Y(n_840) );
INVx2_ASAP7_75t_L g944 ( .A(n_294), .Y(n_944) );
INVx2_ASAP7_75t_SL g1030 ( .A(n_294), .Y(n_1030) );
AND2x4_ASAP7_75t_L g1072 ( .A(n_294), .B(n_356), .Y(n_1072) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
AND2x4_ASAP7_75t_L g314 ( .A(n_295), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g327 ( .A(n_296), .B(n_297), .Y(n_327) );
AND2x2_ASAP7_75t_L g306 ( .A(n_299), .B(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g582 ( .A(n_299), .Y(n_582) );
INVx1_ASAP7_75t_L g646 ( .A(n_299), .Y(n_646) );
BUFx4f_ASAP7_75t_L g920 ( .A(n_299), .Y(n_920) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx2_ASAP7_75t_L g325 ( .A(n_300), .Y(n_325) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_300), .Y(n_455) );
INVx2_ASAP7_75t_SL g561 ( .A(n_300), .Y(n_561) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_300), .Y(n_593) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_300), .Y(n_686) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_300), .Y(n_839) );
BUFx3_ASAP7_75t_L g1071 ( .A(n_300), .Y(n_1071) );
INVx1_ASAP7_75t_L g344 ( .A(n_301), .Y(n_344) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g1016 ( .A(n_303), .Y(n_1016) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g332 ( .A(n_304), .Y(n_332) );
INVx1_ASAP7_75t_L g458 ( .A(n_304), .Y(n_458) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_304), .Y(n_471) );
INVx1_ASAP7_75t_L g584 ( .A(n_304), .Y(n_584) );
INVx1_ASAP7_75t_L g343 ( .A(n_305), .Y(n_343) );
INVx1_ASAP7_75t_L g679 ( .A(n_306), .Y(n_679) );
AND2x4_ASAP7_75t_L g333 ( .A(n_307), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g809 ( .A(n_307), .B(n_593), .Y(n_809) );
AOI221xp5_ASAP7_75t_L g1418 ( .A1(n_307), .A2(n_333), .B1(n_336), .B2(n_1406), .C(n_1419), .Y(n_1418) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g341 ( .A(n_308), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g347 ( .A(n_308), .B(n_332), .Y(n_347) );
OR2x2_ASAP7_75t_L g555 ( .A(n_308), .B(n_368), .Y(n_555) );
INVx1_ASAP7_75t_L g315 ( .A(n_309), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_310), .A2(n_345), .B1(n_418), .B2(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx4_ASAP7_75t_L g811 ( .A(n_313), .Y(n_811) );
AOI22xp5_ASAP7_75t_L g1023 ( .A1(n_313), .A2(n_320), .B1(n_1024), .B2(n_1025), .Y(n_1023) );
AND2x4_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
AND2x4_ASAP7_75t_L g320 ( .A(n_314), .B(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g337 ( .A(n_314), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g479 ( .A(n_314), .B(n_438), .Y(n_479) );
AND2x4_ASAP7_75t_L g951 ( .A(n_314), .B(n_316), .Y(n_951) );
AND2x2_ASAP7_75t_L g953 ( .A(n_314), .B(n_321), .Y(n_953) );
INVx1_ASAP7_75t_L g967 ( .A(n_314), .Y(n_967) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_316), .A2(n_321), .B1(n_705), .B2(n_706), .Y(n_704) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g483 ( .A(n_317), .Y(n_483) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g837 ( .A(n_320), .Y(n_837) );
AOI222xp33_ASAP7_75t_SL g1411 ( .A1(n_320), .A2(n_1412), .B1(n_1414), .B2(n_1415), .C1(n_1416), .C2(n_1417), .Y(n_1411) );
INVx2_ASAP7_75t_L g478 ( .A(n_321), .Y(n_478) );
BUFx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_328), .B1(n_333), .B2(n_335), .C(n_336), .Y(n_323) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g452 ( .A(n_327), .Y(n_452) );
INVx1_ASAP7_75t_L g751 ( .A(n_327), .Y(n_751) );
BUFx3_ASAP7_75t_L g821 ( .A(n_327), .Y(n_821) );
INVx1_ASAP7_75t_L g956 ( .A(n_327), .Y(n_956) );
INVx2_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g850 ( .A(n_330), .Y(n_850) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g692 ( .A(n_332), .Y(n_692) );
INVx2_ASAP7_75t_SL g681 ( .A(n_333), .Y(n_681) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_333), .Y(n_816) );
AOI221xp5_ASAP7_75t_L g843 ( .A1(n_333), .A2(n_336), .B1(n_844), .B2(n_845), .C(n_847), .Y(n_843) );
BUFx6f_ASAP7_75t_L g963 ( .A(n_333), .Y(n_963) );
AND2x4_ASAP7_75t_L g336 ( .A(n_334), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_SL g819 ( .A(n_334), .Y(n_819) );
BUFx6f_ASAP7_75t_L g917 ( .A(n_334), .Y(n_917) );
BUFx4f_ASAP7_75t_L g1422 ( .A(n_334), .Y(n_1422) );
INVx1_ASAP7_75t_L g1432 ( .A(n_334), .Y(n_1432) );
OAI22xp33_ASAP7_75t_L g430 ( .A1(n_335), .A2(n_339), .B1(n_407), .B2(n_431), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g815 ( .A1(n_336), .A2(n_805), .B1(n_816), .B2(n_817), .C(n_822), .Y(n_815) );
INVx1_ASAP7_75t_L g1021 ( .A(n_336), .Y(n_1021) );
BUFx3_ASAP7_75t_L g707 ( .A(n_337), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_345), .B2(n_346), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_340), .A2(n_346), .B1(n_800), .B2(n_802), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_340), .A2(n_346), .B1(n_852), .B2(n_853), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_340), .A2(n_346), .B1(n_969), .B2(n_970), .Y(n_968) );
INVx6_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g575 ( .A(n_342), .Y(n_575) );
INVx2_ASAP7_75t_L g587 ( .A(n_342), .Y(n_587) );
INVx1_ASAP7_75t_L g690 ( .A(n_342), .Y(n_690) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x2_ASAP7_75t_L g565 ( .A(n_343), .B(n_344), .Y(n_565) );
INVx4_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g828 ( .A(n_350), .Y(n_828) );
INVx5_ASAP7_75t_L g937 ( .A(n_350), .Y(n_937) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_354), .Y(n_350) );
INVx3_ASAP7_75t_L g395 ( .A(n_352), .Y(n_395) );
INVx1_ASAP7_75t_L g538 ( .A(n_353), .Y(n_538) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI222xp33_ASAP7_75t_L g552 ( .A1(n_355), .A2(n_524), .B1(n_529), .B2(n_540), .C1(n_553), .C2(n_556), .Y(n_552) );
OR2x6_ASAP7_75t_L g637 ( .A(n_355), .B(n_638), .Y(n_637) );
AND2x4_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx2_ASAP7_75t_L g1413 ( .A(n_357), .Y(n_1413) );
NOR3xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_389), .C(n_402), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_376), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B1(n_371), .B2(n_372), .Y(n_360) );
BUFx2_ASAP7_75t_L g776 ( .A(n_362), .Y(n_776) );
BUFx2_ASAP7_75t_L g859 ( .A(n_362), .Y(n_859) );
BUFx2_ASAP7_75t_L g983 ( .A(n_362), .Y(n_983) );
BUFx2_ASAP7_75t_L g1438 ( .A(n_362), .Y(n_1438) );
AND2x4_ASAP7_75t_L g362 ( .A(n_363), .B(n_367), .Y(n_362) );
INVx1_ASAP7_75t_SL g658 ( .A(n_363), .Y(n_658) );
INVx1_ASAP7_75t_L g736 ( .A(n_363), .Y(n_736) );
INVx2_ASAP7_75t_L g898 ( .A(n_363), .Y(n_898) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g424 ( .A(n_364), .Y(n_424) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_364), .Y(n_523) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g497 ( .A(n_365), .Y(n_497) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_365), .Y(n_509) );
AND2x4_ASAP7_75t_L g374 ( .A(n_366), .B(n_375), .Y(n_374) );
AND2x6_ASAP7_75t_L g372 ( .A(n_367), .B(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g378 ( .A(n_367), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g383 ( .A(n_367), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g654 ( .A(n_367), .B(n_539), .Y(n_654) );
AND2x2_ASAP7_75t_L g670 ( .A(n_367), .B(n_384), .Y(n_670) );
AND2x2_ASAP7_75t_L g672 ( .A(n_367), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g676 ( .A(n_367), .B(n_424), .Y(n_676) );
AND2x2_ASAP7_75t_L g781 ( .A(n_367), .B(n_384), .Y(n_781) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_367), .B(n_384), .Y(n_1051) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g438 ( .A(n_368), .Y(n_438) );
INVx2_ASAP7_75t_L g495 ( .A(n_369), .Y(n_495) );
AND2x4_ASAP7_75t_L g546 ( .A(n_369), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g549 ( .A(n_369), .B(n_385), .Y(n_549) );
INVx1_ASAP7_75t_L g405 ( .A(n_370), .Y(n_405) );
INVx1_ASAP7_75t_L g440 ( .A(n_370), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_372), .A2(n_775), .B1(n_776), .B2(n_777), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_372), .A2(n_841), .B1(n_858), .B2(n_859), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_372), .A2(n_982), .B1(n_983), .B2(n_984), .Y(n_981) );
NAND2x1p5_ASAP7_75t_L g401 ( .A(n_373), .B(n_395), .Y(n_401) );
BUFx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx3_ASAP7_75t_L g500 ( .A(n_374), .Y(n_500) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_374), .Y(n_611) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_374), .Y(n_673) );
BUFx2_ASAP7_75t_L g980 ( .A(n_374), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B1(n_382), .B2(n_383), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_378), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_378), .A2(n_383), .B1(n_842), .B2(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_378), .A2(n_781), .B1(n_986), .B2(n_987), .Y(n_985) );
AOI221xp5_ASAP7_75t_L g1049 ( .A1(n_378), .A2(n_1050), .B1(n_1051), .B2(n_1052), .C(n_1053), .Y(n_1049) );
INVx1_ASAP7_75t_L g1436 ( .A(n_378), .Y(n_1436) );
INVx1_ASAP7_75t_L g886 ( .A(n_379), .Y(n_886) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_379), .Y(n_1002) );
BUFx2_ASAP7_75t_L g1037 ( .A(n_379), .Y(n_1037) );
INVx2_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_SL g539 ( .A(n_380), .Y(n_539) );
INVx2_ASAP7_75t_L g1097 ( .A(n_380), .Y(n_1097) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_381), .Y(n_547) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_385), .Y(n_724) );
INVx1_ASAP7_75t_L g883 ( .A(n_385), .Y(n_883) );
INVx1_ASAP7_75t_L g1041 ( .A(n_385), .Y(n_1041) );
BUFx6f_ASAP7_75t_L g1090 ( .A(n_385), .Y(n_1090) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g399 ( .A(n_386), .Y(n_399) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g784 ( .A(n_391), .Y(n_784) );
NAND2x1_ASAP7_75t_SL g391 ( .A(n_392), .B(n_395), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_392), .A2(n_398), .B1(n_480), .B2(n_485), .Y(n_543) );
NAND2x1p5_ASAP7_75t_L g729 ( .A(n_392), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_394), .Y(n_616) );
NAND2x1p5_ASAP7_75t_L g397 ( .A(n_395), .B(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g973 ( .A(n_395), .B(n_616), .Y(n_973) );
AND2x4_ASAP7_75t_L g975 ( .A(n_395), .B(n_976), .Y(n_975) );
AND2x4_ASAP7_75t_L g979 ( .A(n_395), .B(n_980), .Y(n_979) );
BUFx4f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx4f_ASAP7_75t_L g1389 ( .A(n_397), .Y(n_1389) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OR2x6_ASAP7_75t_L g619 ( .A(n_399), .B(n_537), .Y(n_619) );
BUFx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g785 ( .A(n_401), .Y(n_785) );
OAI33xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_406), .A3(n_417), .B1(n_426), .B2(n_430), .B3(n_435), .Y(n_402) );
OAI33xp33_ASAP7_75t_L g786 ( .A1(n_403), .A2(n_435), .A3(n_787), .B1(n_792), .B2(n_795), .B3(n_801), .Y(n_786) );
OAI33xp33_ASAP7_75t_L g863 ( .A1(n_403), .A2(n_435), .A3(n_864), .B1(n_867), .B2(n_870), .B3(n_873), .Y(n_863) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_410), .B1(n_411), .B2(n_416), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g513 ( .A(n_408), .Y(n_513) );
INVx1_ASAP7_75t_L g789 ( .A(n_408), .Y(n_789) );
INVx2_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_411), .A2(n_789), .B1(n_865), .B2(n_866), .Y(n_864) );
BUFx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI221xp5_ASAP7_75t_L g525 ( .A1(n_412), .A2(n_526), .B1(n_527), .B2(n_529), .C(n_530), .Y(n_525) );
INVx2_ASAP7_75t_L g804 ( .A(n_412), .Y(n_804) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
AND2x2_ASAP7_75t_L g434 ( .A(n_414), .B(n_415), .Y(n_434) );
INVx1_ASAP7_75t_L g977 ( .A(n_415), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_422), .B1(n_423), .B2(n_425), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_418), .A2(n_521), .B1(n_793), .B2(n_794), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_418), .A2(n_521), .B1(n_868), .B2(n_869), .Y(n_867) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g656 ( .A(n_420), .Y(n_656) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_420), .Y(n_896) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g506 ( .A(n_421), .Y(n_506) );
BUFx2_ASAP7_75t_L g734 ( .A(n_421), .Y(n_734) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g429 ( .A(n_424), .Y(n_429) );
INVx2_ASAP7_75t_L g606 ( .A(n_424), .Y(n_606) );
HB1xp67_ASAP7_75t_L g1341 ( .A(n_424), .Y(n_1341) );
INVx1_ASAP7_75t_L g1402 ( .A(n_424), .Y(n_1402) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g799 ( .A(n_429), .Y(n_799) );
INVx1_ASAP7_75t_L g1042 ( .A(n_429), .Y(n_1042) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g632 ( .A(n_433), .B(n_537), .Y(n_632) );
OR2x6_ASAP7_75t_L g743 ( .A(n_433), .B(n_537), .Y(n_743) );
OAI22xp33_ASAP7_75t_L g1395 ( .A1(n_433), .A2(n_740), .B1(n_1396), .B2(n_1397), .Y(n_1395) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g511 ( .A(n_434), .Y(n_511) );
INVx3_ASAP7_75t_L g542 ( .A(n_434), .Y(n_542) );
BUFx2_ASAP7_75t_L g623 ( .A(n_434), .Y(n_623) );
CKINVDCx8_ASAP7_75t_R g435 ( .A(n_436), .Y(n_435) );
INVx5_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx6_ASAP7_75t_L g1003 ( .A(n_437), .Y(n_1003) );
OR2x6_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx2_ASAP7_75t_L g532 ( .A(n_439), .Y(n_532) );
BUFx2_ASAP7_75t_L g612 ( .A(n_439), .Y(n_612) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g710 ( .A(n_444), .Y(n_710) );
XNOR2x1_ASAP7_75t_SL g444 ( .A(n_445), .B(n_566), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND4xp75_ASAP7_75t_L g447 ( .A(n_448), .B(n_490), .C(n_552), .D(n_558), .Y(n_447) );
AND2x2_ASAP7_75t_SL g448 ( .A(n_449), .B(n_475), .Y(n_448) );
AOI33xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_453), .A3(n_459), .B1(n_466), .B2(n_467), .B3(n_472), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_451), .A2(n_473), .B1(n_572), .B2(n_585), .Y(n_571) );
INVx2_ASAP7_75t_L g913 ( .A(n_451), .Y(n_913) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx3_ASAP7_75t_L g468 ( .A(n_455), .Y(n_468) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x6_ASAP7_75t_L g557 ( .A(n_458), .B(n_555), .Y(n_557) );
OR2x2_ASAP7_75t_L g641 ( .A(n_458), .B(n_555), .Y(n_641) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g553 ( .A(n_461), .B(n_554), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g700 ( .A1(n_461), .A2(n_701), .B(n_702), .C(n_707), .Y(n_700) );
INVx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g909 ( .A(n_465), .Y(n_909) );
AND2x4_ASAP7_75t_L g965 ( .A(n_465), .B(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g825 ( .A(n_471), .Y(n_825) );
INVx1_ASAP7_75t_L g923 ( .A(n_471), .Y(n_923) );
BUFx6f_ASAP7_75t_L g962 ( .A(n_471), .Y(n_962) );
BUFx6f_ASAP7_75t_L g1066 ( .A(n_471), .Y(n_1066) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_473), .A2(n_750), .B1(n_752), .B2(n_756), .Y(n_749) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g906 ( .A1(n_474), .A2(n_907), .B1(n_913), .B2(n_914), .C(n_924), .Y(n_906) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_480), .B1(n_481), .B2(n_485), .C(n_486), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g1073 ( .A1(n_476), .A2(n_486), .B1(n_1074), .B2(n_1075), .C(n_1076), .Y(n_1073) );
AOI221xp5_ASAP7_75t_L g1368 ( .A1(n_476), .A2(n_486), .B1(n_1074), .B2(n_1369), .C(n_1370), .Y(n_1368) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
OR2x2_ASAP7_75t_L g927 ( .A(n_478), .B(n_479), .Y(n_927) );
INVx2_ASAP7_75t_SL g484 ( .A(n_479), .Y(n_484) );
INVx1_ASAP7_75t_L g489 ( .A(n_479), .Y(n_489) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_482), .Y(n_596) );
INVx2_ASAP7_75t_L g926 ( .A(n_482), .Y(n_926) );
INVx2_ASAP7_75t_L g1074 ( .A(n_482), .Y(n_1074) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
BUFx2_ASAP7_75t_L g594 ( .A(n_486), .Y(n_594) );
NOR3xp33_ASAP7_75t_L g747 ( .A(n_486), .B(n_748), .C(n_749), .Y(n_747) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_489), .B(n_917), .Y(n_928) );
OAI31xp33_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_501), .A3(n_544), .B(n_550), .Y(n_490) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_493), .A2(n_549), .B1(n_720), .B2(n_721), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_493), .A2(n_549), .B1(n_891), .B2(n_892), .Y(n_890) );
AOI221x1_ASAP7_75t_L g1078 ( .A1(n_493), .A2(n_549), .B1(n_1079), .B2(n_1080), .C(n_1081), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_493), .A2(n_549), .B1(n_1348), .B2(n_1349), .Y(n_1347) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
AND2x4_ASAP7_75t_L g499 ( .A(n_494), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g1045 ( .A(n_496), .Y(n_1045) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g663 ( .A(n_497), .Y(n_663) );
INVx8_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AOI221xp5_ASAP7_75t_SL g1088 ( .A1(n_499), .A2(n_1089), .B1(n_1091), .B2(n_1093), .C(n_1094), .Y(n_1088) );
AOI221xp5_ASAP7_75t_SL g1339 ( .A1(n_499), .A2(n_1340), .B1(n_1342), .B2(n_1345), .C(n_1346), .Y(n_1339) );
BUFx6f_ASAP7_75t_L g1038 ( .A(n_500), .Y(n_1038) );
INVx1_ASAP7_75t_L g1344 ( .A(n_500), .Y(n_1344) );
OAI221xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_510), .B1(n_518), .B2(n_525), .C(n_533), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B1(n_507), .B2(n_508), .Y(n_502) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g519 ( .A(n_505), .Y(n_519) );
INVx2_ASAP7_75t_L g1393 ( .A(n_505), .Y(n_1393) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g602 ( .A(n_506), .Y(n_602) );
INVx2_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_SL g631 ( .A(n_509), .Y(n_631) );
INVx4_ASAP7_75t_L g872 ( .A(n_509), .Y(n_872) );
BUFx3_ASAP7_75t_L g998 ( .A(n_509), .Y(n_998) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_513), .B2(n_514), .C(n_515), .Y(n_510) );
OAI22xp33_ASAP7_75t_L g873 ( .A1(n_511), .A2(n_844), .B1(n_852), .B2(n_874), .Y(n_873) );
OAI21xp5_ASAP7_75t_SL g900 ( .A1(n_511), .A2(n_901), .B(n_902), .Y(n_900) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_SL g626 ( .A(n_517), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B1(n_521), .B2(n_524), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_520), .A2(n_526), .B1(n_559), .B2(n_562), .Y(n_558) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g725 ( .A(n_523), .Y(n_725) );
OAI22xp5_ASAP7_75t_SL g1404 ( .A1(n_527), .A2(n_803), .B1(n_1405), .B2(n_1406), .Y(n_1404) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_540), .B(n_541), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_539), .Y(n_535) );
AND2x2_ASAP7_75t_L g615 ( .A(n_536), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AOI21xp33_ASAP7_75t_L g541 ( .A1(n_537), .A2(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_L g730 ( .A(n_537), .Y(n_730) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx2_ASAP7_75t_L g609 ( .A(n_539), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g738 ( .A1(n_542), .A2(n_626), .B1(n_739), .B2(n_740), .C(n_742), .Y(n_738) );
OAI21xp5_ASAP7_75t_SL g1082 ( .A1(n_542), .A2(n_1083), .B(n_1084), .Y(n_1082) );
CKINVDCx6p67_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
AOI221xp5_ASAP7_75t_L g1350 ( .A1(n_546), .A2(n_1351), .B1(n_1352), .B2(n_1353), .C(n_1354), .Y(n_1350) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_547), .Y(n_727) );
INVx3_ASAP7_75t_L g994 ( .A(n_547), .Y(n_994) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_547), .Y(n_1092) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g708 ( .A(n_550), .Y(n_708) );
BUFx8_ASAP7_75t_SL g744 ( .A(n_550), .Y(n_744) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx2_ASAP7_75t_L g1098 ( .A(n_551), .Y(n_1098) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_553), .A2(n_559), .B1(n_761), .B2(n_762), .C(n_763), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g929 ( .A1(n_553), .A2(n_559), .B1(n_930), .B2(n_931), .C(n_932), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g1365 ( .A1(n_553), .A2(n_559), .B1(n_1366), .B2(n_1367), .Y(n_1365) );
AND2x2_ASAP7_75t_L g559 ( .A(n_554), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x6_ASAP7_75t_L g563 ( .A(n_555), .B(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g643 ( .A(n_555), .B(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g645 ( .A(n_555), .B(n_646), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g1362 ( .A1(n_556), .A2(n_562), .B1(n_1363), .B2(n_1364), .Y(n_1362) );
CKINVDCx6p67_ASAP7_75t_R g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g813 ( .A(n_561), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_561), .A2(n_825), .B1(n_897), .B2(n_899), .Y(n_912) );
INVx2_ASAP7_75t_SL g1065 ( .A(n_561), .Y(n_1065) );
CKINVDCx6p67_ASAP7_75t_R g562 ( .A(n_563), .Y(n_562) );
OAI21xp33_ASAP7_75t_L g683 ( .A1(n_564), .A2(n_684), .B(n_685), .Y(n_683) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx4f_ASAP7_75t_L g579 ( .A(n_565), .Y(n_579) );
INVx1_ASAP7_75t_L g695 ( .A(n_565), .Y(n_695) );
INVx1_ASAP7_75t_L g703 ( .A(n_565), .Y(n_703) );
AO22x2_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_647), .B2(n_648), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND4x1_ASAP7_75t_L g569 ( .A(n_570), .B(n_597), .C(n_635), .D(n_639), .Y(n_569) );
NOR3xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_594), .C(n_595), .Y(n_570) );
OAI221xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_576), .B1(n_577), .B2(n_580), .C(n_581), .Y(n_572) );
BUFx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI221xp5_ASAP7_75t_SL g1420 ( .A1(n_574), .A2(n_923), .B1(n_1394), .B2(n_1397), .C(n_1421), .Y(n_1420) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_576), .A2(n_580), .B1(n_622), .B2(n_624), .C(n_626), .Y(n_621) );
BUFx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g589 ( .A(n_579), .Y(n_589) );
INVx2_ASAP7_75t_SL g754 ( .A(n_579), .Y(n_754) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OAI221xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B1(n_589), .B2(n_590), .C(n_591), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_586), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1014) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g644 ( .A(n_587), .Y(n_644) );
INVx2_ASAP7_75t_L g753 ( .A(n_587), .Y(n_753) );
OAI211xp5_ASAP7_75t_L g1026 ( .A1(n_589), .A2(n_1027), .B(n_1028), .C(n_1029), .Y(n_1026) );
BUFx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_SL g947 ( .A(n_593), .Y(n_947) );
OAI31xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_620), .A3(n_633), .B(n_634), .Y(n_597) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_603), .B1(n_604), .B2(n_607), .C(n_608), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g629 ( .A(n_601), .Y(n_629) );
INVx1_ASAP7_75t_L g796 ( .A(n_601), .Y(n_796) );
INVx2_ASAP7_75t_L g871 ( .A(n_601), .Y(n_871) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_602), .A2(n_1045), .B1(n_1086), .B2(n_1087), .Y(n_1085) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_SL g888 ( .A(n_611), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B1(n_617), .B2(n_618), .Y(n_613) );
CKINVDCx11_ASAP7_75t_R g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g791 ( .A(n_623), .Y(n_791) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_SL g627 ( .A1(n_628), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_627) );
AOI31xp33_ASAP7_75t_L g939 ( .A1(n_634), .A2(n_940), .A3(n_954), .B(n_968), .Y(n_939) );
INVx1_ASAP7_75t_L g1032 ( .A(n_634), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_637), .B(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_637), .B(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g1337 ( .A(n_637), .Y(n_1337) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_667), .C(n_677), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_666), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B1(n_658), .B2(n_659), .C(n_660), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_659), .A2(n_688), .B1(n_689), .B2(n_691), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .C(n_665), .Y(n_661) );
AOI33xp33_ASAP7_75t_L g1034 ( .A1(n_665), .A2(n_1035), .A3(n_1036), .B1(n_1039), .B2(n_1043), .B3(n_1046), .Y(n_1034) );
NOR2xp33_ASAP7_75t_SL g667 ( .A(n_668), .B(n_674), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g1388 ( .A(n_670), .Y(n_1388) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_L g1408 ( .A(n_672), .Y(n_1408) );
INVx2_ASAP7_75t_SL g996 ( .A(n_673), .Y(n_996) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI31xp33_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_680), .A3(n_682), .B(n_708), .Y(n_677) );
OAI211xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_687), .B(n_693), .C(n_700), .Y(n_682) );
BUFx3_ASAP7_75t_L g1426 ( .A(n_686), .Y(n_1426) );
OAI221xp5_ASAP7_75t_L g756 ( .A1(n_689), .A2(n_754), .B1(n_757), .B2(n_758), .C(n_759), .Y(n_756) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI211xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B(n_696), .C(n_697), .Y(n_693) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_698), .Y(n_823) );
INVx1_ASAP7_75t_L g959 ( .A(n_698), .Y(n_959) );
NAND2xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_708), .A2(n_807), .B1(n_827), .B2(n_828), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_1006), .B1(n_1103), .B2(n_1104), .Y(n_711) );
INVx1_ASAP7_75t_L g1103 ( .A(n_712), .Y(n_1103) );
XNOR2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_766), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g764 ( .A(n_716), .Y(n_764) );
NAND4xp25_ASAP7_75t_L g716 ( .A(n_717), .B(n_745), .C(n_747), .D(n_760), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_731), .B(n_744), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_726), .B(n_728), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_732) );
BUFx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g1401 ( .A(n_734), .Y(n_1401) );
OAI221xp5_ASAP7_75t_L g752 ( .A1(n_739), .A2(n_742), .B1(n_753), .B2(n_754), .C(n_755), .Y(n_752) );
INVx3_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g1081 ( .A1(n_743), .A2(n_1082), .B(n_1085), .Y(n_1081) );
INVx2_ASAP7_75t_L g1354 ( .A(n_743), .Y(n_1354) );
INVx3_ASAP7_75t_L g1063 ( .A(n_750), .Y(n_1063) );
OAI21xp33_ASAP7_75t_L g1018 ( .A1(n_754), .A2(n_1019), .B(n_1020), .Y(n_1018) );
XNOR2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_875), .Y(n_766) );
AO22x2_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_769), .B1(n_829), .B2(n_830), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
XNOR2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
AND2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_806), .Y(n_771) );
NOR3xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_782), .C(n_786), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_778), .Y(n_773) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g801 ( .A1(n_789), .A2(n_802), .B1(n_803), .B2(n_805), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_797), .B1(n_798), .B2(n_800), .Y(n_795) );
AOI211xp5_ASAP7_75t_SL g808 ( .A1(n_797), .A2(n_809), .B(n_810), .C(n_812), .Y(n_808) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND3xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_815), .C(n_826), .Y(n_807) );
AOI211xp5_ASAP7_75t_SL g834 ( .A1(n_809), .A2(n_835), .B(n_836), .C(n_838), .Y(n_834) );
AOI221xp5_ASAP7_75t_L g940 ( .A1(n_809), .A2(n_941), .B1(n_945), .B2(n_948), .C(n_949), .Y(n_940) );
INVx1_ASAP7_75t_L g1415 ( .A(n_811), .Y(n_1415) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g846 ( .A(n_819), .Y(n_846) );
INVxp67_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx3_ASAP7_75t_L g1423 ( .A(n_821), .Y(n_1423) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
AND2x2_ASAP7_75t_L g831 ( .A(n_832), .B(n_855), .Y(n_831) );
NAND3xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_843), .C(n_851), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_835), .A2(n_853), .B1(n_871), .B2(n_872), .Y(n_870) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx4_ASAP7_75t_L g942 ( .A(n_849), .Y(n_942) );
INVx1_ASAP7_75t_L g1428 ( .A(n_850), .Y(n_1428) );
NOR3xp33_ASAP7_75t_SL g855 ( .A(n_856), .B(n_862), .C(n_863), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_860), .Y(n_856) );
INVx2_ASAP7_75t_SL g1000 ( .A(n_872), .Y(n_1000) );
OAI22xp33_ASAP7_75t_L g1391 ( .A1(n_872), .A2(n_1392), .B1(n_1393), .B2(n_1394), .Y(n_1391) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_933), .B1(n_1004), .B2(n_1005), .Y(n_875) );
INVx1_ASAP7_75t_L g1004 ( .A(n_876), .Y(n_1004) );
NAND4xp25_ASAP7_75t_L g877 ( .A(n_878), .B(n_904), .C(n_906), .D(n_929), .Y(n_877) );
OAI21xp5_ASAP7_75t_SL g878 ( .A1(n_879), .A2(n_893), .B(n_903), .Y(n_878) );
AOI21xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_884), .B(n_889), .Y(n_880) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_891), .A2(n_892), .B1(n_919), .B2(n_921), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_895), .A2(n_897), .B1(n_898), .B2(n_899), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVxp67_ASAP7_75t_SL g1005 ( .A(n_933), .Y(n_1005) );
XNOR2x1_ASAP7_75t_SL g933 ( .A(n_934), .B(n_935), .Y(n_933) );
OAI22xp33_ASAP7_75t_L g1158 ( .A1(n_934), .A2(n_1159), .B1(n_1161), .B2(n_1162), .Y(n_1158) );
AND2x2_ASAP7_75t_L g935 ( .A(n_936), .B(n_971), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g936 ( .A1(n_937), .A2(n_938), .B(n_939), .Y(n_936) );
BUFx2_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx2_ASAP7_75t_SL g952 ( .A(n_953), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g954 ( .A1(n_955), .A2(n_957), .B1(n_963), .B2(n_964), .C(n_965), .Y(n_954) );
INVx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx1_ASAP7_75t_SL g966 ( .A(n_967), .Y(n_966) );
AND4x1_ASAP7_75t_L g971 ( .A(n_972), .B(n_981), .C(n_985), .D(n_988), .Y(n_971) );
AOI221xp5_ASAP7_75t_L g972 ( .A1(n_973), .A2(n_974), .B1(n_975), .B2(n_978), .C(n_979), .Y(n_972) );
AOI221xp5_ASAP7_75t_L g1048 ( .A1(n_973), .A2(n_975), .B1(n_979), .B2(n_1024), .C(n_1025), .Y(n_1048) );
AOI21xp5_ASAP7_75t_L g1439 ( .A1(n_973), .A2(n_979), .B(n_1416), .Y(n_1439) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
AOI33xp33_ASAP7_75t_L g988 ( .A1(n_989), .A2(n_992), .A3(n_997), .B1(n_999), .B2(n_1001), .B3(n_1003), .Y(n_988) );
INVx2_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx2_ASAP7_75t_SL g993 ( .A(n_994), .Y(n_993) );
INVx2_ASAP7_75t_L g1047 ( .A(n_994), .Y(n_1047) );
INVx2_ASAP7_75t_SL g995 ( .A(n_996), .Y(n_995) );
INVx2_ASAP7_75t_L g1407 ( .A(n_1003), .Y(n_1407) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1006), .Y(n_1104) );
AOI22xp5_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1008), .B1(n_1056), .B2(n_1101), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
HB1xp67_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1010), .Y(n_1055) );
NAND4xp75_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .C(n_1033), .D(n_1049), .Y(n_1010) );
OAI31xp33_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1022), .A3(n_1031), .B(n_1032), .Y(n_1012) );
AOI31xp33_ASAP7_75t_L g1338 ( .A1(n_1032), .A2(n_1339), .A3(n_1347), .B(n_1350), .Y(n_1338) );
AND2x2_ASAP7_75t_SL g1033 ( .A(n_1034), .B(n_1048), .Y(n_1033) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1057), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVxp67_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
NOR4xp75_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1077), .C(n_1099), .D(n_1100), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1073), .Y(n_1061) );
AOI33xp33_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1064), .A3(n_1067), .B1(n_1068), .B2(n_1070), .B3(n_1072), .Y(n_1062) );
AOI33xp33_ASAP7_75t_L g1356 ( .A1(n_1063), .A2(n_1072), .A3(n_1357), .B1(n_1358), .B2(n_1360), .B3(n_1361), .Y(n_1356) );
AOI21x1_ASAP7_75t_L g1077 ( .A1(n_1078), .A2(n_1088), .B(n_1098), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1097), .Y(n_1095) );
INVx2_ASAP7_75t_L g1434 ( .A(n_1098), .Y(n_1434) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
OAI221xp5_ASAP7_75t_L g1105 ( .A1(n_1106), .A2(n_1332), .B1(n_1333), .B2(n_1372), .C(n_1376), .Y(n_1105) );
AOI211xp5_ASAP7_75t_SL g1106 ( .A1(n_1107), .A2(n_1216), .B(n_1230), .C(n_1291), .Y(n_1106) );
A2O1A1Ixp33_ASAP7_75t_L g1107 ( .A1(n_1108), .A2(n_1178), .B(n_1185), .C(n_1188), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_1109), .A2(n_1137), .B1(n_1139), .B2(n_1168), .Y(n_1108) );
NOR4xp25_ASAP7_75t_L g1185 ( .A(n_1109), .B(n_1153), .C(n_1168), .D(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1109), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1133), .Y(n_1109) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1110), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1110), .B(n_1192), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1110), .B(n_1134), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1130), .Y(n_1110) );
INVxp67_ASAP7_75t_SL g1181 ( .A(n_1111), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1111), .B(n_1167), .Y(n_1183) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1111), .Y(n_1198) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1111), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1111), .B(n_1134), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1124), .Y(n_1111) );
AND2x4_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1119), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1115), .B(n_1120), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1118), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g1444 ( .A(n_1116), .Y(n_1444) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1118), .Y(n_1128) );
AND2x4_ASAP7_75t_L g1121 ( .A(n_1119), .B(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1163 ( .A(n_1120), .B(n_1123), .Y(n_1163) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1127), .Y(n_1125) );
AND2x4_ASAP7_75t_L g1129 ( .A(n_1126), .B(n_1128), .Y(n_1129) );
AND2x4_ASAP7_75t_L g1145 ( .A(n_1126), .B(n_1127), .Y(n_1145) );
HB1xp67_ASAP7_75t_L g1445 ( .A(n_1127), .Y(n_1445) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1129), .Y(n_1147) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1130), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1130), .B(n_1181), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1132), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1133), .B(n_1156), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1133), .B(n_1197), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1133), .B(n_1252), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1133), .B(n_1183), .Y(n_1270) );
OAI22xp33_ASAP7_75t_L g1273 ( .A1(n_1133), .A2(n_1274), .B1(n_1276), .B2(n_1279), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1133), .B(n_1267), .Y(n_1310) );
CKINVDCx5p33_ASAP7_75t_R g1133 ( .A(n_1134), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1134), .B(n_1165), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1134), .B(n_1180), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1134), .B(n_1155), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1134), .B(n_1197), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1134), .B(n_1203), .Y(n_1255) );
NOR2xp33_ASAP7_75t_L g1278 ( .A(n_1134), .B(n_1166), .Y(n_1278) );
AND2x4_ASAP7_75t_SL g1134 ( .A(n_1135), .B(n_1136), .Y(n_1134) );
INVxp67_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1153), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1149), .Y(n_1139) );
NAND2xp5_ASAP7_75t_SL g1208 ( .A(n_1140), .B(n_1209), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1140), .B(n_1175), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1140), .B(n_1186), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1140), .B(n_1187), .Y(n_1317) );
CKINVDCx6p67_ASAP7_75t_R g1140 ( .A(n_1141), .Y(n_1140) );
CKINVDCx5p33_ASAP7_75t_R g1204 ( .A(n_1141), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1141), .B(n_1149), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1141), .B(n_1207), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1141), .B(n_1209), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1141), .B(n_1150), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1294 ( .A(n_1141), .B(n_1173), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1141), .B(n_1302), .Y(n_1301) );
OR2x2_ASAP7_75t_L g1311 ( .A(n_1141), .B(n_1149), .Y(n_1311) );
OR2x6_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1143), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_1142), .B(n_1143), .Y(n_1232) );
OAI22xp5_ASAP7_75t_SL g1143 ( .A1(n_1144), .A2(n_1146), .B1(n_1147), .B2(n_1148), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
BUFx3_ASAP7_75t_L g1222 ( .A(n_1145), .Y(n_1222) );
INVx2_ASAP7_75t_L g1157 ( .A(n_1147), .Y(n_1157) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1147), .Y(n_1223) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1149), .Y(n_1193) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1150), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1150), .B(n_1187), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1150), .B(n_1175), .Y(n_1201) );
BUFx6f_ASAP7_75t_L g1244 ( .A(n_1150), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1152), .Y(n_1150) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1153), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1164), .Y(n_1153) );
NOR2x1p5_ASAP7_75t_L g1252 ( .A(n_1154), .B(n_1253), .Y(n_1252) );
INVxp67_ASAP7_75t_L g1302 ( .A(n_1154), .Y(n_1302) );
INVx2_ASAP7_75t_SL g1154 ( .A(n_1155), .Y(n_1154) );
BUFx3_ASAP7_75t_L g1171 ( .A(n_1155), .Y(n_1171) );
BUFx2_ASAP7_75t_L g1192 ( .A(n_1155), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1155), .B(n_1213), .Y(n_1258) );
INVx2_ASAP7_75t_SL g1155 ( .A(n_1156), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1156), .B(n_1187), .Y(n_1207) );
BUFx3_ASAP7_75t_L g1226 ( .A(n_1159), .Y(n_1226) );
BUFx6f_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
HB1xp67_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1163), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1164), .B(n_1171), .Y(n_1236) );
INVxp67_ASAP7_75t_L g1303 ( .A(n_1164), .Y(n_1303) );
AOI311xp33_ASAP7_75t_L g1263 ( .A1(n_1165), .A2(n_1204), .A3(n_1264), .B(n_1266), .C(n_1273), .Y(n_1263) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
O2A1O1Ixp33_ASAP7_75t_L g1260 ( .A1(n_1166), .A2(n_1173), .B(n_1261), .C(n_1262), .Y(n_1260) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1167), .B(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1172), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1321 ( .A(n_1170), .B(n_1294), .Y(n_1321) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1171), .B(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1173), .Y(n_1235) );
INVx2_ASAP7_75t_L g1298 ( .A(n_1173), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1175), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1174), .B(n_1187), .Y(n_1209) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1175), .Y(n_1187) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1175), .Y(n_1213) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1175), .Y(n_1237) );
AOI211xp5_ASAP7_75t_SL g1250 ( .A1(n_1175), .A2(n_1251), .B(n_1254), .C(n_1260), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1177), .Y(n_1175) );
NOR2xp33_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1182), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1180), .B(n_1215), .Y(n_1214) );
NAND3xp33_ASAP7_75t_L g1257 ( .A(n_1180), .B(n_1258), .C(n_1259), .Y(n_1257) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1180), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1180), .B(n_1184), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1184), .Y(n_1182) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1183), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1183), .B(n_1215), .Y(n_1282) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1186), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1186), .B(n_1192), .Y(n_1265) );
AOI21xp5_ASAP7_75t_L g1188 ( .A1(n_1189), .A2(n_1204), .B(n_1205), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_1190), .A2(n_1194), .B1(n_1199), .B2(n_1202), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1193), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1192), .B(n_1201), .Y(n_1200) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1192), .B(n_1243), .Y(n_1242) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1192), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1267 ( .A(n_1192), .B(n_1268), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1196), .Y(n_1194) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1201), .Y(n_1315) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1202), .Y(n_1304) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
AOI221xp5_ASAP7_75t_L g1320 ( .A1(n_1204), .A2(n_1321), .B1(n_1322), .B2(n_1323), .C(n_1327), .Y(n_1320) );
A2O1A1Ixp33_ASAP7_75t_L g1205 ( .A1(n_1206), .A2(n_1208), .B(n_1210), .C(n_1212), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1209), .Y(n_1307) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_1210), .A2(n_1261), .B1(n_1287), .B2(n_1288), .Y(n_1286) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1214), .Y(n_1212) );
NAND2xp67_ASAP7_75t_L g1324 ( .A(n_1213), .B(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1214), .Y(n_1329) );
AOI32xp33_ASAP7_75t_L g1230 ( .A1(n_1216), .A2(n_1231), .A3(n_1250), .B1(n_1263), .B2(n_1281), .Y(n_1230) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
OAI211xp5_ASAP7_75t_L g1254 ( .A1(n_1217), .A2(n_1255), .B(n_1256), .C(n_1257), .Y(n_1254) );
INVx3_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
AOI211xp5_ASAP7_75t_L g1314 ( .A1(n_1219), .A2(n_1315), .B(n_1316), .C(n_1318), .Y(n_1314) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
CKINVDCx5p33_ASAP7_75t_R g1332 ( .A(n_1222), .Y(n_1332) );
OAI22xp33_ASAP7_75t_L g1224 ( .A1(n_1225), .A2(n_1226), .B1(n_1227), .B2(n_1228), .Y(n_1224) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
AOI211xp5_ASAP7_75t_L g1231 ( .A1(n_1232), .A2(n_1233), .B(n_1238), .C(n_1241), .Y(n_1231) );
OAI22xp5_ASAP7_75t_L g1233 ( .A1(n_1234), .A2(n_1235), .B1(n_1236), .B2(n_1237), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1237), .B(n_1239), .Y(n_1238) );
INVx3_ASAP7_75t_L g1285 ( .A(n_1237), .Y(n_1285) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1240), .Y(n_1262) );
OAI222xp33_ASAP7_75t_L g1241 ( .A1(n_1242), .A2(n_1243), .B1(n_1244), .B2(n_1245), .C1(n_1246), .C2(n_1248), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g1296 ( .A1(n_1242), .A2(n_1248), .B1(n_1297), .B2(n_1299), .Y(n_1296) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1243), .Y(n_1331) );
CKINVDCx14_ASAP7_75t_R g1259 ( .A(n_1244), .Y(n_1259) );
A2O1A1Ixp33_ASAP7_75t_L g1327 ( .A1(n_1245), .A2(n_1328), .B(n_1329), .C(n_1330), .Y(n_1327) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1251), .Y(n_1326) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1255), .Y(n_1322) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1261), .Y(n_1287) );
AOI221xp5_ASAP7_75t_L g1309 ( .A1(n_1261), .A2(n_1267), .B1(n_1276), .B2(n_1310), .C(n_1311), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1261), .B(n_1289), .Y(n_1319) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
AOI21xp33_ASAP7_75t_SL g1266 ( .A1(n_1267), .A2(n_1269), .B(n_1271), .Y(n_1266) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1267), .Y(n_1295) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1270), .B(n_1275), .Y(n_1313) );
CKINVDCx5p33_ASAP7_75t_R g1271 ( .A(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
HB1xp67_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_1280), .B(n_1331), .Y(n_1330) );
A2O1A1Ixp33_ASAP7_75t_SL g1281 ( .A1(n_1282), .A2(n_1283), .B(n_1286), .C(n_1290), .Y(n_1281) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
AOI21xp33_ASAP7_75t_L g1305 ( .A1(n_1288), .A2(n_1306), .B(n_1307), .Y(n_1305) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
NAND3xp33_ASAP7_75t_SL g1291 ( .A(n_1292), .B(n_1308), .C(n_1320), .Y(n_1291) );
AOI211xp5_ASAP7_75t_L g1292 ( .A1(n_1293), .A2(n_1295), .B(n_1296), .C(n_1305), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
NAND3xp33_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1303), .C(n_1304), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
NOR3xp33_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1312), .C(n_1314), .Y(n_1308) );
INVxp67_ASAP7_75t_SL g1312 ( .A(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
NAND2xp5_ASAP7_75t_SL g1323 ( .A(n_1324), .B(n_1326), .Y(n_1323) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1325), .Y(n_1328) );
HB1xp67_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
XOR2x2_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1371), .Y(n_1334) );
NOR3xp33_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1338), .C(n_1355), .Y(n_1335) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
NAND4xp25_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1362), .C(n_1365), .D(n_1368), .Y(n_1355) );
INVx2_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
CKINVDCx5p33_ASAP7_75t_R g1378 ( .A(n_1379), .Y(n_1378) );
A2O1A1Ixp33_ASAP7_75t_L g1442 ( .A1(n_1380), .A2(n_1443), .B(n_1445), .C(n_1446), .Y(n_1442) );
INVxp33_ASAP7_75t_SL g1381 ( .A(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1384), .Y(n_1440) );
HB1xp67_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1386), .B(n_1409), .Y(n_1385) );
NOR2xp33_ASAP7_75t_L g1386 ( .A(n_1387), .B(n_1390), .Y(n_1386) );
OAI22xp5_ASAP7_75t_L g1398 ( .A1(n_1399), .A2(n_1400), .B1(n_1402), .B2(n_1403), .Y(n_1398) );
INVx2_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
AOI21xp5_ASAP7_75t_SL g1409 ( .A1(n_1410), .A2(n_1433), .B(n_1435), .Y(n_1409) );
NAND4xp25_ASAP7_75t_SL g1410 ( .A(n_1411), .B(n_1418), .C(n_1420), .D(n_1424), .Y(n_1410) );
INVx2_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
OAI221xp5_ASAP7_75t_L g1424 ( .A1(n_1425), .A2(n_1427), .B1(n_1428), .B2(n_1429), .C(n_1430), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
HB1xp67_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
endmodule