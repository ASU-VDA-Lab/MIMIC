module fake_netlist_5_1737_n_756 (n_137, n_91, n_82, n_122, n_10, n_140, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_756);

input n_137;
input n_91;
input n_82;
input n_122;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_756;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_688;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_658;
wire n_281;
wire n_647;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_208;
wire n_142;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_144;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_656;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_401;
wire n_187;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_26),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_51),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_40),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_36),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_66),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_13),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

NOR2xp67_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_37),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_47),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_21),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_44),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_38),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_95),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_41),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_50),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_59),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_56),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_34),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_31),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_11),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_22),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_114),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_92),
.B(n_35),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_5),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_46),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_91),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_77),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_137),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_61),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_102),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_75),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_97),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_64),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_65),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_18),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_90),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_57),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_71),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_43),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_88),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_17),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_49),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_23),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_39),
.Y(n_196)
);

BUFx8_ASAP7_75t_SL g197 ( 
.A(n_166),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

BUFx8_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_152),
.B(n_0),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_143),
.B(n_0),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_141),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_158),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_161),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_164),
.B(n_1),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_2),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_179),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_181),
.B(n_3),
.Y(n_227)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_142),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

BUFx8_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

OAI22x1_ASAP7_75t_L g234 ( 
.A1(n_196),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_148),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_150),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_151),
.B(n_4),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_153),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_197),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_213),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_R g242 ( 
.A(n_230),
.B(n_184),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_237),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_149),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_228),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_201),
.B(n_166),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_228),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_210),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_228),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_236),
.Y(n_253)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_R g255 ( 
.A(n_201),
.B(n_154),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_208),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_236),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_R g259 ( 
.A(n_221),
.B(n_6),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_200),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_236),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_236),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_214),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_239),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_200),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_202),
.B(n_155),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_239),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_239),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_203),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_203),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_216),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_215),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_209),
.A2(n_190),
.B1(n_191),
.B2(n_194),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_212),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_R g280 ( 
.A(n_212),
.B(n_159),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_233),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_233),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_208),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_199),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_199),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_223),
.Y(n_286)
);

NOR3xp33_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_217),
.C(n_209),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_286),
.B(n_225),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_266),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_225),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_202),
.Y(n_294)
);

NOR3xp33_ASAP7_75t_L g295 ( 
.A(n_247),
.B(n_238),
.C(n_205),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_254),
.B(n_244),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_255),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_254),
.B(n_226),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_223),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_244),
.B(n_226),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_255),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_266),
.A2(n_221),
.B1(n_227),
.B2(n_222),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_260),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_206),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_L g306 ( 
.A(n_253),
.B(n_222),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

NAND2x1_ASAP7_75t_L g308 ( 
.A(n_245),
.B(n_204),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_L g309 ( 
.A(n_258),
.B(n_224),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_267),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_250),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_259),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_261),
.B(n_231),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_262),
.B(n_238),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_279),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_265),
.B(n_206),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_251),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

NOR3xp33_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_205),
.C(n_229),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_270),
.Y(n_323)
);

NOR3xp33_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_229),
.C(n_224),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_242),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_271),
.B(n_227),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_246),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_219),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_242),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_280),
.B(n_167),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_241),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_249),
.B(n_219),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_240),
.Y(n_335)
);

BUFx6f_ASAP7_75t_SL g336 ( 
.A(n_284),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_252),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_243),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_281),
.B(n_215),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_285),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_282),
.B(n_218),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_286),
.B(n_172),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_269),
.B(n_231),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_242),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_275),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_275),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_286),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_L g348 ( 
.A(n_241),
.B(n_173),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_275),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_266),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_293),
.B(n_294),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_174),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_299),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_322),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_310),
.B(n_198),
.Y(n_357)
);

AND2x4_ASAP7_75t_SL g358 ( 
.A(n_323),
.B(n_218),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_313),
.B(n_218),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_323),
.B(n_175),
.Y(n_360)
);

AND2x6_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_204),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_329),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_312),
.A2(n_182),
.B1(n_186),
.B2(n_189),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_307),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_290),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_312),
.A2(n_195),
.B1(n_232),
.B2(n_220),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_313),
.B(n_218),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_291),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_297),
.B(n_234),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_300),
.B(n_220),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_287),
.A2(n_295),
.B1(n_306),
.B2(n_309),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_300),
.B(n_220),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_328),
.B(n_220),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_298),
.A2(n_207),
.B(n_204),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_291),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_350),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_291),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_311),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_288),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_316),
.B(n_232),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_329),
.Y(n_384)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_317),
.Y(n_385)
);

NAND2x1p5_ASAP7_75t_L g386 ( 
.A(n_333),
.B(n_207),
.Y(n_386)
);

BUFx8_ASAP7_75t_SL g387 ( 
.A(n_336),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_302),
.A2(n_232),
.B1(n_207),
.B2(n_78),
.Y(n_388)
);

BUFx8_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_296),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_292),
.B(n_7),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_305),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_304),
.A2(n_76),
.B(n_138),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_337),
.Y(n_394)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_317),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_317),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_302),
.B(n_19),
.Y(n_397)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_325),
.B(n_7),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_301),
.B(n_8),
.Y(n_399)
);

A2O1A1Ixp33_ASAP7_75t_L g400 ( 
.A1(n_287),
.A2(n_321),
.B(n_326),
.C(n_349),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_311),
.Y(n_401)
);

O2A1O1Ixp33_ASAP7_75t_L g402 ( 
.A1(n_314),
.A2(n_289),
.B(n_321),
.C(n_334),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_331),
.B(n_344),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_303),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_315),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_345),
.B(n_20),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_346),
.B(n_24),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_330),
.A2(n_80),
.B1(n_136),
.B2(n_135),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_319),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_320),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_308),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_347),
.B(n_8),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_340),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_339),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_324),
.B(n_9),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_351),
.B(n_342),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_380),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_383),
.A2(n_332),
.B(n_341),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_372),
.A2(n_353),
.B1(n_400),
.B2(n_397),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_327),
.Y(n_421)
);

BUFx8_ASAP7_75t_L g422 ( 
.A(n_362),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_355),
.B(n_335),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_352),
.B(n_324),
.Y(n_425)
);

BUFx8_ASAP7_75t_L g426 ( 
.A(n_362),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_401),
.A2(n_348),
.B(n_338),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_L g428 ( 
.A1(n_402),
.A2(n_415),
.B(n_363),
.C(n_357),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_392),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_352),
.B(n_327),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_376),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_406),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_355),
.B(n_10),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_355),
.B(n_12),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_374),
.A2(n_81),
.B(n_133),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_357),
.B(n_12),
.Y(n_436)
);

CKINVDCx10_ASAP7_75t_R g437 ( 
.A(n_387),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_354),
.A2(n_82),
.B1(n_132),
.B2(n_131),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_390),
.A2(n_74),
.B1(n_129),
.B2(n_128),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_371),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_384),
.B(n_25),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_390),
.A2(n_79),
.B1(n_127),
.B2(n_126),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_359),
.B(n_14),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_379),
.B(n_27),
.Y(n_444)
);

OAI21xp33_ASAP7_75t_L g445 ( 
.A1(n_391),
.A2(n_416),
.B(n_370),
.Y(n_445)
);

AOI21x1_ASAP7_75t_L g446 ( 
.A1(n_373),
.A2(n_72),
.B(n_125),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_368),
.B(n_15),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_410),
.Y(n_448)
);

CKINVDCx8_ASAP7_75t_R g449 ( 
.A(n_384),
.Y(n_449)
);

OR2x6_ASAP7_75t_L g450 ( 
.A(n_394),
.B(n_16),
.Y(n_450)
);

NOR3xp33_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_16),
.C(n_17),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_358),
.B(n_28),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_356),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_388),
.A2(n_33),
.B1(n_42),
.B2(n_45),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_411),
.B(n_48),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_396),
.Y(n_456)
);

OAI22x1_ASAP7_75t_L g457 ( 
.A1(n_399),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_457)
);

NOR2xp67_ASAP7_75t_SL g458 ( 
.A(n_385),
.B(n_55),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_403),
.B(n_60),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_395),
.A2(n_67),
.B(n_68),
.Y(n_460)
);

NOR3xp33_ASAP7_75t_L g461 ( 
.A(n_360),
.B(n_69),
.C(n_70),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_366),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_364),
.B(n_83),
.C(n_84),
.Y(n_463)
);

O2A1O1Ixp33_ASAP7_75t_L g464 ( 
.A1(n_367),
.A2(n_85),
.B(n_87),
.C(n_89),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_398),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_395),
.A2(n_93),
.B(n_94),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_396),
.B(n_403),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_365),
.B(n_96),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_423),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_446),
.Y(n_471)
);

CKINVDCx11_ASAP7_75t_R g472 ( 
.A(n_449),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_430),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_427),
.A2(n_408),
.B(n_407),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_417),
.B(n_381),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_432),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_418),
.Y(n_477)
);

BUFx12f_ASAP7_75t_L g478 ( 
.A(n_422),
.Y(n_478)
);

AOI22x1_ASAP7_75t_L g479 ( 
.A1(n_419),
.A2(n_386),
.B1(n_377),
.B2(n_393),
.Y(n_479)
);

NAND2x1p5_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_376),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_456),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_468),
.A2(n_375),
.B(n_378),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_448),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_425),
.B(n_405),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_431),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_456),
.Y(n_486)
);

NAND2x1p5_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_444),
.Y(n_487)
);

OA21x2_ASAP7_75t_L g488 ( 
.A1(n_428),
.A2(n_409),
.B(n_412),
.Y(n_488)
);

BUFx2_ASAP7_75t_SL g489 ( 
.A(n_456),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_444),
.B(n_376),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_455),
.A2(n_369),
.B(n_361),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_437),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_431),
.Y(n_493)
);

AO21x2_ASAP7_75t_L g494 ( 
.A1(n_420),
.A2(n_361),
.B(n_99),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_443),
.A2(n_361),
.B(n_100),
.Y(n_495)
);

AO21x2_ASAP7_75t_L g496 ( 
.A1(n_447),
.A2(n_98),
.B(n_103),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_421),
.B(n_105),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_465),
.B(n_106),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_462),
.Y(n_499)
);

AO21x2_ASAP7_75t_L g500 ( 
.A1(n_461),
.A2(n_107),
.B(n_108),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_436),
.B(n_414),
.Y(n_501)
);

NAND2x1p5_ASAP7_75t_L g502 ( 
.A(n_458),
.B(n_109),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_435),
.A2(n_111),
.B(n_113),
.Y(n_503)
);

OR3x4_ASAP7_75t_SL g504 ( 
.A(n_424),
.B(n_389),
.C(n_116),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_452),
.Y(n_505)
);

BUFx2_ASAP7_75t_R g506 ( 
.A(n_441),
.Y(n_506)
);

AO21x2_ASAP7_75t_L g507 ( 
.A1(n_463),
.A2(n_115),
.B(n_117),
.Y(n_507)
);

INVx6_ASAP7_75t_L g508 ( 
.A(n_422),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_445),
.B(n_119),
.Y(n_509)
);

BUFx8_ASAP7_75t_L g510 ( 
.A(n_426),
.Y(n_510)
);

NAND2x1p5_ASAP7_75t_L g511 ( 
.A(n_438),
.B(n_120),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_467),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_426),
.Y(n_513)
);

BUFx2_ASAP7_75t_R g514 ( 
.A(n_457),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_453),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_464),
.A2(n_122),
.B(n_123),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_509),
.A2(n_451),
.B1(n_434),
.B2(n_433),
.Y(n_517)
);

OAI22xp33_ASAP7_75t_L g518 ( 
.A1(n_501),
.A2(n_450),
.B1(n_439),
.B2(n_442),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_505),
.B(n_450),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_473),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_483),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_475),
.B(n_440),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_484),
.B(n_454),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_499),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_499),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_501),
.A2(n_389),
.B1(n_460),
.B2(n_466),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_508),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_469),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_470),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_486),
.Y(n_531)
);

NAND2x1p5_ASAP7_75t_L g532 ( 
.A(n_488),
.B(n_124),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_509),
.A2(n_139),
.B1(n_497),
.B2(n_484),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_487),
.A2(n_480),
.B1(n_490),
.B2(n_505),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_492),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_515),
.A2(n_477),
.B(n_511),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_487),
.B(n_498),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_476),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_486),
.Y(n_539)
);

OAI21x1_ASAP7_75t_SL g540 ( 
.A1(n_488),
.A2(n_515),
.B(n_479),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_477),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_498),
.B(n_505),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_511),
.A2(n_512),
.B1(n_480),
.B2(n_500),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_485),
.Y(n_544)
);

INVxp33_ASAP7_75t_L g545 ( 
.A(n_472),
.Y(n_545)
);

CKINVDCx11_ASAP7_75t_R g546 ( 
.A(n_478),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_485),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_SL g548 ( 
.A1(n_508),
.A2(n_511),
.B1(n_513),
.B2(n_510),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_480),
.B(n_512),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_490),
.B(n_485),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_493),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_493),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_491),
.A2(n_482),
.B(n_474),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_512),
.A2(n_500),
.B1(n_488),
.B2(n_494),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_489),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_486),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_493),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_R g558 ( 
.A(n_524),
.B(n_471),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_542),
.B(n_512),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_R g560 ( 
.A(n_535),
.B(n_472),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_520),
.B(n_512),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_542),
.B(n_481),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_529),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_519),
.B(n_481),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_549),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_535),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_529),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_528),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_530),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_537),
.B(n_490),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_530),
.Y(n_571)
);

AND2x2_ASAP7_75t_SL g572 ( 
.A(n_554),
.B(n_517),
.Y(n_572)
);

CKINVDCx16_ASAP7_75t_R g573 ( 
.A(n_528),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_538),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_521),
.B(n_486),
.Y(n_575)
);

CKINVDCx9p33_ASAP7_75t_R g576 ( 
.A(n_523),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_522),
.B(n_486),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_528),
.Y(n_578)
);

OA21x2_ASAP7_75t_L g579 ( 
.A1(n_553),
.A2(n_516),
.B(n_495),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_531),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_R g581 ( 
.A(n_546),
.B(n_492),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_519),
.B(n_514),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_R g583 ( 
.A(n_524),
.B(n_508),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_SL g584 ( 
.A(n_548),
.B(n_502),
.C(n_504),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_531),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_538),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_R g587 ( 
.A(n_544),
.B(n_508),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_525),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_519),
.B(n_550),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_526),
.Y(n_590)
);

AO21x2_ASAP7_75t_L g591 ( 
.A1(n_540),
.A2(n_494),
.B(n_495),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_518),
.B(n_506),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_533),
.A2(n_513),
.B1(n_493),
.B2(n_478),
.Y(n_593)
);

BUFx4f_ASAP7_75t_SL g594 ( 
.A(n_531),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_525),
.B(n_493),
.Y(n_595)
);

OR2x6_ASAP7_75t_SL g596 ( 
.A(n_534),
.B(n_510),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_526),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_541),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_550),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_541),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_539),
.B(n_556),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_536),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_547),
.Y(n_603)
);

NOR3xp33_ASAP7_75t_SL g604 ( 
.A(n_551),
.B(n_510),
.C(n_500),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_547),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_555),
.B(n_507),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_606),
.B(n_532),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_565),
.B(n_543),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_561),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_598),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_559),
.B(n_532),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_562),
.B(n_544),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_578),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_589),
.B(n_574),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_598),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_589),
.B(n_532),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_586),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_605),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_603),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_564),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_590),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_592),
.B(n_544),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_563),
.B(n_496),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_597),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_592),
.B(n_527),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_567),
.B(n_556),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_600),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_572),
.A2(n_584),
.B1(n_593),
.B2(n_558),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_578),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_580),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_602),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_602),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_599),
.B(n_496),
.Y(n_633)
);

OAI221xp5_ASAP7_75t_L g634 ( 
.A1(n_604),
.A2(n_502),
.B1(n_545),
.B2(n_551),
.C(n_552),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_571),
.B(n_496),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_601),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_576),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_572),
.A2(n_502),
.B1(n_552),
.B2(n_557),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_570),
.B(n_494),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_625),
.A2(n_582),
.B(n_576),
.Y(n_640)
);

OAI211xp5_ASAP7_75t_L g641 ( 
.A1(n_628),
.A2(n_583),
.B(n_604),
.C(n_587),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_617),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_631),
.B(n_591),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_631),
.B(n_632),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_632),
.B(n_591),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_639),
.B(n_579),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_617),
.B(n_569),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_609),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_621),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_621),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_624),
.B(n_579),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_636),
.B(n_588),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_624),
.B(n_579),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_629),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_627),
.B(n_583),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_627),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_618),
.B(n_575),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_618),
.B(n_577),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_614),
.B(n_573),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_628),
.B(n_634),
.C(n_608),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_610),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_610),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_629),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_639),
.B(n_595),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_607),
.B(n_471),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_614),
.B(n_596),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_615),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_615),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_648),
.B(n_611),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_642),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_664),
.B(n_607),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_644),
.B(n_613),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_649),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_650),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_646),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_664),
.B(n_633),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_656),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_644),
.B(n_613),
.Y(n_678)
);

CKINVDCx16_ASAP7_75t_R g679 ( 
.A(n_666),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_661),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_662),
.Y(n_681)
);

INVxp33_ASAP7_75t_L g682 ( 
.A(n_659),
.Y(n_682)
);

OAI222xp33_ASAP7_75t_L g683 ( 
.A1(n_679),
.A2(n_637),
.B1(n_633),
.B2(n_655),
.C1(n_666),
.C2(n_638),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_676),
.B(n_646),
.Y(n_684)
);

OAI22xp33_ASAP7_75t_L g685 ( 
.A1(n_682),
.A2(n_640),
.B1(n_660),
.B2(n_637),
.Y(n_685)
);

NAND4xp75_ASAP7_75t_L g686 ( 
.A(n_673),
.B(n_655),
.C(n_654),
.D(n_643),
.Y(n_686)
);

OAI32xp33_ASAP7_75t_L g687 ( 
.A1(n_682),
.A2(n_652),
.A3(n_558),
.B1(n_663),
.B2(n_665),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_669),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_678),
.Y(n_689)
);

OAI22xp33_ASAP7_75t_SL g690 ( 
.A1(n_671),
.A2(n_654),
.B1(n_663),
.B2(n_620),
.Y(n_690)
);

OAI32xp33_ASAP7_75t_L g691 ( 
.A1(n_674),
.A2(n_677),
.A3(n_670),
.B1(n_681),
.B2(n_680),
.Y(n_691)
);

OAI21xp33_ASAP7_75t_L g692 ( 
.A1(n_687),
.A2(n_675),
.B(n_641),
.Y(n_692)
);

NAND3xp33_ASAP7_75t_L g693 ( 
.A(n_685),
.B(n_645),
.C(n_643),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_691),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_689),
.B(n_678),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_684),
.B(n_675),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_694),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_693),
.Y(n_698)
);

OAI21xp33_ASAP7_75t_L g699 ( 
.A1(n_692),
.A2(n_690),
.B(n_622),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_695),
.B(n_688),
.Y(n_700)
);

NOR2x1_ASAP7_75t_L g701 ( 
.A(n_696),
.B(n_686),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_695),
.Y(n_702)
);

NAND2x1p5_ASAP7_75t_L g703 ( 
.A(n_701),
.B(n_663),
.Y(n_703)
);

AOI211xp5_ASAP7_75t_L g704 ( 
.A1(n_698),
.A2(n_683),
.B(n_638),
.C(n_560),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_697),
.B(n_689),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_703),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_705),
.B(n_699),
.Y(n_707)
);

AOI221xp5_ASAP7_75t_L g708 ( 
.A1(n_707),
.A2(n_704),
.B1(n_702),
.B2(n_700),
.C(n_581),
.Y(n_708)
);

AOI321xp33_ASAP7_75t_L g709 ( 
.A1(n_706),
.A2(n_612),
.A3(n_645),
.B1(n_678),
.B2(n_672),
.C(n_611),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_706),
.B(n_566),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_710),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_709),
.Y(n_712)
);

INVxp33_ASAP7_75t_SL g713 ( 
.A(n_708),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_710),
.B(n_672),
.Y(n_714)
);

NOR2x1_ASAP7_75t_L g715 ( 
.A(n_710),
.B(n_581),
.Y(n_715)
);

AO22x2_ASAP7_75t_L g716 ( 
.A1(n_708),
.A2(n_670),
.B1(n_630),
.B2(n_560),
.Y(n_716)
);

OAI211xp5_ASAP7_75t_L g717 ( 
.A1(n_715),
.A2(n_587),
.B(n_630),
.C(n_626),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_711),
.B(n_658),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_714),
.Y(n_719)
);

XOR2xp5_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_568),
.Y(n_720)
);

AOI21xp33_ASAP7_75t_L g721 ( 
.A1(n_713),
.A2(n_665),
.B(n_647),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_712),
.B(n_658),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_712),
.B(n_657),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_719),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_723),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_722),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_720),
.Y(n_727)
);

BUFx12f_ASAP7_75t_L g728 ( 
.A(n_717),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_718),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_725),
.Y(n_730)
);

XNOR2xp5_ASAP7_75t_L g731 ( 
.A(n_724),
.B(n_721),
.Y(n_731)
);

XOR2xp5_ASAP7_75t_L g732 ( 
.A(n_727),
.B(n_531),
.Y(n_732)
);

NAND4xp75_ASAP7_75t_L g733 ( 
.A(n_726),
.B(n_647),
.C(n_557),
.D(n_657),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_729),
.Y(n_734)
);

XNOR2xp5_ASAP7_75t_L g735 ( 
.A(n_728),
.B(n_616),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_728),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_725),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_736),
.A2(n_734),
.B1(n_737),
.B2(n_730),
.Y(n_738)
);

AO22x2_ASAP7_75t_L g739 ( 
.A1(n_732),
.A2(n_733),
.B1(n_731),
.B2(n_735),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_730),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_736),
.A2(n_594),
.B1(n_585),
.B2(n_580),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_730),
.B(n_653),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_736),
.A2(n_594),
.B1(n_585),
.B2(n_635),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_736),
.A2(n_667),
.B1(n_668),
.B2(n_619),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_736),
.A2(n_623),
.B1(n_635),
.B2(n_619),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_740),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_738),
.B(n_616),
.Y(n_747)
);

AO22x2_ASAP7_75t_L g748 ( 
.A1(n_742),
.A2(n_668),
.B1(n_623),
.B2(n_651),
.Y(n_748)
);

XOR2x1_ASAP7_75t_L g749 ( 
.A(n_739),
.B(n_531),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_741),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_747),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_746),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_752),
.B(n_749),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_SL g754 ( 
.A1(n_753),
.A2(n_750),
.B1(n_751),
.B2(n_744),
.Y(n_754)
);

AOI221xp5_ASAP7_75t_L g755 ( 
.A1(n_754),
.A2(n_748),
.B1(n_743),
.B2(n_745),
.C(n_507),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_755),
.A2(n_507),
.B1(n_471),
.B2(n_503),
.Y(n_756)
);


endmodule