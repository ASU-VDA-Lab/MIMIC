module real_aes_11473_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_916, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_916;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_635;
wire n_287;
wire n_357;
wire n_386;
wire n_905;
wire n_792;
wire n_518;
wire n_254;
wire n_673;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_733;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
wire n_862;
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_0), .A2(n_87), .B1(n_522), .B2(n_523), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_1), .B(n_190), .Y(n_574) );
AOI22x1_ASAP7_75t_SL g109 ( .A1(n_2), .A2(n_76), .B1(n_110), .B2(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_3), .B(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_4), .B(n_131), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_5), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_6), .A2(n_40), .B1(n_162), .B2(n_520), .Y(n_635) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_7), .B(n_89), .Y(n_505) );
INVx1_ASAP7_75t_L g910 ( .A(n_7), .Y(n_910) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_8), .B(n_142), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_9), .B(n_123), .Y(n_150) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_10), .A2(n_65), .B1(n_162), .B2(n_201), .Y(n_533) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_11), .B(n_145), .C(n_162), .Y(n_595) );
NAND2x1p5_ASAP7_75t_L g226 ( .A(n_12), .B(n_123), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_13), .B(n_181), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_14), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_15), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_16), .B(n_135), .Y(n_559) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_17), .A2(n_883), .B1(n_885), .B2(n_886), .Y(n_882) );
INVxp33_ASAP7_75t_L g885 ( .A(n_17), .Y(n_885) );
AND2x2_ASAP7_75t_L g200 ( .A(n_18), .B(n_201), .Y(n_200) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_19), .B(n_138), .C(n_142), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_20), .A2(n_28), .B1(n_142), .B2(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_21), .B(n_561), .Y(n_609) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_22), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_23), .B(n_263), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_24), .B(n_189), .Y(n_188) );
NAND2xp33_ASAP7_75t_L g219 ( .A(n_25), .B(n_130), .Y(n_219) );
NAND2xp33_ASAP7_75t_L g143 ( .A(n_26), .B(n_130), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g912 ( .A(n_27), .Y(n_912) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_29), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_30), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_31), .B(n_551), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_32), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_33), .A2(n_84), .B1(n_876), .B2(n_877), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_33), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_34), .A2(n_55), .B1(n_130), .B2(n_201), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_35), .B(n_138), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_36), .B(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g504 ( .A(n_37), .Y(n_504) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_38), .A2(n_68), .B(n_126), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_39), .A2(n_164), .B(n_206), .C(n_207), .Y(n_205) );
NAND2xp33_ASAP7_75t_L g260 ( .A(n_41), .B(n_168), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_42), .B(n_162), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_43), .Y(n_279) );
AND2x6_ASAP7_75t_L g148 ( .A(n_44), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g535 ( .A(n_45), .B(n_263), .Y(n_535) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_45), .Y(n_884) );
NAND2x1p5_ASAP7_75t_L g596 ( .A(n_46), .B(n_263), .Y(n_596) );
OAI22x1_ASAP7_75t_SL g857 ( .A1(n_47), .A2(n_49), .B1(n_858), .B2(n_859), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_47), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_48), .B(n_161), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g858 ( .A(n_49), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_50), .B(n_141), .Y(n_140) );
NAND2xp33_ASAP7_75t_L g186 ( .A(n_51), .B(n_168), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_52), .B(n_135), .Y(n_611) );
INVx1_ASAP7_75t_L g149 ( .A(n_53), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_54), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_56), .B(n_168), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_57), .B(n_263), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_58), .B(n_142), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_59), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_60), .B(n_142), .Y(n_549) );
NAND2x1_ASAP7_75t_L g615 ( .A(n_61), .B(n_263), .Y(n_615) );
AND2x2_ASAP7_75t_L g209 ( .A(n_62), .B(n_189), .Y(n_209) );
AND2x2_ASAP7_75t_L g906 ( .A(n_63), .B(n_907), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_64), .B(n_145), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_66), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_67), .B(n_543), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_69), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_70), .Y(n_546) );
NAND2xp33_ASAP7_75t_L g242 ( .A(n_71), .B(n_135), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g894 ( .A(n_72), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_73), .B(n_145), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_74), .A2(n_79), .B1(n_142), .B2(n_520), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_75), .B(n_218), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_76), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_77), .Y(n_582) );
BUFx10_ASAP7_75t_L g861 ( .A(n_78), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_80), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_SL g526 ( .A(n_81), .Y(n_526) );
NAND2xp33_ASAP7_75t_L g247 ( .A(n_82), .B(n_142), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_83), .Y(n_638) );
INVx1_ASAP7_75t_L g877 ( .A(n_84), .Y(n_877) );
NAND2xp5_ASAP7_75t_SL g129 ( .A(n_85), .B(n_130), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_86), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_88), .Y(n_208) );
AND2x2_ASAP7_75t_L g909 ( .A(n_89), .B(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g126 ( .A(n_90), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_91), .B(n_145), .Y(n_594) );
BUFx2_ASAP7_75t_L g501 ( .A(n_92), .Y(n_501) );
OR2x2_ASAP7_75t_L g870 ( .A(n_92), .B(n_502), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_92), .B(n_503), .Y(n_899) );
INVx1_ASAP7_75t_L g908 ( .A(n_92), .Y(n_908) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_93), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_94), .B(n_168), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_95), .B(n_225), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_96), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_97), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g907 ( .A(n_98), .Y(n_907) );
INVx1_ASAP7_75t_L g199 ( .A(n_99), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_100), .Y(n_160) );
AND2x2_ASAP7_75t_L g173 ( .A(n_101), .B(n_123), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_102), .B(n_171), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_103), .B(n_189), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_900), .B(n_911), .Y(n_104) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_862), .B(n_865), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_856), .B(n_860), .Y(n_106) );
AOI22xp33_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_499), .B1(n_506), .B2(n_507), .Y(n_107) );
INVx1_ASAP7_75t_L g864 ( .A(n_108), .Y(n_864) );
XNOR2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
XNOR2x1_ASAP7_75t_L g508 ( .A(n_109), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g880 ( .A(n_112), .B(n_875), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_112), .A2(n_874), .B1(n_875), .B2(n_879), .Y(n_887) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g879 ( .A(n_113), .Y(n_879) );
NAND2x1p5_ASAP7_75t_L g113 ( .A(n_114), .B(n_416), .Y(n_113) );
AND5x1_ASAP7_75t_L g114 ( .A(n_115), .B(n_319), .C(n_358), .D(n_384), .E(n_399), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_286), .Y(n_115) );
OAI221xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_210), .B1(n_227), .B2(n_237), .C(n_265), .Y(n_116) );
OR2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_151), .Y(n_117) );
INVx1_ASAP7_75t_L g383 ( .A(n_118), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_118), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_118), .B(n_268), .Y(n_467) );
AOI322xp5_ASAP7_75t_L g480 ( .A1(n_118), .A2(n_349), .A3(n_402), .B1(n_481), .B2(n_483), .C1(n_484), .C2(n_487), .Y(n_480) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g368 ( .A(n_119), .B(n_235), .Y(n_368) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_120), .Y(n_236) );
INVx1_ASAP7_75t_L g303 ( .A(n_120), .Y(n_303) );
AND2x2_ASAP7_75t_L g308 ( .A(n_120), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g318 ( .A(n_120), .B(n_232), .Y(n_318) );
AND2x2_ASAP7_75t_L g326 ( .A(n_120), .B(n_174), .Y(n_326) );
INVx1_ASAP7_75t_L g340 ( .A(n_120), .Y(n_340) );
OAI21x1_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_127), .B(n_150), .Y(n_120) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_121), .A2(n_254), .B(n_262), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g282 ( .A1(n_121), .A2(n_254), .B(n_262), .Y(n_282) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_121), .A2(n_588), .B(n_596), .Y(n_587) );
OAI21x1_ASAP7_75t_L g646 ( .A1(n_121), .A2(n_588), .B(n_596), .Y(n_646) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g633 ( .A(n_122), .B(n_146), .Y(n_633) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx4_ASAP7_75t_L g154 ( .A(n_123), .Y(n_154) );
BUFx4f_ASAP7_75t_L g176 ( .A(n_123), .Y(n_176) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_123), .A2(n_240), .B(n_248), .Y(n_239) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_123), .A2(n_240), .B(n_248), .Y(n_285) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_123), .A2(n_240), .B(n_248), .Y(n_290) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_123), .Y(n_599) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g264 ( .A(n_124), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_124), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g190 ( .A(n_125), .Y(n_190) );
OAI21x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_139), .B(n_146), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_133), .B(n_136), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_130), .B(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
INVx1_ASAP7_75t_L g225 ( .A(n_131), .Y(n_225) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_132), .Y(n_135) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_132), .Y(n_142) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_132), .Y(n_162) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
INVx1_ASAP7_75t_L g203 ( .A(n_132), .Y(n_203) );
INVx1_ASAP7_75t_L g276 ( .A(n_134), .Y(n_276) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
INVx2_ASAP7_75t_L g244 ( .A(n_135), .Y(n_244) );
INVx2_ASAP7_75t_L g522 ( .A(n_135), .Y(n_522) );
INVx1_ASAP7_75t_L g565 ( .A(n_135), .Y(n_565) );
INVx2_ASAP7_75t_L g580 ( .A(n_135), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_135), .B(n_582), .Y(n_581) );
OAI21xp33_ASAP7_75t_L g165 ( .A1(n_136), .A2(n_166), .B(n_169), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_136), .A2(n_187), .B1(n_635), .B2(n_636), .Y(n_634) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_137), .Y(n_136) );
INVx3_ASAP7_75t_L g183 ( .A(n_137), .Y(n_183) );
BUFx2_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_137), .A2(n_259), .B(n_260), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_137), .A2(n_549), .B(n_550), .Y(n_548) );
AOI21x1_ASAP7_75t_L g610 ( .A1(n_137), .A2(n_611), .B(n_612), .Y(n_610) );
BUFx12f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx5_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
INVx5_ASAP7_75t_L g164 ( .A(n_138), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_138), .A2(n_275), .B(n_276), .C(n_277), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_138), .A2(n_563), .B1(n_564), .B2(n_566), .Y(n_562) );
OAI321xp33_ASAP7_75t_L g571 ( .A1(n_138), .A2(n_142), .A3(n_522), .B1(n_572), .B2(n_573), .C(n_574), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_143), .B(n_144), .Y(n_139) );
INVx2_ASAP7_75t_L g206 ( .A(n_141), .Y(n_206) );
INVx2_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_142), .B(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g218 ( .A(n_142), .Y(n_218) );
INVx2_ASAP7_75t_L g223 ( .A(n_142), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_142), .A2(n_145), .B(n_546), .C(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_145), .A2(n_246), .B(n_247), .Y(n_245) );
AOI21x1_ASAP7_75t_L g255 ( .A1(n_145), .A2(n_256), .B(n_257), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_146), .A2(n_178), .B(n_184), .Y(n_177) );
OAI21x1_ASAP7_75t_L g215 ( .A1(n_146), .A2(n_216), .B(n_220), .Y(n_215) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_146), .A2(n_241), .B(n_245), .Y(n_240) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_146), .A2(n_274), .B(n_278), .Y(n_273) );
AO31x2_ASAP7_75t_L g517 ( .A1(n_146), .A2(n_154), .A3(n_518), .B(n_524), .Y(n_517) );
INVx8_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_147), .A2(n_156), .B(n_165), .Y(n_155) );
NOR2xp67_ASAP7_75t_L g194 ( .A(n_147), .B(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g530 ( .A(n_147), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_147), .A2(n_574), .B(n_584), .Y(n_583) );
INVx8_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx2_ASAP7_75t_L g261 ( .A(n_148), .Y(n_261) );
INVx1_ASAP7_75t_L g553 ( .A(n_148), .Y(n_553) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_148), .A2(n_558), .B(n_562), .Y(n_557) );
OAI21x1_ASAP7_75t_L g588 ( .A1(n_148), .A2(n_589), .B(n_593), .Y(n_588) );
INVx1_ASAP7_75t_L g469 ( .A(n_151), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_191), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_174), .Y(n_152) );
INVx1_ASAP7_75t_L g307 ( .A(n_153), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_153), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_SL g351 ( .A(n_153), .Y(n_351) );
AO21x2_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_173), .Y(n_153) );
INVx3_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_154), .A2(n_155), .B(n_173), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_163), .Y(n_156) );
NOR2xp67_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx5_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
CKINVDCx6p67_ASAP7_75t_R g187 ( .A(n_164), .Y(n_187) );
AOI21x1_ASAP7_75t_L g558 ( .A1(n_164), .A2(n_559), .B(n_560), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_164), .A2(n_576), .B(n_581), .Y(n_575) );
AOI21x1_ASAP7_75t_L g607 ( .A1(n_164), .A2(n_608), .B(n_609), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
NOR2xp33_ASAP7_75t_SL g169 ( .A(n_170), .B(n_172), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_170), .B(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g520 ( .A(n_171), .Y(n_520) );
INVx2_ASAP7_75t_L g551 ( .A(n_171), .Y(n_551) );
INVx2_ASAP7_75t_L g561 ( .A(n_171), .Y(n_561) );
OR2x2_ASAP7_75t_L g302 ( .A(n_174), .B(n_303), .Y(n_302) );
BUFx3_ASAP7_75t_L g356 ( .A(n_174), .Y(n_356) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g235 ( .A(n_175), .Y(n_235) );
AND2x2_ASAP7_75t_L g333 ( .A(n_175), .B(n_232), .Y(n_333) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_188), .Y(n_175) );
OAI21x1_ASAP7_75t_L g214 ( .A1(n_176), .A2(n_215), .B(n_226), .Y(n_214) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_176), .A2(n_273), .B(n_281), .Y(n_272) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_176), .A2(n_273), .B(n_281), .Y(n_295) );
OA21x2_ASAP7_75t_L g314 ( .A1(n_176), .A2(n_215), .B(n_226), .Y(n_314) );
O2A1O1Ixp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_182), .C(n_183), .Y(n_178) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
O2A1O1Ixp5_ASAP7_75t_L g220 ( .A1(n_183), .A2(n_221), .B(n_222), .C(n_224), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_183), .A2(n_222), .B(n_279), .C(n_280), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_183), .A2(n_187), .B1(n_519), .B2(n_521), .Y(n_518) );
OA22x2_ASAP7_75t_L g531 ( .A1(n_183), .A2(n_187), .B1(n_532), .B2(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_187), .A2(n_217), .B(n_219), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_187), .A2(n_242), .B(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g529 ( .A(n_189), .Y(n_529) );
BUFx5_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g525 ( .A(n_190), .Y(n_525) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_190), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_191), .B(n_235), .Y(n_496) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVxp67_ASAP7_75t_SL g300 ( .A(n_192), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_192), .B(n_235), .Y(n_341) );
INVx1_ASAP7_75t_L g366 ( .A(n_192), .Y(n_366) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g231 ( .A(n_193), .Y(n_231) );
AOI21x1_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_196), .B(n_209), .Y(n_193) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_195), .A2(n_557), .B(n_567), .Y(n_556) );
OAI21x1_ASAP7_75t_L g605 ( .A1(n_195), .A2(n_606), .B(n_615), .Y(n_605) );
OAI21x1_ASAP7_75t_L g662 ( .A1(n_195), .A2(n_606), .B(n_615), .Y(n_662) );
OAI21x1_ASAP7_75t_L g697 ( .A1(n_195), .A2(n_557), .B(n_567), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_205), .Y(n_196) );
OAI21x1_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_200), .B(n_204), .Y(n_197) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g523 ( .A(n_203), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g593 ( .A1(n_206), .A2(n_594), .B(n_595), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_210), .A2(n_453), .B1(n_456), .B2(n_457), .Y(n_452) );
INVx1_ASAP7_75t_L g456 ( .A(n_210), .Y(n_456) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2x1_ASAP7_75t_L g336 ( .A(n_211), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g284 ( .A(n_212), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g324 ( .A(n_212), .B(n_285), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_212), .B(n_313), .Y(n_362) );
OR2x2_ASAP7_75t_L g414 ( .A(n_212), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g296 ( .A(n_213), .B(n_252), .Y(n_296) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g251 ( .A(n_214), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_229), .B(n_233), .Y(n_228) );
INVx1_ASAP7_75t_L g408 ( .A(n_229), .Y(n_408) );
NAND2xp67_ASAP7_75t_L g439 ( .A(n_229), .B(n_326), .Y(n_439) );
INVx1_ASAP7_75t_L g482 ( .A(n_229), .Y(n_482) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
INVx1_ASAP7_75t_L g317 ( .A(n_230), .Y(n_317) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g268 ( .A(n_231), .B(n_232), .Y(n_268) );
INVx1_ASAP7_75t_L g309 ( .A(n_231), .Y(n_309) );
AND2x2_ASAP7_75t_L g350 ( .A(n_231), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g370 ( .A(n_234), .B(n_267), .Y(n_370) );
OR2x2_ASAP7_75t_L g398 ( .A(n_234), .B(n_299), .Y(n_398) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
INVx2_ASAP7_75t_L g375 ( .A(n_235), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_235), .B(n_307), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_249), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_238), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g355 ( .A(n_238), .B(n_356), .Y(n_355) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_238), .B(n_299), .C(n_305), .D(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g400 ( .A(n_238), .B(n_292), .Y(n_400) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g311 ( .A(n_239), .Y(n_311) );
AND2x2_ASAP7_75t_L g492 ( .A(n_239), .B(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g436 ( .A(n_249), .Y(n_436) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g305 ( .A(n_251), .B(n_293), .Y(n_305) );
BUFx2_ASAP7_75t_L g330 ( .A(n_251), .Y(n_330) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_251), .B(n_391), .Y(n_431) );
INVx2_ASAP7_75t_L g313 ( .A(n_252), .Y(n_313) );
OR2x2_ASAP7_75t_L g427 ( .A(n_252), .B(n_272), .Y(n_427) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_258), .B(n_261), .Y(n_254) );
OAI21x1_ASAP7_75t_L g606 ( .A1(n_261), .A2(n_607), .B(n_610), .Y(n_606) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_266), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_268), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g385 ( .A(n_268), .B(n_301), .Y(n_385) );
AND2x2_ASAP7_75t_L g478 ( .A(n_268), .B(n_454), .Y(n_478) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_283), .Y(n_269) );
INVx2_ASAP7_75t_L g485 ( .A(n_270), .Y(n_485) );
BUFx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_271), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_282), .Y(n_271) );
INVx1_ASAP7_75t_L g329 ( .A(n_272), .Y(n_329) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp33_ASAP7_75t_R g373 ( .A(n_284), .B(n_328), .Y(n_373) );
INVx1_ASAP7_75t_L g472 ( .A(n_284), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_285), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g379 ( .A(n_285), .Y(n_379) );
OAI21xp33_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_297), .B(n_304), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
O2A1O1Ixp5_ASAP7_75t_L g358 ( .A1(n_288), .A2(n_359), .B(n_363), .C(n_369), .Y(n_358) );
NOR2x1p5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g335 ( .A(n_290), .Y(n_335) );
BUFx2_ASAP7_75t_L g346 ( .A(n_290), .Y(n_346) );
INVx2_ASAP7_75t_SL g415 ( .A(n_290), .Y(n_415) );
INVx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
AND2x4_ASAP7_75t_L g321 ( .A(n_293), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_295), .Y(n_361) );
AND2x2_ASAP7_75t_L g344 ( .A(n_296), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g491 ( .A(n_296), .Y(n_491) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g474 ( .A(n_299), .Y(n_474) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g395 ( .A(n_302), .Y(n_395) );
INVx1_ASAP7_75t_SL g405 ( .A(n_302), .Y(n_405) );
OR2x2_ASAP7_75t_L g441 ( .A(n_302), .B(n_365), .Y(n_441) );
OR2x2_ASAP7_75t_L g463 ( .A(n_302), .B(n_451), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B1(n_310), .B2(n_315), .Y(n_304) );
INVx2_ASAP7_75t_L g397 ( .A(n_305), .Y(n_397) );
INVx1_ASAP7_75t_L g347 ( .A(n_306), .Y(n_347) );
AND2x4_ASAP7_75t_L g429 ( .A(n_306), .B(n_375), .Y(n_429) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
BUFx2_ASAP7_75t_SL g458 ( .A(n_307), .Y(n_458) );
AND2x4_ASAP7_75t_L g332 ( .A(n_308), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g423 ( .A(n_308), .Y(n_423) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
OR2x6_ASAP7_75t_SL g426 ( .A(n_311), .B(n_427), .Y(n_426) );
OAI211xp5_ASAP7_75t_L g476 ( .A1(n_311), .A2(n_477), .B(n_480), .C(n_488), .Y(n_476) );
AND2x2_ASAP7_75t_L g483 ( .A(n_311), .B(n_431), .Y(n_483) );
INVx2_ASAP7_75t_L g392 ( .A(n_312), .Y(n_392) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx2_ASAP7_75t_L g322 ( .A(n_313), .Y(n_322) );
INVx2_ASAP7_75t_L g380 ( .A(n_314), .Y(n_380) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx2_ASAP7_75t_L g401 ( .A(n_317), .Y(n_401) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_318), .Y(n_357) );
INVx2_ASAP7_75t_L g376 ( .A(n_318), .Y(n_376) );
OR2x2_ASAP7_75t_L g433 ( .A(n_318), .B(n_366), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_342), .Y(n_319) );
OAI332xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_323), .A3(n_325), .B1(n_327), .B2(n_330), .B3(n_331), .C1(n_334), .C2(n_338), .Y(n_320) );
INVx2_ASAP7_75t_L g393 ( .A(n_321), .Y(n_393) );
AND2x4_ASAP7_75t_SL g353 ( .A(n_322), .B(n_337), .Y(n_353) );
BUFx2_ASAP7_75t_L g460 ( .A(n_322), .Y(n_460) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI311xp33_ASAP7_75t_L g369 ( .A1(n_324), .A2(n_370), .A3(n_371), .B1(n_372), .C1(n_382), .Y(n_369) );
AND2x2_ASAP7_75t_L g386 ( .A(n_324), .B(n_387), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_325), .A2(n_389), .B1(n_393), .B2(n_394), .Y(n_388) );
AND2x4_ASAP7_75t_L g349 ( .A(n_326), .B(n_350), .Y(n_349) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g391 ( .A(n_329), .Y(n_391) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_330), .B(n_355), .C(n_357), .Y(n_354) );
AOI22xp33_ASAP7_75t_SL g430 ( .A1(n_330), .A2(n_381), .B1(n_431), .B2(n_432), .Y(n_430) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
OR2x2_ASAP7_75t_L g425 ( .A(n_335), .B(n_392), .Y(n_425) );
BUFx2_ASAP7_75t_L g371 ( .A(n_337), .Y(n_371) );
INVx1_ASAP7_75t_L g387 ( .A(n_337), .Y(n_387) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
OR2x2_ASAP7_75t_L g498 ( .A(n_339), .B(n_496), .Y(n_498) );
INVx1_ASAP7_75t_L g455 ( .A(n_340), .Y(n_455) );
INVx1_ASAP7_75t_L g411 ( .A(n_341), .Y(n_411) );
OAI221xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_347), .B1(n_348), .B2(n_352), .C(n_354), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g381 ( .A(n_350), .B(n_356), .Y(n_381) );
AND2x2_ASAP7_75t_L g404 ( .A(n_350), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g464 ( .A(n_350), .Y(n_464) );
INVx2_ASAP7_75t_L g437 ( .A(n_353), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_353), .A2(n_460), .B1(n_478), .B2(n_479), .Y(n_477) );
AND2x2_ASAP7_75t_L g494 ( .A(n_357), .B(n_495), .Y(n_494) );
INVx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_361), .Y(n_413) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_361), .Y(n_471) );
INVx1_ASAP7_75t_L g493 ( .A(n_362), .Y(n_493) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_377), .B2(n_381), .Y(n_372) );
INVx3_ASAP7_75t_L g475 ( .A(n_374), .Y(n_475) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
AOI321xp33_ASAP7_75t_L g399 ( .A1(n_375), .A2(n_400), .A3(n_401), .B1(n_402), .B2(n_404), .C(n_406), .Y(n_399) );
OR2x2_ASAP7_75t_L g407 ( .A(n_375), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g448 ( .A(n_375), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g410 ( .A(n_376), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g403 ( .A(n_378), .Y(n_403) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_378), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
AOI211xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B(n_388), .C(n_396), .Y(n_384) );
AOI222xp33_ASAP7_75t_L g488 ( .A1(n_385), .A2(n_489), .B1(n_492), .B2(n_494), .C1(n_497), .C2(n_916), .Y(n_488) );
NAND2x1_ASAP7_75t_L g428 ( .A(n_386), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g402 ( .A(n_387), .B(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI32xp33_ASAP7_75t_L g473 ( .A1(n_392), .A2(n_427), .A3(n_463), .B1(n_474), .B2(n_475), .Y(n_473) );
NOR2xp67_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g487 ( .A(n_398), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_401), .B(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_403), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_409), .B(n_412), .Y(n_406) );
INVx1_ASAP7_75t_L g479 ( .A(n_407), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_409), .A2(n_441), .B1(n_442), .B2(n_445), .Y(n_440) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g444 ( .A(n_414), .Y(n_444) );
INVx1_ASAP7_75t_L g451 ( .A(n_415), .Y(n_451) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_476), .Y(n_416) );
NAND4xp75_ASAP7_75t_L g417 ( .A(n_418), .B(n_434), .C(n_447), .D(n_465), .Y(n_417) );
AND3x1_ASAP7_75t_L g418 ( .A(n_419), .B(n_428), .C(n_430), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_424), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
NAND2xp33_ASAP7_75t_SL g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx2_ASAP7_75t_L g443 ( .A(n_427), .Y(n_443) );
OR2x2_ASAP7_75t_L g450 ( .A(n_427), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_438), .B(n_440), .Y(n_434) );
NAND2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND2x1_ASAP7_75t_SL g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI21x1_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_452), .B(n_459), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NOR2x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NOR2x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_470), .B(n_473), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_499), .A2(n_506), .B1(n_508), .B2(n_864), .Y(n_863) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g506 ( .A(n_501), .B(n_502), .Y(n_506) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g904 ( .A(n_504), .B(n_905), .C(n_908), .Y(n_904) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2x1_ASAP7_75t_L g510 ( .A(n_511), .B(n_761), .Y(n_510) );
NAND4xp25_ASAP7_75t_L g511 ( .A(n_512), .B(n_665), .C(n_712), .D(n_749), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_602), .B(n_616), .Y(n_512) );
AO22x1_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_554), .B1(n_585), .B2(n_601), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_536), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_515), .B(n_537), .Y(n_678) );
AND2x2_ASAP7_75t_L g781 ( .A(n_515), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_516), .B(n_733), .Y(n_732) );
INVxp67_ASAP7_75t_L g817 ( .A(n_516), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_527), .Y(n_516) );
AND2x2_ASAP7_75t_L g597 ( .A(n_517), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g623 ( .A(n_517), .Y(n_623) );
INVx1_ASAP7_75t_L g644 ( .A(n_517), .Y(n_644) );
INVx1_ASAP7_75t_L g674 ( .A(n_517), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g543 ( .A(n_525), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_525), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g672 ( .A(n_527), .Y(n_672) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_527), .Y(n_690) );
INVx1_ASAP7_75t_L g717 ( .A(n_527), .Y(n_717) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_527), .Y(n_747) );
INVx1_ASAP7_75t_L g796 ( .A(n_527), .Y(n_796) );
OAI21x1_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_531), .B(n_534), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
OA21x2_ASAP7_75t_L g598 ( .A1(n_531), .A2(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVxp67_ASAP7_75t_L g600 ( .A(n_535), .Y(n_600) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g812 ( .A(n_537), .B(n_597), .Y(n_812) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NOR2xp67_ASAP7_75t_L g643 ( .A(n_538), .B(n_644), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g791 ( .A(n_538), .B(n_716), .C(n_792), .Y(n_791) );
AND2x2_ASAP7_75t_L g795 ( .A(n_538), .B(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g619 ( .A(n_539), .B(n_598), .Y(n_619) );
AND2x2_ASAP7_75t_L g718 ( .A(n_539), .B(n_682), .Y(n_718) );
AND2x2_ASAP7_75t_L g726 ( .A(n_539), .B(n_644), .Y(n_726) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g676 ( .A(n_540), .B(n_587), .Y(n_676) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g650 ( .A(n_541), .Y(n_650) );
AND2x2_ASAP7_75t_L g760 ( .A(n_541), .B(n_587), .Y(n_760) );
NAND2x1p5_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
OAI21x1_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_548), .B(n_552), .Y(n_544) );
AND2x2_ASAP7_75t_L g753 ( .A(n_554), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_568), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_555), .B(n_663), .Y(n_668) );
INVx1_ASAP7_75t_L g736 ( .A(n_555), .Y(n_736) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g627 ( .A(n_556), .Y(n_627) );
INVxp67_ASAP7_75t_L g591 ( .A(n_561), .Y(n_591) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_565), .B(n_613), .Y(n_612) );
BUFx2_ASAP7_75t_L g601 ( .A(n_568), .Y(n_601) );
AND2x4_ASAP7_75t_L g778 ( .A(n_568), .B(n_723), .Y(n_778) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_569), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g730 ( .A(n_569), .B(n_662), .Y(n_730) );
AND2x2_ASAP7_75t_L g844 ( .A(n_569), .B(n_739), .Y(n_844) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g630 ( .A(n_570), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g641 ( .A(n_570), .Y(n_641) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_575), .B(n_583), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI32xp33_ASAP7_75t_L g653 ( .A1(n_585), .A2(n_647), .A3(n_654), .B1(n_655), .B2(n_658), .Y(n_653) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_597), .Y(n_585) );
NOR2xp67_ASAP7_75t_L g620 ( .A(n_586), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g648 ( .A(n_586), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_586), .B(n_674), .Y(n_711) );
OAI32xp33_ASAP7_75t_L g763 ( .A1(n_586), .A2(n_671), .A3(n_764), .B1(n_767), .B2(n_769), .Y(n_763) );
NOR3xp33_ASAP7_75t_L g798 ( .A(n_586), .B(n_664), .C(n_799), .Y(n_798) );
BUFx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_592), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_597), .B(n_748), .Y(n_853) );
AND2x2_ASAP7_75t_L g645 ( .A(n_598), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g654 ( .A(n_601), .Y(n_654) );
INVx1_ASAP7_75t_L g822 ( .A(n_601), .Y(n_822) );
OR2x2_ASAP7_75t_L g849 ( .A(n_602), .B(n_765), .Y(n_849) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g625 ( .A(n_603), .B(n_626), .Y(n_625) );
BUFx2_ASAP7_75t_L g669 ( .A(n_603), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_603), .B(n_626), .Y(n_766) );
AND2x2_ASAP7_75t_L g788 ( .A(n_603), .B(n_689), .Y(n_788) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g652 ( .A(n_604), .B(n_631), .Y(n_652) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_604), .Y(n_842) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g704 ( .A(n_605), .Y(n_704) );
INVx4_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_653), .Y(n_616) );
AOI322xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_624), .A3(n_628), .B1(n_639), .B2(n_642), .C1(n_647), .C2(n_651), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx2_ASAP7_75t_L g710 ( .A(n_619), .Y(n_710) );
AND2x2_ASAP7_75t_L g837 ( .A(n_619), .B(n_681), .Y(n_837) );
INVxp67_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g826 ( .A(n_622), .B(n_650), .Y(n_826) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x4_ASAP7_75t_L g649 ( .A(n_623), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g681 ( .A(n_623), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_625), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g640 ( .A(n_626), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g830 ( .A(n_626), .B(n_735), .Y(n_830) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_SL g664 ( .A(n_627), .Y(n_664) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_629), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g722 ( .A(n_630), .B(n_723), .Y(n_722) );
BUFx3_ASAP7_75t_L g786 ( .A(n_630), .Y(n_786) );
AND2x2_ASAP7_75t_L g807 ( .A(n_630), .B(n_724), .Y(n_807) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_631), .Y(n_657) );
INVx2_ASAP7_75t_L g663 ( .A(n_631), .Y(n_663) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g739 ( .A(n_632), .Y(n_739) );
AOI21x1_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_637), .Y(n_632) );
AND2x2_ASAP7_75t_L g696 ( .A(n_641), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g707 ( .A(n_641), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g765 ( .A(n_641), .B(n_739), .Y(n_765) );
INVxp67_ASAP7_75t_SL g780 ( .A(n_641), .Y(n_780) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g757 ( .A(n_644), .Y(n_757) );
AND2x4_ASAP7_75t_L g825 ( .A(n_645), .B(n_826), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_645), .B(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g682 ( .A(n_646), .Y(n_682) );
AND2x4_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx2_ASAP7_75t_L g691 ( .A(n_649), .Y(n_691) );
AND2x2_ASAP7_75t_L g727 ( .A(n_649), .B(n_717), .Y(n_727) );
BUFx2_ASAP7_75t_L g790 ( .A(n_649), .Y(n_790) );
INVx1_ASAP7_75t_L g847 ( .A(n_649), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_650), .B(n_682), .Y(n_733) );
INVx2_ASAP7_75t_L g684 ( .A(n_652), .Y(n_684) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g794 ( .A1(n_656), .A2(n_726), .B1(n_795), .B2(n_797), .C(n_798), .Y(n_794) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_657), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g797 ( .A(n_657), .Y(n_797) );
INVx1_ASAP7_75t_L g686 ( .A(n_658), .Y(n_686) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_664), .Y(n_659) );
INVx2_ASAP7_75t_L g771 ( .A(n_660), .Y(n_771) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVx2_ASAP7_75t_L g699 ( .A(n_661), .Y(n_699) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g700 ( .A(n_663), .Y(n_700) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_663), .Y(n_729) );
AND2x2_ASAP7_75t_L g683 ( .A(n_664), .B(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g719 ( .A(n_664), .B(n_698), .Y(n_719) );
AND2x2_ASAP7_75t_L g803 ( .A(n_664), .B(n_706), .Y(n_803) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_670), .B1(n_677), .B2(n_683), .C(n_685), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_668), .B(n_780), .Y(n_779) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
OR2x2_ASAP7_75t_L g679 ( .A(n_671), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g767 ( .A(n_671), .B(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g725 ( .A(n_672), .B(n_726), .Y(n_725) );
NOR2x1_ASAP7_75t_L g821 ( .A(n_672), .B(n_757), .Y(n_821) );
NOR2x1_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g693 ( .A(n_674), .Y(n_693) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_674), .Y(n_714) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g740 ( .A(n_676), .B(n_717), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NOR2x1p5_ASAP7_75t_L g827 ( .A(n_680), .B(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g689 ( .A(n_682), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_684), .B(n_696), .Y(n_815) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_692), .B2(n_694), .C(n_701), .Y(n_685) );
OAI222xp33_ASAP7_75t_L g850 ( .A1(n_687), .A2(n_752), .B1(n_851), .B2(n_852), .C1(n_853), .C2(n_854), .Y(n_850) );
OR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_691), .Y(n_687) );
OR2x2_ASAP7_75t_L g692 ( .A(n_688), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
OR2x6_ASAP7_75t_L g835 ( .A(n_691), .B(n_796), .Y(n_835) );
INVx2_ASAP7_75t_L g808 ( .A(n_692), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_698), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_695), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g708 ( .A(n_697), .Y(n_708) );
INVx2_ASAP7_75t_L g724 ( .A(n_697), .Y(n_724) );
INVx1_ASAP7_75t_L g752 ( .A(n_698), .Y(n_752) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx2_ASAP7_75t_L g706 ( .A(n_699), .Y(n_706) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_699), .Y(n_754) );
AND2x2_ASAP7_75t_L g819 ( .A(n_699), .B(n_718), .Y(n_819) );
AND2x2_ASAP7_75t_L g735 ( .A(n_700), .B(n_704), .Y(n_735) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_705), .B(n_709), .Y(n_701) );
BUFx2_ASAP7_75t_L g793 ( .A(n_704), .Y(n_793) );
INVxp67_ASAP7_75t_SL g855 ( .A(n_704), .Y(n_855) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
AND2x2_ASAP7_75t_L g737 ( .A(n_707), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g770 ( .A(n_707), .Y(n_770) );
NOR2x1p5_ASAP7_75t_SL g709 ( .A(n_710), .B(n_711), .Y(n_709) );
AOI211xp5_ASAP7_75t_SL g712 ( .A1(n_713), .A2(n_719), .B(n_720), .C(n_741), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx2_ASAP7_75t_L g806 ( .A(n_715), .Y(n_806) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
AO22x1_ASAP7_75t_L g820 ( .A1(n_716), .A2(n_821), .B1(n_822), .B2(n_823), .Y(n_820) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g768 ( .A(n_718), .Y(n_768) );
AND2x2_ASAP7_75t_L g831 ( .A(n_718), .B(n_817), .Y(n_831) );
INVx1_ASAP7_75t_L g743 ( .A(n_719), .Y(n_743) );
NAND2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_731), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_725), .B1(n_727), .B2(n_728), .Y(n_721) );
INVx2_ASAP7_75t_SL g742 ( .A(n_722), .Y(n_742) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g848 ( .A(n_725), .Y(n_848) );
AND2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g799 ( .A(n_730), .Y(n_799) );
AOI32xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_734), .A3(n_736), .B1(n_737), .B2(n_740), .Y(n_731) );
INVx1_ASAP7_75t_L g748 ( .A(n_733), .Y(n_748) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx2_ASAP7_75t_L g774 ( .A(n_735), .Y(n_774) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g805 ( .A(n_740), .Y(n_805) );
AOI21xp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B(n_744), .Y(n_741) );
OAI321xp33_ASAP7_75t_L g784 ( .A1(n_742), .A2(n_785), .A3(n_787), .B1(n_789), .B2(n_791), .C(n_794), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_748), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND2x1p5_ASAP7_75t_L g759 ( .A(n_746), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI21xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_753), .B(n_755), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AND2x4_ASAP7_75t_L g755 ( .A(n_756), .B(n_758), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g783 ( .A(n_760), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_809), .Y(n_761) );
NOR4xp25_ASAP7_75t_L g762 ( .A(n_763), .B(n_772), .C(n_784), .D(n_800), .Y(n_762) );
OR2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVx2_ASAP7_75t_L g802 ( .A(n_765), .Y(n_802) );
OR2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
INVx2_ASAP7_75t_L g823 ( .A(n_770), .Y(n_823) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
A2O1A1Ixp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .B(n_779), .C(n_781), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI21xp33_ASAP7_75t_L g829 ( .A1(n_776), .A2(n_830), .B(n_831), .Y(n_829) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx4_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
OAI21xp33_ASAP7_75t_L g834 ( .A1(n_785), .A2(n_835), .B(n_836), .Y(n_834) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_786), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g813 ( .A(n_792), .B(n_807), .Y(n_813) );
INVxp67_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_L g828 ( .A(n_795), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_797), .A2(n_802), .B1(n_825), .B2(n_827), .Y(n_824) );
AO22x1_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_804), .B1(n_807), .B2(n_808), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g852 ( .A(n_802), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
NOR3xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_832), .C(n_850), .Y(n_809) );
NAND4xp25_ASAP7_75t_L g810 ( .A(n_811), .B(n_818), .C(n_824), .D(n_829), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_813), .B1(n_814), .B2(n_816), .Y(n_811) );
INVxp67_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
BUFx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_830), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g851 ( .A(n_831), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_838), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_845), .B1(n_848), .B2(n_849), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_841), .B(n_843), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx4_ASAP7_75t_SL g856 ( .A(n_857), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_857), .B(n_863), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_861), .Y(n_860) );
NOR2x1_ASAP7_75t_R g867 ( .A(n_861), .B(n_868), .Y(n_867) );
INVx2_ASAP7_75t_SL g898 ( .A(n_861), .Y(n_898) );
OAI21xp5_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_871), .B(n_888), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx4_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
BUFx6f_ASAP7_75t_L g892 ( .A(n_869), .Y(n_892) );
BUFx6f_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_881), .B1(n_882), .B2(n_887), .Y(n_871) );
OAI21xp5_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_878), .B(n_880), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g873 ( .A(n_874), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_882), .Y(n_881) );
CKINVDCx5p33_ASAP7_75t_R g886 ( .A(n_883), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_884), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_893), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
BUFx6f_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
BUFx12f_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
OR2x2_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_901), .Y(n_900) );
BUFx12f_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx4_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
BUFx4f_ASAP7_75t_L g914 ( .A(n_903), .Y(n_914) );
AND2x2_ASAP7_75t_SL g903 ( .A(n_904), .B(n_909), .Y(n_903) );
INVx4_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .Y(n_911) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
endmodule