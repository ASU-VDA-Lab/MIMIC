module real_aes_7770_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_756;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g169 ( .A1(n_0), .A2(n_170), .B(n_173), .C(n_177), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_1), .B(n_161), .Y(n_180) );
INVx1_ASAP7_75t_L g444 ( .A(n_2), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_3), .B(n_171), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_4), .A2(n_134), .B(n_137), .C(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_5), .A2(n_129), .B(n_561), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_6), .A2(n_129), .B(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_7), .B(n_161), .Y(n_567) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_8), .A2(n_163), .B(n_235), .Y(n_234) );
AND2x6_ASAP7_75t_L g134 ( .A(n_9), .B(n_135), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_10), .A2(n_134), .B(n_137), .C(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g528 ( .A(n_11), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_12), .B(n_39), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_13), .B(n_176), .Y(n_539) );
INVx1_ASAP7_75t_L g155 ( .A(n_14), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_15), .B(n_171), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_16), .A2(n_172), .B(n_547), .C(n_549), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_17), .B(n_161), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_18), .B(n_149), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g136 ( .A1(n_19), .A2(n_137), .B(n_140), .C(n_148), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g576 ( .A1(n_20), .A2(n_175), .B(n_243), .C(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_21), .B(n_176), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_22), .B(n_176), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_23), .Y(n_509) );
INVx1_ASAP7_75t_L g489 ( .A(n_24), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_25), .A2(n_137), .B(n_148), .C(n_238), .Y(n_237) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_26), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_27), .Y(n_535) );
INVx1_ASAP7_75t_L g503 ( .A(n_28), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_29), .A2(n_129), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g132 ( .A(n_30), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_31), .A2(n_187), .B(n_188), .C(n_192), .Y(n_186) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_32), .A2(n_104), .B1(n_450), .B2(n_459), .C1(n_761), .C2(n_766), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_32), .A2(n_33), .B1(n_108), .B2(n_109), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_32), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_33), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_34), .A2(n_175), .B(n_564), .C(n_566), .Y(n_563) );
INVxp67_ASAP7_75t_L g504 ( .A(n_35), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_36), .B(n_240), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_37), .A2(n_137), .B(n_148), .C(n_488), .Y(n_487) );
CKINVDCx14_ASAP7_75t_R g562 ( .A(n_38), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_40), .A2(n_177), .B(n_526), .C(n_527), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_41), .B(n_128), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_42), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_43), .B(n_171), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_44), .B(n_129), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_45), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_46), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_47), .A2(n_187), .B(n_192), .C(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g174 ( .A(n_48), .Y(n_174) );
INVx1_ASAP7_75t_L g218 ( .A(n_49), .Y(n_218) );
INVx1_ASAP7_75t_L g575 ( .A(n_50), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_51), .B(n_129), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_52), .Y(n_157) );
CKINVDCx14_ASAP7_75t_R g524 ( .A(n_53), .Y(n_524) );
AOI22xp5_ASAP7_75t_SL g460 ( .A1(n_54), .A2(n_442), .B1(n_461), .B2(n_758), .Y(n_460) );
INVx1_ASAP7_75t_L g135 ( .A(n_55), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_56), .B(n_129), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_57), .B(n_161), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_58), .A2(n_147), .B(n_203), .C(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g154 ( .A(n_59), .Y(n_154) );
INVx1_ASAP7_75t_SL g565 ( .A(n_60), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_61), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_62), .B(n_171), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_63), .B(n_161), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_64), .B(n_172), .Y(n_253) );
INVx1_ASAP7_75t_L g512 ( .A(n_65), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g167 ( .A(n_66), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_67), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_68), .A2(n_137), .B(n_192), .C(n_201), .Y(n_200) );
CKINVDCx16_ASAP7_75t_R g227 ( .A(n_69), .Y(n_227) );
INVx1_ASAP7_75t_L g458 ( .A(n_70), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_71), .A2(n_129), .B(n_523), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_72), .A2(n_94), .B1(n_114), .B2(n_115), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_72), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_73), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_74), .A2(n_102), .B1(n_471), .B2(n_472), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_74), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_75), .A2(n_129), .B(n_544), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_76), .A2(n_128), .B(n_499), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_77), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_78), .A2(n_468), .B1(n_469), .B2(n_470), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_78), .Y(n_468) );
INVx1_ASAP7_75t_L g545 ( .A(n_79), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_80), .B(n_145), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_81), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_82), .A2(n_129), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g548 ( .A(n_83), .Y(n_548) );
INVx2_ASAP7_75t_L g152 ( .A(n_84), .Y(n_152) );
INVx1_ASAP7_75t_L g538 ( .A(n_85), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_86), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_87), .B(n_176), .Y(n_254) );
OR2x2_ASAP7_75t_L g441 ( .A(n_88), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g463 ( .A(n_88), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_89), .A2(n_137), .B(n_192), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_90), .B(n_129), .Y(n_185) );
INVx1_ASAP7_75t_L g189 ( .A(n_91), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_92), .B(n_447), .Y(n_446) );
INVxp67_ASAP7_75t_L g230 ( .A(n_93), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_94), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_95), .A2(n_467), .B1(n_473), .B2(n_474), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_95), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_96), .B(n_163), .Y(n_529) );
INVx1_ASAP7_75t_L g202 ( .A(n_97), .Y(n_202) );
INVx1_ASAP7_75t_L g249 ( .A(n_98), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_99), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g578 ( .A(n_100), .Y(n_578) );
AND2x2_ASAP7_75t_L g220 ( .A(n_101), .B(n_151), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_102), .Y(n_471) );
OAI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_439), .B(n_446), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_107), .B1(n_110), .B2(n_111), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_108), .B(n_162), .Y(n_540) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_113), .B1(n_116), .B2(n_117), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_116), .A2(n_117), .B1(n_465), .B2(n_466), .Y(n_464) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_SL g117 ( .A(n_118), .B(n_394), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_329), .Y(n_118) );
NAND4xp25_ASAP7_75t_SL g119 ( .A(n_120), .B(n_274), .C(n_298), .D(n_321), .Y(n_119) );
AOI221xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_211), .B1(n_245), .B2(n_258), .C(n_261), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_181), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_123), .A2(n_159), .B1(n_212), .B2(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_123), .B(n_182), .Y(n_332) );
AND2x2_ASAP7_75t_L g351 ( .A(n_123), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_123), .B(n_335), .Y(n_421) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_159), .Y(n_123) );
AND2x2_ASAP7_75t_L g289 ( .A(n_124), .B(n_182), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_124), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g312 ( .A(n_124), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g317 ( .A(n_124), .B(n_160), .Y(n_317) );
INVx2_ASAP7_75t_L g349 ( .A(n_124), .Y(n_349) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_124), .Y(n_393) );
AND2x2_ASAP7_75t_L g410 ( .A(n_124), .B(n_287), .Y(n_410) );
INVx5_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g328 ( .A(n_125), .B(n_287), .Y(n_328) );
AND2x4_ASAP7_75t_L g342 ( .A(n_125), .B(n_159), .Y(n_342) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_125), .Y(n_346) );
AND2x2_ASAP7_75t_L g366 ( .A(n_125), .B(n_281), .Y(n_366) );
AND2x2_ASAP7_75t_L g416 ( .A(n_125), .B(n_183), .Y(n_416) );
AND2x2_ASAP7_75t_L g426 ( .A(n_125), .B(n_160), .Y(n_426) );
OR2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_156), .Y(n_125) );
AOI21xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_136), .B(n_149), .Y(n_126) );
BUFx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_134), .Y(n_129) );
NAND2x1p5_ASAP7_75t_L g250 ( .A(n_130), .B(n_134), .Y(n_250) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx1_ASAP7_75t_L g147 ( .A(n_131), .Y(n_147) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g138 ( .A(n_132), .Y(n_138) );
INVx1_ASAP7_75t_L g244 ( .A(n_132), .Y(n_244) );
INVx1_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_133), .Y(n_143) );
INVx3_ASAP7_75t_L g172 ( .A(n_133), .Y(n_172) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
INVx1_ASAP7_75t_L g240 ( .A(n_133), .Y(n_240) );
BUFx3_ASAP7_75t_L g148 ( .A(n_134), .Y(n_148) );
INVx4_ASAP7_75t_SL g179 ( .A(n_134), .Y(n_179) );
INVx5_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx3_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_138), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_144), .B(n_146), .Y(n_140) );
INVx2_ASAP7_75t_L g145 ( .A(n_142), .Y(n_145) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx4_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_145), .A2(n_189), .B(n_190), .C(n_191), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_145), .A2(n_191), .B(n_218), .C(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_145), .A2(n_512), .B(n_513), .C(n_514), .Y(n_511) );
O2A1O1Ixp5_ASAP7_75t_L g537 ( .A1(n_145), .A2(n_514), .B(n_538), .C(n_539), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_146), .A2(n_171), .B(n_489), .C(n_490), .Y(n_488) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_147), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_150), .B(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g158 ( .A(n_151), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_151), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_151), .A2(n_215), .B(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_151), .A2(n_250), .B(n_486), .C(n_487), .Y(n_485) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_151), .A2(n_522), .B(n_529), .Y(n_521) );
AND2x2_ASAP7_75t_SL g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AND2x2_ASAP7_75t_L g164 ( .A(n_152), .B(n_153), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_158), .A2(n_534), .B(n_540), .Y(n_533) );
AND2x2_ASAP7_75t_L g282 ( .A(n_159), .B(n_182), .Y(n_282) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_159), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_159), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g372 ( .A(n_159), .Y(n_372) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g260 ( .A(n_160), .B(n_197), .Y(n_260) );
AND2x2_ASAP7_75t_L g287 ( .A(n_160), .B(n_198), .Y(n_287) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_165), .B(n_180), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_162), .B(n_194), .Y(n_193) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_162), .A2(n_199), .B(n_209), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_162), .B(n_210), .Y(n_209) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_162), .A2(n_248), .B(n_255), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_162), .B(n_492), .Y(n_491) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_162), .A2(n_508), .B(n_515), .Y(n_507) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_163), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_163), .A2(n_236), .B(n_237), .Y(n_235) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g257 ( .A(n_164), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_SL g166 ( .A1(n_167), .A2(n_168), .B(n_169), .C(n_179), .Y(n_166) );
INVx2_ASAP7_75t_L g187 ( .A(n_168), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_168), .A2(n_179), .B(n_227), .C(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_SL g499 ( .A1(n_168), .A2(n_179), .B(n_500), .C(n_501), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_SL g523 ( .A1(n_168), .A2(n_179), .B(n_524), .C(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_SL g544 ( .A1(n_168), .A2(n_179), .B(n_545), .C(n_546), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g561 ( .A1(n_168), .A2(n_179), .B(n_562), .C(n_563), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_SL g574 ( .A1(n_168), .A2(n_179), .B(n_575), .C(n_576), .Y(n_574) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_171), .B(n_230), .Y(n_229) );
OAI22xp33_ASAP7_75t_L g502 ( .A1(n_171), .A2(n_204), .B1(n_503), .B2(n_504), .Y(n_502) );
INVx5_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_172), .B(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_175), .B(n_565), .Y(n_564) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g526 ( .A(n_176), .Y(n_526) );
INVx2_ASAP7_75t_L g514 ( .A(n_177), .Y(n_514) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_178), .Y(n_191) );
INVx1_ASAP7_75t_L g549 ( .A(n_178), .Y(n_549) );
INVx1_ASAP7_75t_L g192 ( .A(n_179), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_181), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_195), .Y(n_181) );
OR2x2_ASAP7_75t_L g313 ( .A(n_182), .B(n_196), .Y(n_313) );
AND2x2_ASAP7_75t_L g350 ( .A(n_182), .B(n_260), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_182), .B(n_281), .Y(n_361) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_182), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_182), .B(n_317), .Y(n_434) );
INVx5_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx2_ASAP7_75t_L g259 ( .A(n_183), .Y(n_259) );
AND2x2_ASAP7_75t_L g268 ( .A(n_183), .B(n_196), .Y(n_268) );
AND2x2_ASAP7_75t_L g384 ( .A(n_183), .B(n_279), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_183), .B(n_317), .Y(n_406) );
OR2x6_ASAP7_75t_L g183 ( .A(n_184), .B(n_193), .Y(n_183) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_196), .Y(n_352) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_197), .Y(n_304) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
BUFx2_ASAP7_75t_L g281 ( .A(n_198), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_208), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_205), .C(n_206), .Y(n_201) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_204), .B(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_204), .B(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g566 ( .A(n_207), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_221), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_212), .B(n_294), .Y(n_413) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_213), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g265 ( .A(n_213), .B(n_266), .Y(n_265) );
INVx5_ASAP7_75t_SL g273 ( .A(n_213), .Y(n_273) );
OR2x2_ASAP7_75t_L g296 ( .A(n_213), .B(n_266), .Y(n_296) );
OR2x2_ASAP7_75t_L g306 ( .A(n_213), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g369 ( .A(n_213), .B(n_223), .Y(n_369) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_213), .B(n_222), .Y(n_407) );
NOR4xp25_ASAP7_75t_L g428 ( .A(n_213), .B(n_349), .C(n_429), .D(n_430), .Y(n_428) );
AND2x2_ASAP7_75t_L g438 ( .A(n_213), .B(n_270), .Y(n_438) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_220), .Y(n_213) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g263 ( .A(n_222), .B(n_259), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_222), .B(n_265), .Y(n_432) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_232), .Y(n_222) );
OR2x2_ASAP7_75t_L g272 ( .A(n_223), .B(n_273), .Y(n_272) );
INVx3_ASAP7_75t_L g279 ( .A(n_223), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_223), .B(n_247), .Y(n_291) );
INVxp67_ASAP7_75t_L g294 ( .A(n_223), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_223), .B(n_266), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_223), .B(n_233), .Y(n_360) );
AND2x2_ASAP7_75t_L g375 ( .A(n_223), .B(n_270), .Y(n_375) );
OR2x2_ASAP7_75t_L g404 ( .A(n_223), .B(n_233), .Y(n_404) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_231), .Y(n_223) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_224), .A2(n_543), .B(n_550), .Y(n_542) );
OA21x2_ASAP7_75t_L g559 ( .A1(n_224), .A2(n_560), .B(n_567), .Y(n_559) );
OA21x2_ASAP7_75t_L g572 ( .A1(n_224), .A2(n_573), .B(n_579), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_232), .B(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_232), .B(n_273), .Y(n_412) );
OR2x2_ASAP7_75t_L g433 ( .A(n_232), .B(n_310), .Y(n_433) );
INVx1_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
OR2x2_ASAP7_75t_L g246 ( .A(n_233), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g270 ( .A(n_233), .B(n_266), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_233), .B(n_247), .Y(n_285) );
AND2x2_ASAP7_75t_L g355 ( .A(n_233), .B(n_279), .Y(n_355) );
AND2x2_ASAP7_75t_L g389 ( .A(n_233), .B(n_273), .Y(n_389) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_234), .B(n_273), .Y(n_292) );
AND2x2_ASAP7_75t_L g320 ( .A(n_234), .B(n_247), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_241), .B(n_242), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_242), .A2(n_253), .B(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_245), .B(n_328), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_246), .A2(n_335), .B1(n_371), .B2(n_388), .C(n_390), .Y(n_387) );
INVx5_ASAP7_75t_SL g266 ( .A(n_247), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_250), .B(n_251), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_250), .A2(n_509), .B(n_510), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_250), .A2(n_535), .B(n_536), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g497 ( .A(n_257), .Y(n_497) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
OAI33xp33_ASAP7_75t_L g286 ( .A1(n_259), .A2(n_287), .A3(n_288), .B1(n_290), .B2(n_293), .B3(n_297), .Y(n_286) );
OR2x2_ASAP7_75t_L g302 ( .A(n_259), .B(n_303), .Y(n_302) );
AOI322xp5_ASAP7_75t_L g411 ( .A1(n_259), .A2(n_328), .A3(n_335), .B1(n_412), .B2(n_413), .C1(n_414), .C2(n_417), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_259), .B(n_287), .Y(n_429) );
A2O1A1Ixp33_ASAP7_75t_SL g435 ( .A1(n_259), .A2(n_287), .B(n_436), .C(n_438), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g274 ( .A1(n_260), .A2(n_275), .B1(n_280), .B2(n_283), .C(n_286), .Y(n_274) );
INVx1_ASAP7_75t_L g367 ( .A(n_260), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_260), .B(n_416), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_264), .B1(n_267), .B2(n_269), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g344 ( .A(n_265), .B(n_279), .Y(n_344) );
AND2x2_ASAP7_75t_L g402 ( .A(n_265), .B(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g310 ( .A(n_266), .B(n_273), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_266), .B(n_279), .Y(n_338) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_268), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_268), .B(n_346), .Y(n_400) );
OAI321xp33_ASAP7_75t_L g419 ( .A1(n_268), .A2(n_341), .A3(n_420), .B1(n_421), .B2(n_422), .C(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g386 ( .A(n_269), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_270), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g325 ( .A(n_270), .B(n_273), .Y(n_325) );
AOI321xp33_ASAP7_75t_L g383 ( .A1(n_270), .A2(n_287), .A3(n_384), .B1(n_385), .B2(n_386), .C(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g300 ( .A(n_272), .B(n_285), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_273), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_273), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_273), .B(n_359), .Y(n_396) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g319 ( .A(n_277), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g284 ( .A(n_278), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g392 ( .A(n_279), .Y(n_392) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_282), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g315 ( .A(n_287), .Y(n_315) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_289), .B(n_324), .Y(n_373) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
OR2x2_ASAP7_75t_L g337 ( .A(n_292), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g382 ( .A(n_292), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_293), .A2(n_340), .B1(n_343), .B2(n_345), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g437 ( .A(n_296), .B(n_360), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_301), .B1(n_305), .B2(n_311), .C(n_314), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx2_ASAP7_75t_L g335 ( .A(n_304), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_SL g381 ( .A(n_307), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_309), .B(n_359), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_309), .A2(n_377), .B(n_379), .Y(n_376) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g422 ( .A(n_310), .B(n_404), .Y(n_422) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_SL g324 ( .A(n_313), .Y(n_324) );
AOI21xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B(n_318), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g368 ( .A(n_320), .B(n_369), .Y(n_368) );
INVxp67_ASAP7_75t_L g430 ( .A(n_320), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_325), .B(n_326), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_324), .B(n_342), .Y(n_378) );
INVxp67_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g399 ( .A(n_328), .Y(n_399) );
NAND5xp2_ASAP7_75t_L g329 ( .A(n_330), .B(n_347), .C(n_356), .D(n_376), .E(n_383), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_336), .C(n_339), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g371 ( .A(n_335), .Y(n_371) );
CKINVDCx16_ASAP7_75t_R g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_343), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g385 ( .A(n_345), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_351), .B(n_353), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_348), .A2(n_402), .B1(n_405), .B2(n_407), .C(n_408), .Y(n_401) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AOI321xp33_ASAP7_75t_L g356 ( .A1(n_349), .A2(n_357), .A3(n_361), .B1(n_362), .B2(n_368), .C(n_370), .Y(n_356) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g427 ( .A(n_361), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_363), .B(n_367), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g379 ( .A(n_364), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
NOR2xp67_ASAP7_75t_SL g391 ( .A(n_365), .B(n_372), .Y(n_391) );
AOI321xp33_ASAP7_75t_SL g423 ( .A1(n_368), .A2(n_424), .A3(n_425), .B1(n_426), .B2(n_427), .C(n_428), .Y(n_423) );
O2A1O1Ixp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B(n_373), .C(n_374), .Y(n_370) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_381), .B(n_389), .Y(n_418) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND3xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .C(n_393), .Y(n_390) );
NOR3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_419), .C(n_431), .Y(n_394) );
OAI211xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_397), .B(n_401), .C(n_411), .Y(n_395) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_399), .B(n_400), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_400), .A2(n_432), .B1(n_433), .B2(n_434), .C(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g420 ( .A(n_402), .Y(n_420) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g424 ( .A(n_422), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
CKINVDCx14_ASAP7_75t_R g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g449 ( .A(n_441), .Y(n_449) );
INVx1_ASAP7_75t_SL g765 ( .A(n_441), .Y(n_765) );
BUFx2_ASAP7_75t_L g768 ( .A(n_441), .Y(n_768) );
NOR2x2_ASAP7_75t_L g760 ( .A(n_442), .B(n_463), .Y(n_760) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
CKINVDCx6p67_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_SL g763 ( .A(n_455), .B(n_457), .Y(n_763) );
OA21x2_ASAP7_75t_L g767 ( .A1(n_455), .A2(n_456), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVxp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_464), .B1(n_475), .B2(n_477), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g476 ( .A(n_463), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_465), .A2(n_466), .B1(n_478), .B2(n_479), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g474 ( .A(n_467), .Y(n_474) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OR4x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_648), .C(n_695), .D(n_735), .Y(n_479) );
NAND3xp33_ASAP7_75t_SL g480 ( .A(n_481), .B(n_594), .C(n_623), .Y(n_480) );
AOI211xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_517), .B(n_551), .C(n_587), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_482), .A2(n_607), .B(n_624), .C(n_628), .Y(n_623) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_493), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_484), .B(n_586), .Y(n_585) );
INVx3_ASAP7_75t_SL g590 ( .A(n_484), .Y(n_590) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_484), .Y(n_602) );
AND2x4_ASAP7_75t_L g606 ( .A(n_484), .B(n_558), .Y(n_606) );
AND2x2_ASAP7_75t_L g617 ( .A(n_484), .B(n_507), .Y(n_617) );
OR2x2_ASAP7_75t_L g641 ( .A(n_484), .B(n_554), .Y(n_641) );
AND2x2_ASAP7_75t_L g654 ( .A(n_484), .B(n_559), .Y(n_654) );
AND2x2_ASAP7_75t_L g694 ( .A(n_484), .B(n_680), .Y(n_694) );
AND2x2_ASAP7_75t_L g701 ( .A(n_484), .B(n_664), .Y(n_701) );
AND2x2_ASAP7_75t_L g731 ( .A(n_484), .B(n_494), .Y(n_731) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_491), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_493), .B(n_658), .Y(n_670) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_506), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_494), .B(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g608 ( .A(n_494), .B(n_506), .Y(n_608) );
BUFx3_ASAP7_75t_L g616 ( .A(n_494), .Y(n_616) );
OR2x2_ASAP7_75t_L g637 ( .A(n_494), .B(n_520), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_494), .B(n_658), .Y(n_748) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .B(n_505), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_496), .A2(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g555 ( .A(n_498), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_505), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_506), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g601 ( .A(n_506), .Y(n_601) );
AND2x2_ASAP7_75t_L g664 ( .A(n_506), .B(n_559), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_506), .A2(n_667), .B1(n_669), .B2(n_671), .C(n_672), .Y(n_666) );
AND2x2_ASAP7_75t_L g680 ( .A(n_506), .B(n_554), .Y(n_680) );
AND2x2_ASAP7_75t_L g706 ( .A(n_506), .B(n_590), .Y(n_706) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g586 ( .A(n_507), .B(n_559), .Y(n_586) );
BUFx2_ASAP7_75t_L g720 ( .A(n_507), .Y(n_720) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI32xp33_ASAP7_75t_L g686 ( .A1(n_518), .A2(n_647), .A3(n_661), .B1(n_687), .B2(n_688), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .Y(n_518) );
AND2x2_ASAP7_75t_L g627 ( .A(n_519), .B(n_571), .Y(n_627) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g609 ( .A(n_520), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_520), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g681 ( .A(n_520), .B(n_571), .Y(n_681) );
AND2x2_ASAP7_75t_L g692 ( .A(n_520), .B(n_584), .Y(n_692) );
BUFx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g593 ( .A(n_521), .B(n_572), .Y(n_593) );
AND2x2_ASAP7_75t_L g597 ( .A(n_521), .B(n_572), .Y(n_597) );
AND2x2_ASAP7_75t_L g632 ( .A(n_521), .B(n_583), .Y(n_632) );
AND2x2_ASAP7_75t_L g639 ( .A(n_521), .B(n_541), .Y(n_639) );
OAI211xp5_ASAP7_75t_L g644 ( .A1(n_521), .A2(n_590), .B(n_601), .C(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g698 ( .A(n_521), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_521), .B(n_532), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_530), .B(n_581), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_530), .B(n_597), .Y(n_687) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g592 ( .A(n_531), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_541), .Y(n_531) );
AND2x2_ASAP7_75t_L g584 ( .A(n_532), .B(n_542), .Y(n_584) );
OR2x2_ASAP7_75t_L g599 ( .A(n_532), .B(n_542), .Y(n_599) );
AND2x2_ASAP7_75t_L g622 ( .A(n_532), .B(n_583), .Y(n_622) );
INVx1_ASAP7_75t_L g626 ( .A(n_532), .Y(n_626) );
AND2x2_ASAP7_75t_L g645 ( .A(n_532), .B(n_582), .Y(n_645) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_532), .A2(n_610), .B1(n_656), .B2(n_657), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_532), .B(n_698), .Y(n_722) );
AND2x2_ASAP7_75t_L g737 ( .A(n_532), .B(n_597), .Y(n_737) );
INVx4_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx3_ASAP7_75t_L g569 ( .A(n_533), .Y(n_569) );
AND2x2_ASAP7_75t_L g611 ( .A(n_533), .B(n_542), .Y(n_611) );
AND2x2_ASAP7_75t_L g613 ( .A(n_533), .B(n_571), .Y(n_613) );
AND3x2_ASAP7_75t_L g675 ( .A(n_533), .B(n_639), .C(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g710 ( .A(n_541), .B(n_582), .Y(n_710) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g571 ( .A(n_542), .B(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_542), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_542), .B(n_581), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_542), .B(n_622), .C(n_698), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_568), .B1(n_580), .B2(n_585), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_554), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g662 ( .A(n_554), .Y(n_662) );
OAI31xp33_ASAP7_75t_L g678 ( .A1(n_557), .A2(n_679), .A3(n_680), .B(n_681), .Y(n_678) );
AND2x2_ASAP7_75t_L g703 ( .A(n_557), .B(n_590), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_557), .B(n_616), .Y(n_749) );
AND2x2_ASAP7_75t_L g658 ( .A(n_558), .B(n_590), .Y(n_658) );
AND2x2_ASAP7_75t_L g719 ( .A(n_558), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g589 ( .A(n_559), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g647 ( .A(n_559), .Y(n_647) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
CKINVDCx16_ASAP7_75t_R g668 ( .A(n_569), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_570), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AOI221x1_ASAP7_75t_SL g635 ( .A1(n_571), .A2(n_636), .B1(n_638), .B2(n_640), .C(n_642), .Y(n_635) );
INVx2_ASAP7_75t_L g583 ( .A(n_572), .Y(n_583) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_572), .Y(n_677) );
INVx1_ASAP7_75t_L g665 ( .A(n_580), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_581), .B(n_598), .Y(n_690) );
INVx1_ASAP7_75t_SL g753 ( .A(n_581), .Y(n_753) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g671 ( .A(n_584), .B(n_597), .Y(n_671) );
INVx1_ASAP7_75t_L g739 ( .A(n_585), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_585), .B(n_668), .Y(n_752) );
INVx2_ASAP7_75t_SL g591 ( .A(n_586), .Y(n_591) );
AND2x2_ASAP7_75t_L g634 ( .A(n_586), .B(n_590), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_586), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_586), .B(n_661), .Y(n_688) );
AOI21xp33_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_591), .B(n_592), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_589), .B(n_661), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_589), .B(n_616), .Y(n_757) );
OR2x2_ASAP7_75t_L g629 ( .A(n_590), .B(n_608), .Y(n_629) );
AND2x2_ASAP7_75t_L g728 ( .A(n_590), .B(n_719), .Y(n_728) );
OAI22xp5_ASAP7_75t_SL g603 ( .A1(n_591), .A2(n_604), .B1(n_609), .B2(n_612), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_591), .B(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g651 ( .A(n_593), .B(n_599), .Y(n_651) );
INVx1_ASAP7_75t_L g715 ( .A(n_593), .Y(n_715) );
AOI311xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_600), .A3(n_602), .B(n_603), .C(n_614), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_598), .A2(n_730), .B1(n_742), .B2(n_745), .C(n_747), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_598), .B(n_753), .Y(n_755) );
INVx2_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g652 ( .A(n_600), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g642 ( .A1(n_601), .A2(n_643), .B(n_644), .C(n_646), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_SL g711 ( .A1(n_605), .A2(n_607), .B(n_712), .C(n_713), .Y(n_711) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_606), .B(n_680), .Y(n_746) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
OAI221xp5_ASAP7_75t_L g628 ( .A1(n_609), .A2(n_629), .B1(n_630), .B2(n_633), .C(n_635), .Y(n_628) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g631 ( .A(n_611), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g714 ( .A(n_611), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_618), .Y(n_614) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_615), .A2(n_673), .B(n_674), .C(n_678), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_616), .B(n_617), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_616), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_616), .B(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVxp67_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g638 ( .A(n_622), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_626), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g740 ( .A(n_629), .Y(n_740) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_632), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g667 ( .A(n_632), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g744 ( .A(n_632), .Y(n_744) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g685 ( .A(n_634), .B(n_661), .Y(n_685) );
INVx1_ASAP7_75t_SL g679 ( .A(n_641), .Y(n_679) );
INVx1_ASAP7_75t_L g656 ( .A(n_647), .Y(n_656) );
NAND3xp33_ASAP7_75t_SL g648 ( .A(n_649), .B(n_666), .C(n_682), .Y(n_648) );
AOI322xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .A3(n_653), .B1(n_655), .B2(n_659), .C1(n_663), .C2(n_665), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g702 ( .A1(n_650), .A2(n_703), .B(n_704), .C(n_711), .Y(n_702) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_653), .A2(n_674), .B1(n_705), .B2(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g663 ( .A(n_661), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g700 ( .A(n_661), .B(n_701), .Y(n_700) );
AOI32xp33_ASAP7_75t_L g751 ( .A1(n_661), .A2(n_752), .A3(n_753), .B1(n_754), .B2(n_756), .Y(n_751) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g673 ( .A(n_664), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_664), .A2(n_717), .B1(n_721), .B2(n_723), .C(n_726), .Y(n_716) );
AND2x2_ASAP7_75t_L g730 ( .A(n_664), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g733 ( .A(n_668), .B(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g743 ( .A(n_668), .B(n_744), .Y(n_743) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g734 ( .A(n_677), .B(n_698), .Y(n_734) );
AOI211xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_685), .B(n_686), .C(n_689), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B(n_693), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI211xp5_ASAP7_75t_SL g695 ( .A1(n_696), .A2(n_699), .B(n_702), .C(n_716), .Y(n_695) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_710), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g725 ( .A(n_722), .Y(n_725) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI21xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_729), .B(n_732), .Y(n_726) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OAI211xp5_ASAP7_75t_SL g735 ( .A1(n_736), .A2(n_738), .B(n_741), .C(n_751), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI21xp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B(n_750), .Y(n_747) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx3_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
NAND2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
endmodule