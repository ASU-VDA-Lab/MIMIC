module fake_jpeg_1490_n_571 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_571);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_571;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_56),
.Y(n_157)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_58),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_28),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_62),
.Y(n_171)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_87),
.Y(n_121)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_78),
.B(n_98),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_51),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_92),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

BUFx2_ASAP7_75t_R g91 ( 
.A(n_43),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_91),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_20),
.B(n_18),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_39),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_100),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_20),
.B(n_15),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

BUFx8_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_43),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_19),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_106),
.B(n_23),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_44),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_109),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_44),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_111),
.B(n_54),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_40),
.B1(n_50),
.B2(n_46),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_115),
.A2(n_45),
.B1(n_35),
.B2(n_61),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_106),
.B(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_116),
.B(n_127),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_23),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_72),
.A2(n_49),
.B1(n_37),
.B2(n_36),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_130),
.A2(n_154),
.B1(n_24),
.B2(n_29),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_58),
.B(n_49),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_131),
.B(n_144),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_53),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_77),
.A2(n_36),
.B1(n_33),
.B2(n_19),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_146),
.A2(n_56),
.B1(n_40),
.B2(n_32),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_53),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_155),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_159),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_74),
.A2(n_33),
.B1(n_37),
.B2(n_45),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_68),
.B(n_50),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_75),
.B(n_32),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_156),
.B(n_174),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_89),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_94),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_177),
.Y(n_195)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_84),
.B(n_26),
.Y(n_170)
);

OR2x2_ASAP7_75t_SL g241 ( 
.A(n_170),
.B(n_1),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_59),
.B(n_46),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_82),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_120),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_178),
.B(n_216),
.Y(n_269)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_180),
.A2(n_186),
.B1(n_188),
.B2(n_224),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_182),
.A2(n_129),
.B1(n_122),
.B2(n_110),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_183),
.B(n_193),
.Y(n_278)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_185),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_124),
.A2(n_24),
.B1(n_29),
.B2(n_35),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_114),
.B(n_107),
.C(n_79),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_187),
.B(n_221),
.C(n_151),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_189),
.Y(n_290)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_190),
.Y(n_288)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_192),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_142),
.B(n_136),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_196),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_139),
.B(n_15),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_197),
.B(n_201),
.Y(n_298)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_198),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_171),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_199),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_200),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_121),
.B(n_69),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_125),
.B(n_83),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_203),
.B(n_231),
.Y(n_299)
);

CKINVDCx12_ASAP7_75t_R g204 ( 
.A(n_118),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_204),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_132),
.Y(n_205)
);

INVx11_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_123),
.Y(n_206)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_206),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_95),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_226),
.Y(n_252)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_208),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_153),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_209),
.B(n_214),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_210),
.Y(n_277)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_119),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_211),
.Y(n_255)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_213),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_137),
.B(n_15),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_215),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_168),
.A2(n_86),
.B1(n_85),
.B2(n_70),
.Y(n_216)
);

INVx4_ASAP7_75t_SL g217 ( 
.A(n_147),
.Y(n_217)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_219),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_126),
.B(n_71),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_220),
.B(n_230),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_170),
.B(n_140),
.C(n_113),
.Y(n_221)
);

AO22x2_ASAP7_75t_L g222 ( 
.A1(n_160),
.A2(n_76),
.B1(n_67),
.B2(n_104),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_222),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_145),
.A2(n_64),
.B1(n_55),
.B2(n_26),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_160),
.B(n_110),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_154),
.A2(n_22),
.B1(n_44),
.B2(n_2),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_118),
.B(n_0),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_112),
.B(n_22),
.CI(n_2),
.CON(n_227),
.SN(n_227)
);

AOI32xp33_ASAP7_75t_L g284 ( 
.A1(n_227),
.A2(n_148),
.A3(n_128),
.B1(n_7),
.B2(n_8),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_118),
.B(n_1),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_232),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_153),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_135),
.B(n_1),
.Y(n_231)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_135),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_233),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_112),
.Y(n_234)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_234),
.Y(n_287)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_141),
.Y(n_235)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_235),
.Y(n_297)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_143),
.Y(n_236)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_236),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_130),
.A2(n_54),
.B1(n_2),
.B2(n_3),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_173),
.B1(n_172),
.B2(n_122),
.Y(n_247)
);

OR2x4_ASAP7_75t_L g238 ( 
.A(n_146),
.B(n_1),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_241),
.B(n_2),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_239),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_143),
.B(n_150),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_216),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_243),
.B(n_257),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_176),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_244),
.A2(n_223),
.B(n_222),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_247),
.A2(n_251),
.B1(n_286),
.B2(n_294),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_224),
.A2(n_150),
.B1(n_173),
.B2(n_117),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_250),
.A2(n_239),
.B1(n_213),
.B2(n_185),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_117),
.B1(n_134),
.B2(n_129),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_145),
.C(n_151),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_254),
.B(n_275),
.C(n_5),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_265),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_243),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_147),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_273),
.B(n_279),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_148),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_183),
.B(n_147),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_238),
.A2(n_182),
.B1(n_222),
.B2(n_203),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_202),
.B(n_148),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_292),
.B(n_296),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_188),
.A2(n_134),
.B1(n_128),
.B2(n_133),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_295),
.A2(n_190),
.B1(n_208),
.B2(n_196),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_242),
.B(n_133),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_300),
.B(n_339),
.Y(n_371)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_302),
.Y(n_351)
);

AND2x6_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_241),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_310),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_293),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_305),
.B(n_309),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_181),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_308),
.Y(n_350)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_307),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_195),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_278),
.B(n_184),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_264),
.Y(n_310)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_285),
.Y(n_312)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_312),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_254),
.B(n_240),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_314),
.B(n_319),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_315),
.A2(n_289),
.B(n_264),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_267),
.A2(n_200),
.B(n_227),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_316),
.A2(n_317),
.B(n_290),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_257),
.A2(n_227),
.B(n_199),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_244),
.A2(n_205),
.B1(n_211),
.B2(n_218),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_318),
.A2(n_290),
.B1(n_256),
.B2(n_260),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_252),
.B(n_187),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_178),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_320),
.B(n_325),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_270),
.B(n_179),
.Y(n_321)
);

XNOR2x1_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_339),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_266),
.A2(n_191),
.B1(n_236),
.B2(n_235),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_322),
.A2(n_324),
.B1(n_330),
.B2(n_331),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_323),
.A2(n_326),
.B1(n_289),
.B2(n_253),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_263),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_294),
.A2(n_206),
.B1(n_194),
.B2(n_217),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_249),
.B(n_210),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_327),
.B(n_332),
.Y(n_363)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_256),
.Y(n_328)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_328),
.Y(n_362)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_246),
.Y(n_329)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_329),
.Y(n_364)
);

OAI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_244),
.A2(n_233),
.B1(n_189),
.B2(n_205),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_248),
.A2(n_198),
.B1(n_5),
.B2(n_7),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_258),
.B(n_3),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_333),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_265),
.B(n_3),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_334),
.B(n_335),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_3),
.Y(n_335)
);

BUFx4f_ASAP7_75t_SL g336 ( 
.A(n_274),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_336),
.Y(n_380)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_297),
.Y(n_337)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_338),
.Y(n_374)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_245),
.Y(n_340)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_340),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_287),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_341),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_280),
.B(n_7),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_343),
.B(n_345),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_255),
.B(n_244),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_262),
.B(n_8),
.C(n_10),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_277),
.C(n_272),
.Y(n_387)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_288),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_288),
.Y(n_366)
);

OA22x2_ASAP7_75t_L g348 ( 
.A1(n_269),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_348),
.B(n_269),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_313),
.A2(n_269),
.B1(n_250),
.B2(n_281),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_353),
.A2(n_375),
.B1(n_336),
.B2(n_307),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_300),
.B(n_268),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_354),
.B(n_383),
.C(n_385),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_355),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_313),
.A2(n_271),
.B1(n_259),
.B2(n_255),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_356),
.A2(n_377),
.B1(n_329),
.B2(n_302),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_358),
.A2(n_379),
.B(n_382),
.Y(n_410)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_301),
.B(n_342),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_370),
.B(n_381),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_371),
.B(n_304),
.Y(n_394)
);

BUFx4f_ASAP7_75t_SL g414 ( 
.A(n_376),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_313),
.A2(n_253),
.B1(n_245),
.B2(n_261),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_335),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_378),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_308),
.B(n_276),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_316),
.A2(n_317),
.B(n_345),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_314),
.B(n_261),
.Y(n_383)
);

AO22x1_ASAP7_75t_L g384 ( 
.A1(n_326),
.A2(n_260),
.B1(n_282),
.B2(n_276),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_338),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_321),
.B(n_282),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_387),
.B(n_12),
.Y(n_427)
);

NAND2xp33_ASAP7_75t_L g389 ( 
.A(n_306),
.B(n_277),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_389),
.B(n_349),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_319),
.B(n_272),
.C(n_11),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_390),
.B(n_334),
.C(n_346),
.Y(n_393)
);

BUFx12_ASAP7_75t_L g392 ( 
.A(n_380),
.Y(n_392)
);

BUFx12_ASAP7_75t_L g440 ( 
.A(n_392),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_393),
.B(n_400),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_394),
.B(n_427),
.Y(n_434)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_396),
.Y(n_447)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_351),
.Y(n_397)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_397),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_412),
.Y(n_432)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_399),
.B(n_403),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_360),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_353),
.A2(n_303),
.B1(n_311),
.B2(n_323),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_402),
.A2(n_404),
.B1(n_406),
.B2(n_411),
.Y(n_428)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_364),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_365),
.A2(n_311),
.B1(n_315),
.B2(n_310),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_340),
.C(n_337),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_405),
.B(n_415),
.C(n_385),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_365),
.A2(n_344),
.B1(n_333),
.B2(n_348),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_373),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_407),
.Y(n_436)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_408),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_348),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_409),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_379),
.A2(n_344),
.B1(n_348),
.B2(n_347),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_413),
.A2(n_422),
.B1(n_384),
.B2(n_375),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_354),
.B(n_312),
.C(n_336),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_374),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_416),
.B(n_419),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_382),
.A2(n_328),
.B(n_12),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_417),
.A2(n_424),
.B(n_367),
.Y(n_433)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_374),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_378),
.B(n_10),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_425),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_355),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_422)
);

INVx6_ASAP7_75t_L g423 ( 
.A(n_372),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_372),
.Y(n_456)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_352),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_377),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_426),
.B(n_363),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_420),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_429),
.B(n_430),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_423),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_433),
.B(n_441),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_410),
.A2(n_357),
.B(n_358),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_435),
.A2(n_439),
.B(n_443),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_437),
.B(n_444),
.Y(n_460)
);

A2O1A1O1Ixp25_ASAP7_75t_L g438 ( 
.A1(n_394),
.A2(n_350),
.B(n_355),
.C(n_386),
.D(n_361),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_438),
.A2(n_362),
.B(n_425),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_410),
.A2(n_417),
.B(n_409),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_412),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_401),
.B(n_350),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_442),
.B(n_457),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_418),
.A2(n_383),
.B(n_386),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_391),
.B(n_361),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_391),
.B(n_390),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_453),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_451),
.A2(n_459),
.B1(n_396),
.B2(n_408),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_452),
.A2(n_352),
.B1(n_384),
.B2(n_13),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_405),
.B(n_387),
.Y(n_453)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_456),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_398),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_415),
.B(n_388),
.C(n_369),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_369),
.C(n_359),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_404),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_418),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_469),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_432),
.A2(n_402),
.B1(n_411),
.B2(n_409),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_463),
.A2(n_466),
.B1(n_470),
.B2(n_486),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_432),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_464),
.B(n_478),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_435),
.A2(n_406),
.B(n_395),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_465),
.A2(n_481),
.B(n_450),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_432),
.A2(n_414),
.B1(n_421),
.B2(n_397),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_444),
.B(n_393),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_467),
.B(n_468),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_434),
.B(n_453),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_437),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_443),
.B(n_422),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_476),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_428),
.A2(n_368),
.B1(n_407),
.B2(n_414),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_475),
.A2(n_484),
.B1(n_452),
.B2(n_447),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_431),
.B(n_388),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_477),
.B(n_480),
.C(n_483),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_458),
.B(n_362),
.C(n_359),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_455),
.A2(n_414),
.B(n_392),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_438),
.B(n_352),
.C(n_392),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_445),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_485),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_455),
.A2(n_439),
.B1(n_428),
.B2(n_436),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_474),
.Y(n_488)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_488),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_489),
.A2(n_500),
.B1(n_508),
.B2(n_509),
.Y(n_515)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_466),
.Y(n_490)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_490),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_476),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_492),
.B(n_493),
.Y(n_524)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_479),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_482),
.A2(n_433),
.B(n_436),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_494),
.A2(n_496),
.B(n_440),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_461),
.B(n_449),
.Y(n_495)
);

MAJx2_ASAP7_75t_L g517 ( 
.A(n_495),
.B(n_505),
.C(n_462),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_482),
.A2(n_465),
.B(n_472),
.Y(n_496)
);

CKINVDCx14_ASAP7_75t_R g497 ( 
.A(n_483),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_497),
.B(n_499),
.Y(n_527)
);

AOI21x1_ASAP7_75t_L g519 ( 
.A1(n_498),
.A2(n_481),
.B(n_473),
.Y(n_519)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_471),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_463),
.A2(n_450),
.B1(n_449),
.B2(n_454),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_460),
.B(n_448),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_477),
.B(n_454),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_507),
.Y(n_511)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_486),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_475),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_462),
.C(n_480),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_510),
.B(n_523),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_505),
.B(n_469),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_513),
.B(n_516),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_468),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_520),
.Y(n_539)
);

BUFx12_ASAP7_75t_L g518 ( 
.A(n_492),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_518),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_519),
.A2(n_522),
.B(n_498),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_496),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_503),
.A2(n_460),
.B1(n_467),
.B2(n_440),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_521),
.A2(n_526),
.B1(n_494),
.B2(n_501),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_507),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_489),
.A2(n_440),
.B1(n_502),
.B2(n_509),
.Y(n_525)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_525),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_503),
.A2(n_490),
.B1(n_500),
.B2(n_508),
.Y(n_526)
);

AO21x1_ASAP7_75t_L g544 ( 
.A1(n_529),
.A2(n_541),
.B(n_542),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_SL g551 ( 
.A(n_530),
.B(n_518),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_512),
.B(n_495),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_532),
.B(n_533),
.Y(n_552)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_524),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_510),
.B(n_487),
.C(n_504),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_534),
.B(n_521),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_511),
.B(n_491),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_520),
.Y(n_543)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_524),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_540),
.Y(n_546)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_527),
.Y(n_540)
);

FAx1_ASAP7_75t_SL g541 ( 
.A(n_517),
.B(n_504),
.CI(n_491),
.CON(n_541),
.SN(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_522),
.A2(n_519),
.B(n_514),
.Y(n_542)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_543),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_538),
.B(n_531),
.C(n_513),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_545),
.B(n_547),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_531),
.B(n_516),
.C(n_511),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_548),
.A2(n_553),
.B(n_535),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_539),
.B(n_515),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_549),
.B(n_550),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_537),
.B(n_526),
.Y(n_550)
);

AND2x4_ASAP7_75t_SL g555 ( 
.A(n_551),
.B(n_544),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_528),
.B(n_530),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_554),
.B(n_555),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_546),
.A2(n_542),
.B1(n_529),
.B2(n_534),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_556),
.A2(n_539),
.B(n_551),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_558),
.A2(n_544),
.B(n_545),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_561),
.B(n_562),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_557),
.B(n_552),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_563),
.A2(n_555),
.B(n_559),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_565),
.B(n_560),
.C(n_518),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_566),
.B(n_564),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_567),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_568),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_541),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_541),
.Y(n_571)
);


endmodule