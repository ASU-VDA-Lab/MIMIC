module fake_aes_11149_n_42 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_42);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_40;
wire n_29;
wire n_39;
BUFx6f_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_8), .B(n_5), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_5), .Y(n_17) );
OAI22xp5_ASAP7_75t_L g18 ( .A1(n_13), .A2(n_8), .B1(n_1), .B2(n_7), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_2), .Y(n_19) );
NOR2x1_ASAP7_75t_L g20 ( .A(n_2), .B(n_6), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_3), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_11), .Y(n_22) );
BUFx2_ASAP7_75t_L g23 ( .A(n_17), .Y(n_23) );
NAND2xp33_ASAP7_75t_L g24 ( .A(n_15), .B(n_14), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
OAI21x1_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_21), .B(n_20), .Y(n_26) );
AO21x2_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_16), .B(n_18), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_26), .B(n_23), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_29), .B(n_23), .Y(n_30) );
INVx1_ASAP7_75t_SL g31 ( .A(n_28), .Y(n_31) );
OAI21xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_16), .B(n_27), .Y(n_32) );
AOI31xp33_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_27), .A3(n_1), .B(n_3), .Y(n_33) );
AOI221xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_27), .B1(n_22), .B2(n_15), .C(n_7), .Y(n_34) );
AOI22xp5_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_27), .B1(n_22), .B2(n_15), .Y(n_35) );
INVx1_ASAP7_75t_SL g36 ( .A(n_33), .Y(n_36) );
AND2x4_ASAP7_75t_L g37 ( .A(n_36), .B(n_0), .Y(n_37) );
AND3x4_ASAP7_75t_L g38 ( .A(n_34), .B(n_0), .C(n_4), .Y(n_38) );
NAND4xp75_ASAP7_75t_L g39 ( .A(n_35), .B(n_4), .C(n_6), .D(n_10), .Y(n_39) );
OR5x1_ASAP7_75t_L g40 ( .A(n_38), .B(n_12), .C(n_15), .D(n_22), .E(n_39), .Y(n_40) );
AO22x2_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_39), .B1(n_36), .B2(n_37), .Y(n_41) );
INVxp67_ASAP7_75t_L g42 ( .A(n_41), .Y(n_42) );
endmodule