module fake_netlist_6_4042_n_1889 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_442, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_443, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_446, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_433, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1889);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_433;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1889;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_1380;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1697;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_527;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_1466;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1737;
wire n_653;
wire n_1464;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_1028;
wire n_576;
wire n_472;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_1884;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_183),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_58),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_69),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_157),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_229),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_453),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_184),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_327),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_28),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_421),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_446),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_149),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_47),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_449),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_105),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_217),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_271),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_21),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_355),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_118),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_323),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_126),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_280),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_255),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_435),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_416),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_342),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_432),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_411),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_90),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_335),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_148),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_436),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_192),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_427),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_309),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_334),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_237),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_286),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_373),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_251),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_431),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_20),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_167),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_112),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_442),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_417),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_410),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_290),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_194),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_73),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_80),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_302),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_24),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_89),
.Y(n_512)
);

BUFx5_ASAP7_75t_L g513 ( 
.A(n_447),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_171),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_31),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_450),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_208),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_250),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_353),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_196),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_234),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_399),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_438),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_295),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_380),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_67),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_347),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_404),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_406),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_333),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_388),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_213),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_389),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_424),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_65),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_273),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_233),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_372),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_164),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_216),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_0),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_265),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_354),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_443),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_289),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_366),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_9),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_48),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_159),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_391),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_420),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_74),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_266),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_387),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_173),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_254),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_209),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_149),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_34),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_132),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_418),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_219),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_257),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_94),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_433),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_47),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_419),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_145),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_276),
.Y(n_569)
);

BUFx8_ASAP7_75t_SL g570 ( 
.A(n_319),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_210),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_171),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_303),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_195),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_113),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_297),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_197),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_2),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_296),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_35),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_202),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_390),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_392),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_359),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_440),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_434),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_350),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_321),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_457),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_215),
.Y(n_590)
);

BUFx5_ASAP7_75t_L g591 ( 
.A(n_95),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_156),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_454),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_123),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_134),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_31),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_345),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_249),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_246),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_17),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_18),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_364),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_80),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_49),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_61),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_337),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_344),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_159),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_20),
.Y(n_609)
);

BUFx8_ASAP7_75t_SL g610 ( 
.A(n_451),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_63),
.Y(n_611)
);

CKINVDCx16_ASAP7_75t_R g612 ( 
.A(n_437),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_384),
.Y(n_613)
);

CKINVDCx16_ASAP7_75t_R g614 ( 
.A(n_352),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_444),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_408),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_14),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_403),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_423),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_17),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_363),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_262),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_98),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_112),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_76),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_18),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_50),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_107),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_365),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_117),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_142),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_62),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_287),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_185),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_107),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_85),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_267),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_151),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_439),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_79),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_119),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_193),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_129),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_152),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_174),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_178),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_430),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_325),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_139),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_236),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_244),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_212),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_258),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_122),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_429),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_320),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_304),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_283),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_422),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_121),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_76),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_409),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_182),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_338),
.Y(n_664)
);

CKINVDCx16_ASAP7_75t_R g665 ( 
.A(n_328),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_269),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_214),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_147),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_15),
.Y(n_669)
);

CKINVDCx14_ASAP7_75t_R g670 ( 
.A(n_13),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_113),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_351),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_324),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_239),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_322),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_376),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_82),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_378),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_102),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_348),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_43),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_426),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_188),
.Y(n_683)
);

BUFx10_ASAP7_75t_L g684 ( 
.A(n_428),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_332),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_441),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_425),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_591),
.Y(n_688)
);

INVxp67_ASAP7_75t_SL g689 ( 
.A(n_683),
.Y(n_689)
);

INVxp33_ASAP7_75t_L g690 ( 
.A(n_654),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_570),
.Y(n_691)
);

CKINVDCx16_ASAP7_75t_R g692 ( 
.A(n_612),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_654),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_512),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_591),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_610),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_500),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_566),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_617),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_591),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_591),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_458),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_462),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_591),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_603),
.Y(n_705)
);

INVxp33_ASAP7_75t_L g706 ( 
.A(n_459),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_603),
.Y(n_707)
);

INVxp33_ASAP7_75t_SL g708 ( 
.A(n_683),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_625),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_625),
.Y(n_710)
);

INVxp33_ASAP7_75t_L g711 ( 
.A(n_479),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_463),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_514),
.Y(n_713)
);

INVxp33_ASAP7_75t_SL g714 ( 
.A(n_460),
.Y(n_714)
);

INVxp33_ASAP7_75t_L g715 ( 
.A(n_515),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_467),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_631),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_513),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_513),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_564),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_568),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_572),
.Y(n_722)
);

CKINVDCx16_ASAP7_75t_R g723 ( 
.A(n_614),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_681),
.Y(n_724)
);

INVxp67_ASAP7_75t_SL g725 ( 
.A(n_471),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_601),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_596),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_468),
.Y(n_728)
);

INVxp33_ASAP7_75t_SL g729 ( 
.A(n_461),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_608),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_624),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_474),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_494),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_476),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_480),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_637),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_627),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_504),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_643),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_644),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_668),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_671),
.Y(n_742)
);

CKINVDCx16_ASAP7_75t_R g743 ( 
.A(n_665),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_478),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_478),
.Y(n_745)
);

INVxp67_ASAP7_75t_SL g746 ( 
.A(n_529),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_529),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_544),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_544),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_581),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_581),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_482),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_588),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_588),
.Y(n_754)
);

INVxp67_ASAP7_75t_SL g755 ( 
.A(n_589),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_483),
.Y(n_756)
);

INVxp33_ASAP7_75t_L g757 ( 
.A(n_535),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_589),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_655),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_513),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_655),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_663),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_670),
.Y(n_763)
);

INVxp67_ASAP7_75t_SL g764 ( 
.A(n_663),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_678),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_484),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_466),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_678),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_465),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_672),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_763),
.B(n_491),
.Y(n_771)
);

BUFx12f_ASAP7_75t_L g772 ( 
.A(n_691),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_738),
.Y(n_773)
);

OA21x2_ASAP7_75t_L g774 ( 
.A1(n_688),
.A2(n_481),
.B(n_473),
.Y(n_774)
);

OA21x2_ASAP7_75t_L g775 ( 
.A1(n_695),
.A2(n_488),
.B(n_485),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_709),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_738),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_710),
.Y(n_778)
);

INVx6_ASAP7_75t_L g779 ( 
.A(n_738),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_769),
.B(n_744),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_745),
.B(n_590),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_747),
.B(n_556),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_700),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_770),
.Y(n_784)
);

XOR2xp5_ASAP7_75t_L g785 ( 
.A(n_694),
.B(n_464),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_708),
.B(n_670),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_690),
.A2(n_604),
.B1(n_469),
.B2(n_472),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_767),
.Y(n_788)
);

AOI22x1_ASAP7_75t_SL g789 ( 
.A1(n_694),
.A2(n_470),
.B1(n_477),
.B2(n_475),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_748),
.B(n_556),
.Y(n_790)
);

INVxp33_ASAP7_75t_SL g791 ( 
.A(n_702),
.Y(n_791)
);

INVx6_ASAP7_75t_L g792 ( 
.A(n_770),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_701),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_704),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_699),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_SL g796 ( 
.A1(n_699),
.A2(n_487),
.B1(n_501),
.B2(n_489),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_749),
.B(n_486),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_713),
.Y(n_798)
);

AOI22x1_ASAP7_75t_SL g799 ( 
.A1(n_717),
.A2(n_502),
.B1(n_509),
.B2(n_508),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_720),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_746),
.B(n_525),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_703),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_721),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_712),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_755),
.B(n_528),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_692),
.A2(n_496),
.B1(n_530),
.B2(n_521),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_716),
.Y(n_807)
);

INVx6_ASAP7_75t_L g808 ( 
.A(n_723),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_743),
.A2(n_629),
.B1(n_658),
.B2(n_573),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_722),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_726),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_730),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_731),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_737),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_739),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_740),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_741),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_742),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_718),
.Y(n_819)
);

INVx5_ASAP7_75t_L g820 ( 
.A(n_719),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_719),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_728),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_760),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_732),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_804),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_804),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_803),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_795),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_822),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_R g830 ( 
.A(n_822),
.B(n_696),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_810),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_791),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_791),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_777),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_786),
.B(n_734),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_772),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_811),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_R g838 ( 
.A(n_795),
.B(n_735),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_777),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_807),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_824),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_786),
.Y(n_842)
);

BUFx10_ASAP7_75t_L g843 ( 
.A(n_808),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_813),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_808),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_802),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_792),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_785),
.Y(n_848)
);

BUFx10_ASAP7_75t_L g849 ( 
.A(n_808),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_771),
.Y(n_850)
);

XNOR2xp5_ASAP7_75t_SL g851 ( 
.A(n_796),
.B(n_690),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_788),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_802),
.B(n_752),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_773),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_784),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_806),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_792),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_815),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_773),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_819),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_792),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_809),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_817),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_R g864 ( 
.A(n_797),
.B(n_756),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_773),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_789),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_799),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_788),
.Y(n_868)
);

INVxp67_ASAP7_75t_SL g869 ( 
.A(n_780),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_771),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_797),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_787),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_783),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_787),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_773),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_801),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_801),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_805),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_793),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_805),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_812),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_819),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_779),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_779),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_812),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_800),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_819),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_R g888 ( 
.A(n_814),
.B(n_766),
.Y(n_888)
);

BUFx10_ASAP7_75t_L g889 ( 
.A(n_800),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_800),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_800),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_816),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_816),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_814),
.B(n_725),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_816),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_781),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_781),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_794),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_816),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_780),
.Y(n_900)
);

NAND2xp33_ASAP7_75t_R g901 ( 
.A(n_774),
.B(n_714),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_823),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_779),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_871),
.B(n_714),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_852),
.Y(n_905)
);

BUFx10_ASAP7_75t_L g906 ( 
.A(n_853),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_852),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_868),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_842),
.B(n_729),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_869),
.B(n_823),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_842),
.B(n_729),
.Y(n_911)
);

AND2x2_ASAP7_75t_SL g912 ( 
.A(n_835),
.B(n_851),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_881),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_828),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_873),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_879),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_831),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_900),
.B(n_733),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_894),
.B(n_736),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_870),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_876),
.B(n_877),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_878),
.B(n_689),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_837),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_844),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_847),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_886),
.B(n_821),
.Y(n_926)
);

INVx6_ASAP7_75t_L g927 ( 
.A(n_843),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_858),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_863),
.Y(n_929)
);

AOI22x1_ASAP7_75t_L g930 ( 
.A1(n_872),
.A2(n_765),
.B1(n_764),
.B2(n_751),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_880),
.Y(n_931)
);

AND2x2_ASAP7_75t_SL g932 ( 
.A(n_874),
.B(n_620),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_830),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_885),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_896),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_834),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_855),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_839),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_887),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_843),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_890),
.B(n_774),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_891),
.B(n_775),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_850),
.B(n_698),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_846),
.B(n_697),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_849),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_883),
.B(n_798),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_849),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_892),
.B(n_775),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_883),
.B(n_884),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_857),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_884),
.Y(n_951)
);

AND2x6_ASAP7_75t_L g952 ( 
.A(n_860),
.B(n_504),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_903),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_SL g954 ( 
.A(n_864),
.B(n_685),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_893),
.B(n_686),
.Y(n_955)
);

BUFx6f_ASAP7_75t_SL g956 ( 
.A(n_845),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_840),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_SL g958 ( 
.A(n_832),
.B(n_717),
.Y(n_958)
);

BUFx10_ASAP7_75t_L g959 ( 
.A(n_825),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_826),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_862),
.B(n_727),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_887),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_895),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_889),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_899),
.B(n_492),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_882),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_897),
.A2(n_532),
.B1(n_538),
.B2(n_531),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_902),
.Y(n_968)
);

BUFx6f_ASAP7_75t_SL g969 ( 
.A(n_836),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_861),
.B(n_757),
.Y(n_970)
);

AO22x2_ASAP7_75t_L g971 ( 
.A1(n_856),
.A2(n_693),
.B1(n_636),
.B2(n_641),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_859),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_859),
.B(n_818),
.Y(n_973)
);

BUFx4f_ASAP7_75t_L g974 ( 
.A(n_865),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_865),
.B(n_705),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_841),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_902),
.Y(n_977)
);

OAI22xp33_ASAP7_75t_L g978 ( 
.A1(n_901),
.A2(n_790),
.B1(n_782),
.B2(n_711),
.Y(n_978)
);

BUFx8_ASAP7_75t_SL g979 ( 
.A(n_848),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_829),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_888),
.B(n_571),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_902),
.B(n_782),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_838),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_833),
.B(n_750),
.Y(n_984)
);

AND2x6_ASAP7_75t_L g985 ( 
.A(n_854),
.B(n_504),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_875),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_866),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_875),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_867),
.Y(n_989)
);

INVx8_ASAP7_75t_L g990 ( 
.A(n_857),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_873),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_898),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_842),
.B(n_724),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_843),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_842),
.B(n_724),
.Y(n_995)
);

AND2x6_ASAP7_75t_L g996 ( 
.A(n_894),
.B(n_504),
.Y(n_996)
);

AO22x2_ASAP7_75t_L g997 ( 
.A1(n_842),
.A2(n_660),
.B1(n_541),
.B2(n_661),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_827),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_827),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_827),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_847),
.B(n_707),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_869),
.B(n_790),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_881),
.Y(n_1003)
);

OR2x6_ASAP7_75t_L g1004 ( 
.A(n_845),
.B(n_753),
.Y(n_1004)
);

CKINVDCx16_ASAP7_75t_R g1005 ( 
.A(n_838),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_827),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_827),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_827),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_827),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_830),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_881),
.Y(n_1011)
);

AND2x6_ASAP7_75t_L g1012 ( 
.A(n_894),
.B(n_527),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_847),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_868),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_843),
.Y(n_1015)
);

AND2x2_ASAP7_75t_SL g1016 ( 
.A(n_835),
.B(n_495),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_850),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_900),
.B(n_757),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_923),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_972),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_970),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_1016),
.A2(n_499),
.B1(n_510),
.B2(n_497),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1002),
.B(n_516),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_905),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_932),
.A2(n_518),
.B1(n_522),
.B2(n_519),
.Y(n_1025)
);

OAI22xp33_ASAP7_75t_SL g1026 ( 
.A1(n_930),
.A2(n_758),
.B1(n_759),
.B2(n_754),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_979),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_919),
.B(n_542),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_960),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_980),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_916),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_916),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_905),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_907),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_924),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_978),
.B(n_545),
.Y(n_1036)
);

AND2x6_ASAP7_75t_L g1037 ( 
.A(n_941),
.B(n_546),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_1013),
.B(n_761),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_917),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_1018),
.Y(n_1040)
);

NAND2x1p5_ASAP7_75t_L g1041 ( 
.A(n_964),
.B(n_776),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_991),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_945),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_928),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_982),
.B(n_550),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_925),
.B(n_1001),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_922),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_1001),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_918),
.B(n_551),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_909),
.B(n_706),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_963),
.B(n_762),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_926),
.B(n_553),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_929),
.Y(n_1053)
);

AO22x2_ASAP7_75t_L g1054 ( 
.A1(n_967),
.A2(n_563),
.B1(n_565),
.B2(n_554),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_998),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_964),
.B(n_768),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_999),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1000),
.Y(n_1058)
);

AO22x2_ASAP7_75t_L g1059 ( 
.A1(n_961),
.A2(n_587),
.B1(n_593),
.B2(n_574),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1006),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1007),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1008),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1009),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_942),
.A2(n_674),
.B1(n_645),
.B2(n_599),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_975),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_975),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_SL g1067 ( 
.A1(n_912),
.A2(n_511),
.B1(n_594),
.B2(n_558),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_992),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_911),
.B(n_598),
.Y(n_1069)
);

AO22x2_ASAP7_75t_L g1070 ( 
.A1(n_904),
.A2(n_602),
.B1(n_616),
.B2(n_615),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_945),
.B(n_778),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_935),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_973),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_973),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_949),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_938),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_948),
.A2(n_622),
.B1(n_633),
.B2(n_619),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_954),
.A2(n_653),
.B1(n_657),
.B2(n_650),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_947),
.B(n_666),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_993),
.B(n_706),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_994),
.B(n_673),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_936),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_966),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_994),
.B(n_682),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_943),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_939),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_962),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_935),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_944),
.B(n_711),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_995),
.B(n_715),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_L g1091 ( 
.A(n_930),
.B(n_984),
.C(n_965),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_986),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_988),
.Y(n_1093)
);

CKINVDCx14_ASAP7_75t_R g1094 ( 
.A(n_914),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_946),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_908),
.B(n_715),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_1015),
.Y(n_1097)
);

INVxp67_ASAP7_75t_L g1098 ( 
.A(n_921),
.Y(n_1098)
);

AO22x2_ASAP7_75t_L g1099 ( 
.A1(n_1014),
.A2(n_596),
.B1(n_2),
.B2(n_0),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_968),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_949),
.B(n_175),
.Y(n_1101)
);

AO22x2_ASAP7_75t_L g1102 ( 
.A1(n_955),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_934),
.B(n_526),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_1003),
.B(n_176),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_977),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_1004),
.Y(n_1106)
);

AO22x2_ASAP7_75t_L g1107 ( 
.A1(n_971),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_951),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_920),
.A2(n_493),
.B1(n_498),
.B2(n_490),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_953),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_931),
.A2(n_505),
.B1(n_506),
.B2(n_503),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_996),
.B(n_507),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_1004),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_906),
.B(n_539),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1011),
.B(n_177),
.Y(n_1115)
);

INVxp67_ASAP7_75t_L g1116 ( 
.A(n_937),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_974),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_997),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_1005),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_997),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_927),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1012),
.A2(n_513),
.B1(n_540),
.B2(n_527),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1012),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_933),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1012),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_981),
.B(n_906),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_985),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_985),
.Y(n_1128)
);

AOI211xp5_ASAP7_75t_L g1129 ( 
.A1(n_958),
.A2(n_548),
.B(n_549),
.C(n_547),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_985),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1017),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_952),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_927),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_952),
.Y(n_1134)
);

NAND2x1p5_ASAP7_75t_L g1135 ( 
.A(n_940),
.B(n_527),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_957),
.B(n_552),
.Y(n_1136)
);

NAND2x1p5_ASAP7_75t_L g1137 ( 
.A(n_950),
.B(n_976),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_952),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_983),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_971),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_990),
.B(n_527),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_956),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_990),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_983),
.B(n_1010),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_959),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_959),
.Y(n_1146)
);

CKINVDCx16_ASAP7_75t_R g1147 ( 
.A(n_969),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_989),
.Y(n_1148)
);

INVxp67_ASAP7_75t_SL g1149 ( 
.A(n_989),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_987),
.B(n_559),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_915),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1016),
.A2(n_517),
.B(n_523),
.C(n_520),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_923),
.Y(n_1153)
);

AO22x2_ASAP7_75t_L g1154 ( 
.A1(n_967),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_913),
.B(n_524),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_923),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_909),
.B(n_560),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_915),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_979),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_915),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_964),
.B(n_540),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_905),
.Y(n_1162)
);

OA22x2_ASAP7_75t_L g1163 ( 
.A1(n_1018),
.A2(n_578),
.B1(n_580),
.B2(n_575),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_970),
.Y(n_1164)
);

OR2x6_ASAP7_75t_L g1165 ( 
.A(n_990),
.B(n_540),
.Y(n_1165)
);

NOR2x1p5_ASAP7_75t_L g1166 ( 
.A(n_940),
.B(n_592),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_970),
.Y(n_1167)
);

INVxp67_ASAP7_75t_SL g1168 ( 
.A(n_910),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_915),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1016),
.A2(n_533),
.B(n_536),
.C(n_534),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_923),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1157),
.A2(n_537),
.B(n_555),
.C(n_543),
.Y(n_1172)
);

AO22x1_ASAP7_75t_L g1173 ( 
.A1(n_1050),
.A2(n_600),
.B1(n_605),
.B2(n_595),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1168),
.A2(n_820),
.B(n_585),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1080),
.B(n_557),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1023),
.A2(n_820),
.B(n_647),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1090),
.B(n_609),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1097),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1047),
.B(n_611),
.Y(n_1179)
);

NAND2xp33_ASAP7_75t_L g1180 ( 
.A(n_1097),
.B(n_1121),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1045),
.A2(n_647),
.B(n_585),
.Y(n_1181)
);

NAND3xp33_ASAP7_75t_L g1182 ( 
.A(n_1025),
.B(n_626),
.C(n_623),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1164),
.B(n_672),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1089),
.B(n_561),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1031),
.B(n_562),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1077),
.A2(n_569),
.B(n_567),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1028),
.A2(n_659),
.B(n_577),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1052),
.A2(n_659),
.B(n_579),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1032),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_1097),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1069),
.A2(n_684),
.B(n_630),
.C(n_632),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1037),
.A2(n_582),
.B(n_576),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1039),
.A2(n_584),
.B1(n_586),
.B2(n_583),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1042),
.B(n_597),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1121),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1096),
.B(n_684),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1091),
.A2(n_607),
.B(n_613),
.C(n_606),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1040),
.B(n_628),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1037),
.A2(n_621),
.B(n_618),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1151),
.B(n_634),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1085),
.B(n_639),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1158),
.B(n_642),
.Y(n_1202)
);

AO21x1_ASAP7_75t_L g1203 ( 
.A1(n_1036),
.A2(n_5),
.B(n_6),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1160),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1021),
.B(n_635),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1169),
.A2(n_687),
.B(n_648),
.C(n_651),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1126),
.B(n_1167),
.Y(n_1207)
);

INVxp67_ASAP7_75t_L g1208 ( 
.A(n_1024),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1019),
.A2(n_652),
.B(n_646),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1044),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1053),
.Y(n_1211)
);

AO22x1_ASAP7_75t_L g1212 ( 
.A1(n_1149),
.A2(n_640),
.B1(n_649),
.B2(n_638),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1022),
.A2(n_680),
.B(n_662),
.C(n_664),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1049),
.B(n_656),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1062),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1153),
.A2(n_675),
.B(n_667),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1063),
.B(n_676),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1035),
.B(n_669),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1150),
.B(n_677),
.Y(n_1219)
);

O2A1O1Ixp5_ASAP7_75t_L g1220 ( 
.A1(n_1152),
.A2(n_180),
.B(n_181),
.C(n_179),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1055),
.A2(n_679),
.B1(n_187),
.B2(n_189),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1033),
.B(n_7),
.Y(n_1222)
);

INVx3_ASAP7_75t_SL g1223 ( 
.A(n_1029),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_SL g1224 ( 
.A(n_1030),
.B(n_1146),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1057),
.B(n_8),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1058),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1098),
.B(n_1162),
.Y(n_1227)
);

OAI321xp33_ASAP7_75t_L g1228 ( 
.A1(n_1067),
.A2(n_10),
.A3(n_12),
.B1(n_8),
.B2(n_9),
.C(n_11),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1034),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1060),
.B(n_1061),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1037),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1136),
.A2(n_190),
.B1(n_191),
.B2(n_186),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1156),
.B(n_13),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1088),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1046),
.B(n_1075),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1171),
.B(n_14),
.Y(n_1236)
);

NOR2x1p5_ASAP7_75t_SL g1237 ( 
.A(n_1123),
.B(n_1125),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1020),
.A2(n_199),
.B1(n_200),
.B2(n_198),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1139),
.B(n_15),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1037),
.B(n_1068),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1075),
.A2(n_203),
.B1(n_204),
.B2(n_201),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1078),
.A2(n_21),
.B(n_16),
.C(n_19),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1101),
.A2(n_206),
.B(n_205),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1082),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1104),
.B(n_207),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1064),
.A2(n_1170),
.B(n_1083),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1076),
.B(n_22),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1114),
.B(n_22),
.Y(n_1248)
);

BUFx2_ASAP7_75t_SL g1249 ( 
.A(n_1133),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1026),
.A2(n_1118),
.B(n_1120),
.C(n_1129),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1038),
.B(n_23),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1073),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1104),
.B(n_1115),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1038),
.B(n_23),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1048),
.A2(n_218),
.B(n_211),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1124),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1086),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1065),
.A2(n_1066),
.B1(n_1051),
.B2(n_1074),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1095),
.A2(n_221),
.B(n_220),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1115),
.B(n_222),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1103),
.B(n_25),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1051),
.B(n_223),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1027),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1121),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1070),
.B(n_25),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1108),
.A2(n_225),
.B1(n_226),
.B2(n_224),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1116),
.B(n_26),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1070),
.B(n_26),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1110),
.A2(n_228),
.B1(n_230),
.B2(n_227),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1144),
.B(n_27),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1092),
.B(n_27),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1046),
.B(n_231),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1140),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1112),
.A2(n_235),
.B(n_232),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1093),
.A2(n_240),
.B1(n_241),
.B2(n_238),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1072),
.B(n_29),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1087),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1117),
.A2(n_33),
.B(n_30),
.C(n_32),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1100),
.B(n_32),
.Y(n_1279)
);

O2A1O1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1111),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_1280)
);

INVxp67_ASAP7_75t_L g1281 ( 
.A(n_1106),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1155),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1056),
.A2(n_243),
.B1(n_245),
.B2(n_242),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1105),
.A2(n_248),
.B(n_247),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1127),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1122),
.A2(n_253),
.B(n_252),
.Y(n_1286)
);

OAI321xp33_ASAP7_75t_L g1287 ( 
.A1(n_1154),
.A2(n_36),
.A3(n_37),
.B1(n_38),
.B2(n_39),
.C(n_40),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_SL g1288 ( 
.A(n_1159),
.B(n_256),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1109),
.B(n_39),
.Y(n_1289)
);

AND2x6_ASAP7_75t_L g1290 ( 
.A(n_1128),
.B(n_259),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1130),
.A2(n_261),
.B(n_260),
.Y(n_1291)
);

NOR2xp67_ASAP7_75t_L g1292 ( 
.A(n_1148),
.B(n_263),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1113),
.B(n_40),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1132),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1079),
.A2(n_1084),
.B(n_1081),
.C(n_1131),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1054),
.B(n_41),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1079),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1134),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1102),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1043),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1054),
.B(n_44),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1138),
.A2(n_268),
.B(n_264),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1081),
.B(n_44),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1084),
.B(n_1059),
.Y(n_1304)
);

OAI321xp33_ASAP7_75t_L g1305 ( 
.A1(n_1154),
.A2(n_45),
.A3(n_46),
.B1(n_48),
.B2(n_49),
.C(n_50),
.Y(n_1305)
);

INVx3_ASAP7_75t_SL g1306 ( 
.A(n_1147),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1059),
.B(n_45),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1141),
.A2(n_272),
.B(n_270),
.Y(n_1308)
);

NOR2xp67_ASAP7_75t_L g1309 ( 
.A(n_1145),
.B(n_274),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1102),
.B(n_46),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1137),
.B(n_51),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1143),
.B(n_51),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1094),
.B(n_52),
.Y(n_1313)
);

BUFx8_ASAP7_75t_SL g1314 ( 
.A(n_1119),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1141),
.A2(n_277),
.B(n_275),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1165),
.A2(n_279),
.B(n_278),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1165),
.A2(n_1041),
.B(n_1161),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1166),
.B(n_281),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1071),
.B(n_52),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1142),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1135),
.A2(n_284),
.B(n_282),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1163),
.B(n_53),
.Y(n_1322)
);

NOR2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1107),
.B(n_285),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1107),
.A2(n_291),
.B(n_288),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1099),
.B(n_54),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1099),
.B(n_55),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1050),
.B(n_56),
.Y(n_1327)
);

O2A1O1Ixp5_ASAP7_75t_L g1328 ( 
.A1(n_1069),
.A2(n_293),
.B(n_294),
.C(n_292),
.Y(n_1328)
);

AO21x1_ASAP7_75t_L g1329 ( 
.A1(n_1036),
.A2(n_56),
.B(n_57),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1248),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1330)
);

AOI221xp5_ASAP7_75t_L g1331 ( 
.A1(n_1177),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.C(n_62),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1210),
.Y(n_1332)
);

OAI22x1_ASAP7_75t_L g1333 ( 
.A1(n_1323),
.A2(n_64),
.B1(n_60),
.B2(n_63),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1208),
.B(n_64),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1246),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1175),
.B(n_66),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1235),
.B(n_298),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1264),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1229),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_R g1340 ( 
.A(n_1256),
.B(n_299),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1211),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1264),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1195),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1327),
.B(n_68),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1197),
.A2(n_301),
.B(n_300),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1253),
.B(n_68),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1314),
.Y(n_1347)
);

O2A1O1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1270),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1215),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1234),
.B(n_70),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1224),
.B(n_1227),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1214),
.B(n_71),
.Y(n_1352)
);

CKINVDCx6p67_ASAP7_75t_R g1353 ( 
.A(n_1223),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1184),
.B(n_72),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1313),
.A2(n_78),
.B1(n_75),
.B2(n_77),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1289),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1189),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1207),
.B(n_81),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1295),
.B(n_81),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1178),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1258),
.B(n_82),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1300),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1219),
.B(n_83),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1280),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1230),
.B(n_84),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1304),
.B(n_86),
.Y(n_1366)
);

O2A1O1Ixp5_ASAP7_75t_L g1367 ( 
.A1(n_1186),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1204),
.B(n_87),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1250),
.A2(n_1286),
.B(n_1191),
.C(n_1261),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1205),
.B(n_88),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1178),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_SL g1372 ( 
.A1(n_1291),
.A2(n_306),
.B(n_307),
.C(n_305),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1226),
.B(n_89),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_R g1374 ( 
.A(n_1263),
.B(n_308),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1179),
.B(n_90),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_SL g1376 ( 
.A1(n_1284),
.A2(n_311),
.B(n_312),
.C(n_310),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1252),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1244),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1185),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1235),
.B(n_91),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1178),
.B(n_93),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1306),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1257),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1217),
.B(n_94),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1190),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1218),
.B(n_95),
.Y(n_1386)
);

CKINVDCx8_ASAP7_75t_R g1387 ( 
.A(n_1249),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1245),
.A2(n_314),
.B(n_313),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1281),
.Y(n_1389)
);

NOR3xp33_ASAP7_75t_SL g1390 ( 
.A(n_1228),
.B(n_96),
.C(n_97),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1196),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1318),
.B(n_1277),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_SL g1393 ( 
.A1(n_1260),
.A2(n_316),
.B(n_317),
.C(n_315),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1318),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1310),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_1395)
);

OR2x6_ASAP7_75t_L g1396 ( 
.A(n_1317),
.B(n_318),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1277),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1198),
.B(n_102),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1311),
.B(n_103),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_L g1400 ( 
.A(n_1173),
.B(n_1282),
.C(n_1242),
.Y(n_1400)
);

AO32x1_ASAP7_75t_L g1401 ( 
.A1(n_1299),
.A2(n_103),
.A3(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1194),
.A2(n_104),
.B1(n_106),
.B2(n_108),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1285),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1200),
.B(n_108),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1243),
.A2(n_329),
.B(n_326),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1174),
.A2(n_331),
.B(n_330),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1183),
.B(n_109),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1262),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1293),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1294),
.Y(n_1410)
);

NAND3xp33_ASAP7_75t_SL g1411 ( 
.A(n_1324),
.B(n_110),
.C(n_111),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1201),
.B(n_114),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1320),
.A2(n_1307),
.B(n_1268),
.C(n_1265),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1202),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1298),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1325),
.A2(n_115),
.B(n_116),
.C(n_117),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1276),
.B(n_118),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1290),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1240),
.A2(n_339),
.B(n_336),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1290),
.Y(n_1420)
);

BUFx2_ASAP7_75t_SL g1421 ( 
.A(n_1309),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1206),
.A2(n_341),
.B(n_340),
.Y(n_1422)
);

BUFx2_ASAP7_75t_R g1423 ( 
.A(n_1272),
.Y(n_1423)
);

O2A1O1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1326),
.A2(n_119),
.B(n_120),
.C(n_121),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1233),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1247),
.B(n_1225),
.Y(n_1426)
);

NAND2x1p5_ASAP7_75t_L g1427 ( 
.A(n_1312),
.B(n_343),
.Y(n_1427)
);

AND3x1_ASAP7_75t_SL g1428 ( 
.A(n_1287),
.B(n_120),
.C(n_122),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1303),
.B(n_123),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1271),
.B(n_124),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1222),
.Y(n_1431)
);

INVx3_ASAP7_75t_SL g1432 ( 
.A(n_1290),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1251),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1220),
.A2(n_125),
.B(n_127),
.C(n_128),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1290),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1236),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_SL g1437 ( 
.A(n_1203),
.B(n_127),
.C(n_128),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1279),
.Y(n_1438)
);

NOR3xp33_ASAP7_75t_L g1439 ( 
.A(n_1182),
.B(n_1322),
.C(n_1212),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1254),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1172),
.A2(n_129),
.B(n_130),
.C(n_131),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1319),
.B(n_130),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1180),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1296),
.Y(n_1444)
);

AO21x1_ASAP7_75t_L g1445 ( 
.A1(n_1274),
.A2(n_131),
.B(n_132),
.Y(n_1445)
);

O2A1O1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1278),
.A2(n_133),
.B(n_134),
.C(n_135),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1237),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1267),
.B(n_133),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1187),
.A2(n_349),
.B(n_346),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1301),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1239),
.B(n_135),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1328),
.Y(n_1452)
);

INVx3_ASAP7_75t_SL g1453 ( 
.A(n_1288),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1273),
.Y(n_1454)
);

AO32x1_ASAP7_75t_L g1455 ( 
.A1(n_1238),
.A2(n_136),
.A3(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1297),
.A2(n_136),
.B(n_137),
.C(n_138),
.Y(n_1456)
);

BUFx5_ASAP7_75t_L g1457 ( 
.A(n_1259),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1329),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1292),
.Y(n_1459)
);

AOI33xp33_ASAP7_75t_L g1460 ( 
.A1(n_1231),
.A2(n_140),
.A3(n_141),
.B1(n_142),
.B2(n_143),
.B3(n_144),
.Y(n_1460)
);

NOR2xp67_ASAP7_75t_SL g1461 ( 
.A(n_1305),
.B(n_140),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1193),
.B(n_141),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1360),
.Y(n_1463)
);

NAND2x1p5_ASAP7_75t_L g1464 ( 
.A(n_1385),
.B(n_1283),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1347),
.Y(n_1465)
);

BUFx8_ASAP7_75t_SL g1466 ( 
.A(n_1382),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_1353),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1458),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1418),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1332),
.Y(n_1470)
);

INVx1_ASAP7_75t_SL g1471 ( 
.A(n_1339),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1343),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1362),
.Y(n_1473)
);

INVx4_ASAP7_75t_L g1474 ( 
.A(n_1385),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1389),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1431),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1341),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1349),
.Y(n_1478)
);

BUFx2_ASAP7_75t_SL g1479 ( 
.A(n_1387),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1409),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1357),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1453),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1351),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1392),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1418),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1360),
.Y(n_1486)
);

NAND2x1p5_ASAP7_75t_L g1487 ( 
.A(n_1385),
.B(n_1232),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1400),
.A2(n_1199),
.B1(n_1192),
.B2(n_1221),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1374),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1340),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1418),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1440),
.B(n_1241),
.Y(n_1492)
);

INVx4_ASAP7_75t_L g1493 ( 
.A(n_1360),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1371),
.Y(n_1494)
);

BUFx2_ASAP7_75t_SL g1495 ( 
.A(n_1443),
.Y(n_1495)
);

INVx5_ASAP7_75t_L g1496 ( 
.A(n_1371),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1392),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1444),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1371),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1397),
.Y(n_1500)
);

BUFx4f_ASAP7_75t_SL g1501 ( 
.A(n_1435),
.Y(n_1501)
);

OR2x6_ASAP7_75t_L g1502 ( 
.A(n_1420),
.B(n_1308),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1394),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1420),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1450),
.Y(n_1505)
);

INVx6_ASAP7_75t_L g1506 ( 
.A(n_1337),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1403),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1425),
.B(n_1213),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1350),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1420),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1337),
.Y(n_1511)
);

BUFx12f_ASAP7_75t_L g1512 ( 
.A(n_1399),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1338),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1377),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1334),
.Y(n_1515)
);

BUFx4_ASAP7_75t_SL g1516 ( 
.A(n_1396),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1396),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1342),
.B(n_1255),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1447),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1439),
.A2(n_1451),
.B1(n_1412),
.B2(n_1361),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1433),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1378),
.Y(n_1522)
);

INVx4_ASAP7_75t_L g1523 ( 
.A(n_1432),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_SL g1524 ( 
.A(n_1459),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1383),
.Y(n_1525)
);

INVx6_ASAP7_75t_L g1526 ( 
.A(n_1363),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1410),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1358),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1415),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1436),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1427),
.Y(n_1531)
);

INVx3_ASAP7_75t_SL g1532 ( 
.A(n_1370),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1359),
.B(n_1315),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1346),
.Y(n_1534)
);

NOR2x1_ASAP7_75t_R g1535 ( 
.A(n_1417),
.B(n_1316),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1375),
.Y(n_1536)
);

BUFx4f_ASAP7_75t_L g1537 ( 
.A(n_1386),
.Y(n_1537)
);

BUFx2_ASAP7_75t_SL g1538 ( 
.A(n_1445),
.Y(n_1538)
);

INVx5_ASAP7_75t_L g1539 ( 
.A(n_1398),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1438),
.Y(n_1540)
);

BUFx16f_ASAP7_75t_R g1541 ( 
.A(n_1355),
.Y(n_1541)
);

OAI22xp33_ASAP7_75t_SL g1542 ( 
.A1(n_1344),
.A2(n_1269),
.B1(n_1266),
.B2(n_1275),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1373),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1448),
.Y(n_1544)
);

INVx3_ASAP7_75t_SL g1545 ( 
.A(n_1380),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1368),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1354),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_SL g1548 ( 
.A(n_1454),
.Y(n_1548)
);

INVx5_ASAP7_75t_L g1549 ( 
.A(n_1452),
.Y(n_1549)
);

BUFx2_ASAP7_75t_R g1550 ( 
.A(n_1421),
.Y(n_1550)
);

INVx5_ASAP7_75t_L g1551 ( 
.A(n_1393),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1365),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1333),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1401),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1426),
.B(n_1188),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1430),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1404),
.Y(n_1557)
);

BUFx12f_ASAP7_75t_L g1558 ( 
.A(n_1366),
.Y(n_1558)
);

INVx5_ASAP7_75t_L g1559 ( 
.A(n_1428),
.Y(n_1559)
);

INVx8_ASAP7_75t_L g1560 ( 
.A(n_1423),
.Y(n_1560)
);

CKINVDCx11_ASAP7_75t_R g1561 ( 
.A(n_1379),
.Y(n_1561)
);

CKINVDCx14_ASAP7_75t_R g1562 ( 
.A(n_1407),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1384),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1429),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1381),
.B(n_1302),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1352),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1336),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1462),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1461),
.A2(n_1216),
.B1(n_1209),
.B2(n_1321),
.Y(n_1569)
);

INVx4_ASAP7_75t_L g1570 ( 
.A(n_1457),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1442),
.Y(n_1571)
);

BUFx2_ASAP7_75t_SL g1572 ( 
.A(n_1548),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1478),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1544),
.B(n_1441),
.Y(n_1574)
);

O2A1O1Ixp33_ASAP7_75t_SL g1575 ( 
.A1(n_1492),
.A2(n_1335),
.B(n_1369),
.C(n_1331),
.Y(n_1575)
);

AOI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1520),
.A2(n_1348),
.B1(n_1356),
.B2(n_1402),
.C(n_1414),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_L g1577 ( 
.A(n_1528),
.B(n_1408),
.C(n_1330),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1558),
.B(n_1476),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1479),
.B(n_1413),
.Y(n_1579)
);

O2A1O1Ixp33_ASAP7_75t_SL g1580 ( 
.A1(n_1483),
.A2(n_1434),
.B(n_1372),
.C(n_1364),
.Y(n_1580)
);

NAND2x1p5_ASAP7_75t_L g1581 ( 
.A(n_1496),
.B(n_1388),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1471),
.Y(n_1582)
);

AO21x2_ASAP7_75t_L g1583 ( 
.A1(n_1555),
.A2(n_1411),
.B(n_1376),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1488),
.A2(n_1422),
.B(n_1345),
.Y(n_1584)
);

AO21x2_ASAP7_75t_L g1585 ( 
.A1(n_1468),
.A2(n_1449),
.B(n_1437),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1472),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1468),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1498),
.B(n_1505),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1519),
.A2(n_1367),
.B(n_1181),
.Y(n_1589)
);

NAND2x1p5_ASAP7_75t_L g1590 ( 
.A(n_1496),
.B(n_1523),
.Y(n_1590)
);

AOI21xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1560),
.A2(n_1424),
.B(n_1416),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1507),
.Y(n_1592)
);

O2A1O1Ixp33_ASAP7_75t_SL g1593 ( 
.A1(n_1508),
.A2(n_1456),
.B(n_1446),
.C(n_1395),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_R g1594 ( 
.A(n_1490),
.B(n_1457),
.Y(n_1594)
);

AOI21xp33_ASAP7_75t_L g1595 ( 
.A1(n_1535),
.A2(n_1391),
.B(n_1405),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_SL g1596 ( 
.A1(n_1552),
.A2(n_1419),
.B(n_1406),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1515),
.B(n_356),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1547),
.B(n_1460),
.Y(n_1598)
);

OAI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1537),
.A2(n_1390),
.B1(n_1176),
.B2(n_1455),
.C(n_1457),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1517),
.B(n_357),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1556),
.B(n_143),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1566),
.B(n_1557),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1514),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1480),
.Y(n_1604)
);

OR2x6_ASAP7_75t_L g1605 ( 
.A(n_1479),
.B(n_1455),
.Y(n_1605)
);

O2A1O1Ixp33_ASAP7_75t_SL g1606 ( 
.A1(n_1541),
.A2(n_145),
.B(n_146),
.C(n_147),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1540),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1521),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1534),
.B(n_146),
.Y(n_1609)
);

AO21x2_ASAP7_75t_L g1610 ( 
.A1(n_1554),
.A2(n_148),
.B(n_150),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1565),
.A2(n_413),
.B(n_456),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1517),
.A2(n_412),
.B(n_455),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_SL g1613 ( 
.A1(n_1562),
.A2(n_1553),
.B1(n_1548),
.B2(n_1564),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1568),
.B(n_358),
.Y(n_1614)
);

A2O1A1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1563),
.A2(n_150),
.B(n_151),
.C(n_153),
.Y(n_1615)
);

OAI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1539),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1511),
.B(n_360),
.Y(n_1617)
);

NAND3xp33_ASAP7_75t_L g1618 ( 
.A(n_1561),
.B(n_154),
.C(n_155),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1569),
.A2(n_415),
.B(n_452),
.Y(n_1619)
);

AO31x2_ASAP7_75t_L g1620 ( 
.A1(n_1570),
.A2(n_414),
.A3(n_448),
.B(n_445),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1549),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1522),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1549),
.Y(n_1623)
);

AO21x1_ASAP7_75t_L g1624 ( 
.A1(n_1542),
.A2(n_156),
.B(n_157),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1481),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1527),
.A2(n_1540),
.B(n_1487),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1470),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1503),
.Y(n_1628)
);

AOI222xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1509),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.C1(n_162),
.C2(n_163),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1587),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1626),
.Y(n_1631)
);

NAND2x1p5_ASAP7_75t_L g1632 ( 
.A(n_1621),
.B(n_1623),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1587),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1592),
.B(n_1567),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1621),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1607),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1623),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1625),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1590),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1603),
.B(n_1502),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1579),
.Y(n_1641)
);

BUFx4_ASAP7_75t_R g1642 ( 
.A(n_1628),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1627),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1573),
.Y(n_1644)
);

INVx5_ASAP7_75t_L g1645 ( 
.A(n_1579),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1585),
.B(n_1554),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1622),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1620),
.B(n_1502),
.Y(n_1648)
);

AO21x2_ASAP7_75t_L g1649 ( 
.A1(n_1584),
.A2(n_1533),
.B(n_1538),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1589),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1610),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1620),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1588),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1576),
.A2(n_1506),
.B1(n_1545),
.B2(n_1482),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1620),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1602),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1598),
.B(n_1530),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_SL g1658 ( 
.A(n_1645),
.B(n_1550),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1633),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1630),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1643),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1630),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1642),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1630),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1654),
.B(n_1629),
.C(n_1577),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1653),
.B(n_1582),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1636),
.B(n_1613),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1646),
.B(n_1609),
.Y(n_1668)
);

OAI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1651),
.A2(n_1618),
.B(n_1591),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1648),
.A2(n_1614),
.B(n_1616),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1649),
.A2(n_1624),
.B1(n_1538),
.B2(n_1559),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1656),
.B(n_1546),
.Y(n_1672)
);

OR2x6_ASAP7_75t_L g1673 ( 
.A(n_1648),
.B(n_1641),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_R g1674 ( 
.A(n_1641),
.B(n_1467),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1635),
.Y(n_1675)
);

NAND2xp33_ASAP7_75t_R g1676 ( 
.A(n_1646),
.B(n_1594),
.Y(n_1676)
);

XNOR2xp5_ASAP7_75t_L g1677 ( 
.A(n_1657),
.B(n_1465),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_SL g1678 ( 
.A(n_1645),
.B(n_1523),
.Y(n_1678)
);

CKINVDCx11_ASAP7_75t_R g1679 ( 
.A(n_1641),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1638),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1635),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1656),
.B(n_1543),
.Y(n_1682)
);

OR2x6_ASAP7_75t_L g1683 ( 
.A(n_1673),
.B(n_1648),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1661),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1660),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1659),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1668),
.B(n_1649),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1679),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1681),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1673),
.B(n_1649),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1661),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1673),
.B(n_1631),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1660),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1662),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1662),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1664),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1664),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1667),
.B(n_1635),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1666),
.B(n_1634),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1688),
.B(n_1674),
.Y(n_1700)
);

OA21x2_ASAP7_75t_L g1701 ( 
.A1(n_1685),
.A2(n_1669),
.B(n_1650),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1684),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1685),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1690),
.A2(n_1665),
.B(n_1670),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1688),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1683),
.A2(n_1671),
.B1(n_1645),
.B2(n_1663),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1689),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1703),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1704),
.A2(n_1671),
.B1(n_1645),
.B2(n_1683),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1705),
.B(n_1692),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1702),
.B(n_1687),
.Y(n_1711)
);

OAI211xp5_ASAP7_75t_L g1712 ( 
.A1(n_1700),
.A2(n_1606),
.B(n_1674),
.C(n_1615),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1710),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1711),
.B(n_1702),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1708),
.B(n_1691),
.Y(n_1715)
);

NAND4xp75_ASAP7_75t_L g1716 ( 
.A(n_1712),
.B(n_1701),
.C(n_1690),
.D(n_1692),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1709),
.B(n_1707),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1710),
.B(n_1698),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1713),
.B(n_1699),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1714),
.B(n_1701),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1718),
.B(n_1466),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1721),
.B(n_1716),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1719),
.B(n_1715),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_L g1724 ( 
.A(n_1722),
.B(n_1717),
.C(n_1720),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1724),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1725),
.B(n_1723),
.Y(n_1726)
);

AOI21xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1725),
.A2(n_1560),
.B(n_1578),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1726),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1727),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1728),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1729),
.A2(n_1608),
.B(n_1706),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1728),
.Y(n_1732)
);

A2O1A1Ixp33_ASAP7_75t_L g1733 ( 
.A1(n_1730),
.A2(n_1597),
.B(n_1572),
.C(n_1586),
.Y(n_1733)
);

AOI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1732),
.A2(n_1524),
.B1(n_1604),
.B2(n_1572),
.C(n_1473),
.Y(n_1734)
);

AOI211xp5_ASAP7_75t_L g1735 ( 
.A1(n_1731),
.A2(n_1532),
.B(n_1601),
.C(n_1475),
.Y(n_1735)
);

AOI221x1_ASAP7_75t_L g1736 ( 
.A1(n_1733),
.A2(n_1734),
.B1(n_1735),
.B2(n_161),
.C(n_162),
.Y(n_1736)
);

OAI211xp5_ASAP7_75t_L g1737 ( 
.A1(n_1734),
.A2(n_1489),
.B(n_1539),
.C(n_1474),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1735),
.B(n_1677),
.Y(n_1738)
);

AOI31xp33_ASAP7_75t_L g1739 ( 
.A1(n_1734),
.A2(n_1524),
.A3(n_1617),
.B(n_1501),
.Y(n_1739)
);

OAI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1734),
.A2(n_1658),
.B1(n_1536),
.B2(n_1526),
.C(n_1539),
.Y(n_1740)
);

OAI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1734),
.A2(n_1526),
.B1(n_1678),
.B2(n_1676),
.C(n_1672),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1734),
.A2(n_1639),
.B1(n_1512),
.B2(n_1631),
.Y(n_1742)
);

NOR3xp33_ASAP7_75t_SL g1743 ( 
.A(n_1737),
.B(n_1676),
.C(n_158),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1739),
.A2(n_1575),
.B1(n_1684),
.B2(n_1595),
.C(n_1600),
.Y(n_1744)
);

AOI32xp33_ASAP7_75t_L g1745 ( 
.A1(n_1742),
.A2(n_1617),
.A3(n_1600),
.B1(n_1474),
.B2(n_1639),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1736),
.B(n_1682),
.Y(n_1746)
);

AND4x2_ASAP7_75t_L g1747 ( 
.A(n_1740),
.B(n_160),
.C(n_163),
.D(n_164),
.Y(n_1747)
);

OAI21xp33_ASAP7_75t_SL g1748 ( 
.A1(n_1738),
.A2(n_1689),
.B(n_1683),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1741),
.A2(n_1495),
.B1(n_1496),
.B2(n_1493),
.Y(n_1749)
);

AOI222xp33_ASAP7_75t_L g1750 ( 
.A1(n_1737),
.A2(n_1651),
.B1(n_1571),
.B2(n_1559),
.C1(n_1599),
.C2(n_1645),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1736),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1736),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1751),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1752),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1743),
.A2(n_1571),
.B1(n_1639),
.B2(n_1645),
.Y(n_1755)
);

AO22x2_ASAP7_75t_L g1756 ( 
.A1(n_1746),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1748),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1749),
.Y(n_1758)
);

NOR4xp75_ASAP7_75t_L g1759 ( 
.A(n_1747),
.B(n_166),
.C(n_168),
.D(n_169),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1744),
.B(n_1634),
.Y(n_1760)
);

OAI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1750),
.A2(n_1612),
.B(n_1611),
.Y(n_1761)
);

NAND4xp75_ASAP7_75t_L g1762 ( 
.A(n_1745),
.B(n_168),
.C(n_169),
.D(n_170),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1751),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1751),
.B(n_170),
.Y(n_1764)
);

NAND4xp75_ASAP7_75t_L g1765 ( 
.A(n_1751),
.B(n_172),
.C(n_1516),
.D(n_1574),
.Y(n_1765)
);

INVxp67_ASAP7_75t_SL g1766 ( 
.A(n_1751),
.Y(n_1766)
);

NOR3x1_ASAP7_75t_L g1767 ( 
.A(n_1751),
.B(n_172),
.C(n_1499),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_SL g1768 ( 
.A(n_1751),
.B(n_1493),
.Y(n_1768)
);

NAND5xp2_ASAP7_75t_L g1769 ( 
.A(n_1751),
.B(n_1464),
.C(n_1581),
.D(n_1593),
.E(n_1632),
.Y(n_1769)
);

NOR2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1751),
.B(n_1486),
.Y(n_1770)
);

NAND2x1p5_ASAP7_75t_L g1771 ( 
.A(n_1751),
.B(n_1513),
.Y(n_1771)
);

INVx2_ASAP7_75t_SL g1772 ( 
.A(n_1751),
.Y(n_1772)
);

NOR2x1_ASAP7_75t_L g1773 ( 
.A(n_1751),
.B(n_1495),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1751),
.Y(n_1774)
);

NOR3xp33_ASAP7_75t_L g1775 ( 
.A(n_1751),
.B(n_1531),
.C(n_1485),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1751),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1751),
.A2(n_1571),
.B(n_1500),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1751),
.B(n_1529),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_1756),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1753),
.Y(n_1780)
);

NOR2x1_ASAP7_75t_L g1781 ( 
.A(n_1764),
.B(n_1494),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1759),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1772),
.B(n_1766),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1756),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1754),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1757),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1765),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_R g1788 ( 
.A(n_1763),
.B(n_361),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1773),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1767),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1774),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1776),
.B(n_1768),
.Y(n_1792)
);

INVx1_ASAP7_75t_SL g1793 ( 
.A(n_1762),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1775),
.A2(n_1525),
.B1(n_1513),
.B2(n_1632),
.C(n_1510),
.Y(n_1794)
);

NOR4xp75_ASAP7_75t_L g1795 ( 
.A(n_1778),
.B(n_1504),
.C(n_1491),
.D(n_1485),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1771),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1770),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1758),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1777),
.B(n_1477),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_R g1800 ( 
.A(n_1760),
.B(n_362),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1755),
.Y(n_1801)
);

INVx1_ASAP7_75t_SL g1802 ( 
.A(n_1761),
.Y(n_1802)
);

BUFx2_ASAP7_75t_L g1803 ( 
.A(n_1769),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_R g1804 ( 
.A(n_1772),
.B(n_367),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1759),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1759),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1756),
.Y(n_1807)
);

XNOR2xp5_ASAP7_75t_L g1808 ( 
.A(n_1782),
.B(n_1805),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1790),
.B(n_1637),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1779),
.B(n_1513),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1784),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_L g1812 ( 
.A(n_1786),
.B(n_1463),
.C(n_1510),
.Y(n_1812)
);

OAI22x1_ASAP7_75t_L g1813 ( 
.A1(n_1806),
.A2(n_1632),
.B1(n_1504),
.B2(n_1491),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1780),
.Y(n_1814)
);

XNOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1785),
.B(n_368),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_SL g1816 ( 
.A1(n_1807),
.A2(n_1463),
.B1(n_1510),
.B2(n_1506),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1783),
.Y(n_1817)
);

AOI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1791),
.A2(n_1463),
.B1(n_1681),
.B2(n_1637),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1793),
.A2(n_1637),
.B1(n_1686),
.B2(n_1675),
.Y(n_1819)
);

AO21x2_ASAP7_75t_L g1820 ( 
.A1(n_1792),
.A2(n_369),
.B(n_370),
.Y(n_1820)
);

OAI22x1_ASAP7_75t_L g1821 ( 
.A1(n_1787),
.A2(n_1469),
.B1(n_1559),
.B2(n_1497),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1789),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1801),
.A2(n_1469),
.B1(n_1631),
.B2(n_1605),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1780),
.Y(n_1824)
);

AOI22x1_ASAP7_75t_L g1825 ( 
.A1(n_1798),
.A2(n_1484),
.B1(n_374),
.B2(n_375),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1780),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1796),
.A2(n_1596),
.B(n_1580),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1781),
.Y(n_1828)
);

AO21x1_ASAP7_75t_L g1829 ( 
.A1(n_1797),
.A2(n_1697),
.B(n_1696),
.Y(n_1829)
);

AO22x2_ASAP7_75t_L g1830 ( 
.A1(n_1802),
.A2(n_1695),
.B1(n_1694),
.B2(n_1693),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1803),
.Y(n_1831)
);

AOI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1794),
.A2(n_1648),
.B1(n_1605),
.B2(n_1640),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1799),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_SL g1834 ( 
.A1(n_1788),
.A2(n_1518),
.B1(n_1655),
.B2(n_1652),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1804),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1800),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1795),
.A2(n_1652),
.B1(n_1655),
.B2(n_1551),
.Y(n_1837)
);

CKINVDCx20_ASAP7_75t_R g1838 ( 
.A(n_1808),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1811),
.A2(n_1619),
.B(n_1518),
.Y(n_1839)
);

XNOR2xp5_ASAP7_75t_L g1840 ( 
.A(n_1815),
.B(n_371),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1826),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1831),
.B(n_377),
.Y(n_1842)
);

OA21x2_ASAP7_75t_L g1843 ( 
.A1(n_1810),
.A2(n_379),
.B(n_381),
.Y(n_1843)
);

OAI22xp33_ASAP7_75t_SL g1844 ( 
.A1(n_1822),
.A2(n_1817),
.B1(n_1825),
.B2(n_1814),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1824),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1820),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_SL g1847 ( 
.A1(n_1836),
.A2(n_1551),
.B1(n_1640),
.B2(n_1533),
.Y(n_1847)
);

OAI211xp5_ASAP7_75t_L g1848 ( 
.A1(n_1828),
.A2(n_382),
.B(n_383),
.C(n_385),
.Y(n_1848)
);

OA22x2_ASAP7_75t_L g1849 ( 
.A1(n_1809),
.A2(n_1640),
.B1(n_1644),
.B2(n_1647),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1812),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1835),
.B(n_1640),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1833),
.Y(n_1852)
);

OAI22x1_ASAP7_75t_L g1853 ( 
.A1(n_1818),
.A2(n_1551),
.B1(n_1680),
.B2(n_1644),
.Y(n_1853)
);

NOR2x1_ASAP7_75t_L g1854 ( 
.A(n_1819),
.B(n_386),
.Y(n_1854)
);

AO22x2_ASAP7_75t_L g1855 ( 
.A1(n_1816),
.A2(n_393),
.B1(n_394),
.B2(n_395),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1843),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1846),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1838),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1841),
.Y(n_1859)
);

INVxp67_ASAP7_75t_SL g1860 ( 
.A(n_1842),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1840),
.Y(n_1861)
);

INVxp67_ASAP7_75t_SL g1862 ( 
.A(n_1852),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1851),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1845),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1854),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1844),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1850),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1855),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1862),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1858),
.A2(n_1855),
.B1(n_1832),
.B2(n_1834),
.Y(n_1870)
);

INVx1_ASAP7_75t_SL g1871 ( 
.A(n_1868),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1862),
.A2(n_1848),
.B1(n_1827),
.B2(n_1847),
.Y(n_1872)
);

OR3x1_ASAP7_75t_L g1873 ( 
.A(n_1866),
.B(n_1821),
.C(n_1853),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1859),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1864),
.Y(n_1875)
);

OAI21x1_ASAP7_75t_L g1876 ( 
.A1(n_1869),
.A2(n_1856),
.B(n_1865),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1874),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_SL g1878 ( 
.A1(n_1873),
.A2(n_1863),
.B1(n_1867),
.B2(n_1857),
.Y(n_1878)
);

NAND5xp2_ASAP7_75t_L g1879 ( 
.A(n_1877),
.B(n_1875),
.C(n_1861),
.D(n_1860),
.E(n_1871),
.Y(n_1879)
);

INVx4_ASAP7_75t_L g1880 ( 
.A(n_1878),
.Y(n_1880)
);

AOI211xp5_ASAP7_75t_L g1881 ( 
.A1(n_1876),
.A2(n_1872),
.B(n_1870),
.C(n_1829),
.Y(n_1881)
);

XOR2x2_ASAP7_75t_L g1882 ( 
.A(n_1878),
.B(n_1849),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1880),
.Y(n_1883)
);

OAI222xp33_ASAP7_75t_L g1884 ( 
.A1(n_1879),
.A2(n_1823),
.B1(n_1837),
.B2(n_1813),
.C1(n_1830),
.C2(n_1839),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1883),
.A2(n_1882),
.B1(n_1881),
.B2(n_1830),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1884),
.A2(n_1583),
.B1(n_1647),
.B2(n_398),
.Y(n_1886)
);

AO21x2_ASAP7_75t_L g1887 ( 
.A1(n_1885),
.A2(n_396),
.B(n_397),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1887),
.A2(n_1886),
.B1(n_401),
.B2(n_402),
.Y(n_1888)
);

AOI211xp5_ASAP7_75t_L g1889 ( 
.A1(n_1888),
.A2(n_400),
.B(n_405),
.C(n_407),
.Y(n_1889)
);


endmodule