module fake_jpeg_27857_n_187 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_17),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_16),
.B1(n_21),
.B2(n_20),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_29),
.B1(n_24),
.B2(n_25),
.Y(n_45)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_19),
.C(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_42),
.B1(n_35),
.B2(n_27),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_32),
.Y(n_46)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

CKINVDCx11_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_56),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_28),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_33),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_70),
.C(n_23),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_34),
.B(n_23),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_71),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_40),
.C(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_51),
.B1(n_46),
.B2(n_47),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_78),
.B1(n_24),
.B2(n_25),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_39),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_36),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_50),
.B1(n_37),
.B2(n_34),
.Y(n_78)
);

OA21x2_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_58),
.B(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_34),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_84),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_35),
.B1(n_43),
.B2(n_36),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_68),
.B1(n_62),
.B2(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_61),
.B(n_43),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_68),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_62),
.B1(n_68),
.B2(n_57),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_90),
.B1(n_98),
.B2(n_78),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_88),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_81),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_99),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_58),
.B1(n_65),
.B2(n_60),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_85),
.C(n_84),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_94),
.C(n_71),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_105),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_108),
.B1(n_24),
.B2(n_55),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_80),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_122),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_94),
.B1(n_95),
.B2(n_89),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_127),
.B1(n_48),
.B2(n_38),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_109),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_65),
.C(n_31),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_129),
.C(n_117),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_65),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_52),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_69),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_54),
.B1(n_48),
.B2(n_55),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_107),
.B1(n_109),
.B2(n_54),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_31),
.C(n_69),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_139),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_140),
.B(n_22),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_20),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_66),
.B1(n_13),
.B2(n_12),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_66),
.C(n_19),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_66),
.C(n_38),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_R g144 ( 
.A(n_133),
.B(n_122),
.C(n_115),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_13),
.C(n_12),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_152),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_148),
.C(n_27),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_0),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_147),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_22),
.C(n_18),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_143),
.B(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_157),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_142),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_156),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

OAI21x1_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_1),
.B(n_2),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_29),
.B1(n_2),
.B2(n_3),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_162),
.B1(n_159),
.B2(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_149),
.C(n_153),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_22),
.C(n_18),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_166),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_168),
.B(n_169),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_160),
.B1(n_3),
.B2(n_4),
.Y(n_166)
);

OAI221xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_18),
.B1(n_22),
.B2(n_5),
.C(n_6),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_162),
.A2(n_2),
.B(n_4),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_5),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_171),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_176),
.C(n_7),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_6),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_170),
.A2(n_7),
.B(n_8),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

HB1xp67_ASAP7_75t_SL g181 ( 
.A(n_178),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_9),
.C(n_10),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_175),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_183),
.C(n_9),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_177),
.B(n_10),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_184),
.A2(n_185),
.B(n_182),
.C(n_11),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_10),
.Y(n_187)
);


endmodule