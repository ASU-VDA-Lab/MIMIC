module fake_jpeg_5322_n_230 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_SL g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_32),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_38),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_56),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_18),
.B1(n_29),
.B2(n_25),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_35),
.B1(n_37),
.B2(n_30),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_29),
.B1(n_19),
.B2(n_25),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_29),
.B1(n_25),
.B2(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_28),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_33),
.A2(n_17),
.B1(n_20),
.B2(n_26),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_23),
.B1(n_20),
.B2(n_17),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_64),
.Y(n_88)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_45),
.B1(n_51),
.B2(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_48),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_22),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_14),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_81),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_34),
.C(n_31),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_52),
.C(n_59),
.Y(n_82)
);

AO22x1_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_38),
.B1(n_31),
.B2(n_27),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_46),
.B(n_58),
.C(n_38),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_23),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_0),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_91),
.C(n_61),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_89),
.B(n_98),
.C(n_64),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_50),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_85),
.C(n_97),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_41),
.B(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_99),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_67),
.A2(n_78),
.B1(n_75),
.B2(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_41),
.B1(n_55),
.B2(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_43),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_66),
.A3(n_73),
.B1(n_76),
.B2(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_101),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_22),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_54),
.B1(n_53),
.B2(n_38),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_77),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_77),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_43),
.B1(n_54),
.B2(n_74),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_123),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_115),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_117),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_97),
.B1(n_102),
.B2(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_84),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_116),
.A2(n_84),
.B(n_89),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_124),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_121),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_80),
.C(n_43),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_72),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_113),
.C(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_142),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_96),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_137),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_134),
.A2(n_138),
.B1(n_142),
.B2(n_131),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_97),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_105),
.C(n_122),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_100),
.B1(n_102),
.B2(n_93),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_118),
.B1(n_109),
.B2(n_117),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_103),
.B(n_93),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_81),
.B1(n_77),
.B2(n_87),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_72),
.B1(n_27),
.B2(n_24),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_139),
.B(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_144),
.Y(n_162)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_149),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_148),
.B(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_152),
.B1(n_134),
.B2(n_137),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_106),
.B1(n_110),
.B2(n_112),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_159),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_154),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_140),
.C(n_144),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_129),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_126),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_24),
.B1(n_15),
.B2(n_22),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_163),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_86),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_127),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_165),
.C(n_168),
.Y(n_179)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_153),
.B1(n_150),
.B2(n_151),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_135),
.C(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_0),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_130),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_147),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_177),
.B(n_127),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_187),
.C(n_188),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_185),
.Y(n_199)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_177),
.A2(n_152),
.B1(n_147),
.B2(n_150),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_172),
.B1(n_164),
.B2(n_174),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_191),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_8),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_24),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_24),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_190),
.C(n_170),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_15),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_184),
.B(n_171),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_195),
.C(n_198),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_202),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_190),
.B(n_175),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_1),
.Y(n_210)
);

AO22x1_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_178),
.B1(n_0),
.B2(n_2),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_201),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_178),
.C(n_2),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_179),
.C(n_2),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_210),
.B(n_194),
.Y(n_211)
);

AOI31xp67_ASAP7_75t_SL g205 ( 
.A1(n_193),
.A2(n_1),
.A3(n_3),
.B(n_5),
.Y(n_205)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_6),
.B(n_7),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_209),
.Y(n_212)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_203),
.B(n_202),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_216),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_5),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_215),
.B(n_217),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_7),
.B(n_9),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_11),
.B(n_12),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_10),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_12),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_10),
.C(n_11),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_223),
.A2(n_224),
.B(n_226),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_220),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_227),
.A2(n_13),
.B(n_228),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_13),
.Y(n_230)
);


endmodule