module fake_jpeg_30278_n_179 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_27),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_0),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_12),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_79),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_1),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_74),
.Y(n_88)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_95),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_55),
.B1(n_72),
.B2(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_89),
.B1(n_70),
.B2(n_55),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_70),
.B(n_60),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_2),
.B(n_3),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_59),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_68),
.B1(n_54),
.B2(n_64),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_62),
.Y(n_95)
);

CKINVDCx6p67_ASAP7_75t_R g99 ( 
.A(n_78),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_80),
.B1(n_55),
.B2(n_72),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_107),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_67),
.B1(n_66),
.B2(n_65),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_96),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_71),
.B1(n_63),
.B2(n_59),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_2),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_6),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_59),
.B(n_3),
.C(n_4),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_9),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_4),
.B(n_5),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_93),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_26),
.B1(n_49),
.B2(n_48),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_127)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_124),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_6),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_11),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_11),
.B(n_13),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_112),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_20),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_146)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_21),
.B1(n_23),
.B2(n_28),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_141),
.A2(n_152),
.B1(n_157),
.B2(n_43),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_133),
.B(n_126),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_146),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_147),
.B(n_148),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_135),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_120),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_46),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_132),
.B1(n_130),
.B2(n_119),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_40),
.C(n_41),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_141),
.C(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_150),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_151),
.B1(n_149),
.B2(n_154),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_160),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_169),
.A2(n_158),
.B1(n_161),
.B2(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_172),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_167),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_170),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_163),
.B(n_168),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_172),
.Y(n_179)
);


endmodule