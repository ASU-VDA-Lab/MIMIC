module fake_jpeg_2131_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_56),
.Y(n_60)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_50),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_51),
.B1(n_52),
.B2(n_39),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_72),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_45),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_74),
.Y(n_94)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_58),
.B1(n_49),
.B2(n_44),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_56),
.B1(n_59),
.B2(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_78),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_59),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_60),
.C(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_73),
.B(n_72),
.C(n_80),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_87),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_67),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_19),
.C(n_36),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_49),
.B1(n_48),
.B2(n_42),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_93),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_70),
.B1(n_20),
.B2(n_21),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_99),
.B1(n_98),
.B2(n_86),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_0),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_1),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_2),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_105),
.B(n_106),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_3),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_109),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_22),
.C(n_34),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_117),
.C(n_15),
.Y(n_124)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_112),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_27),
.B1(n_30),
.B2(n_29),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_4),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_96),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_116),
.B(n_5),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_26),
.C(n_33),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_17),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_127),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_16),
.B(n_31),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_122),
.B(n_125),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_117),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_14),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.Y(n_140)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_120),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_139),
.B(n_141),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_131),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_132),
.B(n_118),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_123),
.C(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_144),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_143),
.B(n_110),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_124),
.B1(n_136),
.B2(n_28),
.Y(n_148)
);

AOI221x1_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_37),
.B1(n_136),
.B2(n_7),
.C(n_8),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_112),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_5),
.Y(n_151)
);


endmodule