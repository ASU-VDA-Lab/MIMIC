module fake_netlist_6_4932_n_1769 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1769);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1769;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_50),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_43),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_83),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_27),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_128),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_80),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_121),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_9),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_29),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_105),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_76),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_21),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_123),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_16),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_31),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_56),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_70),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_20),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_30),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_49),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_50),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_10),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_29),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_5),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_36),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_92),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_26),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_114),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_7),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_20),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_91),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_148),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_85),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_33),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_27),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_21),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_81),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_8),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_26),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_18),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_137),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_39),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_82),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_34),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_140),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_99),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_40),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_9),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_61),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_19),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_109),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_2),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_136),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_31),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_127),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_142),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_75),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_63),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_32),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_13),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_3),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_0),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_77),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_139),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_160),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_40),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_157),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_100),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_46),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_103),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_44),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_49),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_55),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_144),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_93),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_147),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_28),
.Y(n_250)
);

INVxp33_ASAP7_75t_SL g251 ( 
.A(n_73),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_13),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_52),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_129),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_51),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_122),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_10),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_5),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_23),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_62),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_159),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_12),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_161),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_6),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_33),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_130),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_88),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_34),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_24),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_58),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_110),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_47),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_67),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_36),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_74),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_6),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_64),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_32),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_145),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_44),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_16),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_37),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_117),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_72),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_118),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_39),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_19),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_42),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_15),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_43),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_156),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_146),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_45),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_104),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_41),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_14),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_71),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_151),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_150),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_12),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_47),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_119),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_106),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_54),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_38),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_87),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_7),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_0),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_3),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_158),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_8),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_37),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_15),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_22),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_138),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_48),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_18),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_65),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_162),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_120),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_141),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_111),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_42),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_187),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_250),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_165),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_250),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_250),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_250),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_250),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_166),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_250),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_195),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_197),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_250),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_181),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_221),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_214),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_237),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_193),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_193),
.Y(n_342)
);

INVxp33_ASAP7_75t_SL g343 ( 
.A(n_174),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_240),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_198),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_193),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_193),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_198),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_249),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_193),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_210),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_174),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_196),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_210),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_210),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_210),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_210),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_198),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_288),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_255),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_165),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_200),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_176),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_201),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_207),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_288),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_209),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_300),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_275),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_300),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_209),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_207),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_179),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_202),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_309),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_309),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_319),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_216),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_323),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_168),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_209),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_219),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_290),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_184),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_188),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_190),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_199),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_296),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_203),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_226),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_290),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_212),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_217),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_220),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_227),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_209),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_263),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_241),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_290),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_242),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_245),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_333),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_331),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_340),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_342),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_340),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_346),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_345),
.B(n_237),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_346),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_347),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_347),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_345),
.B(n_273),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_363),
.A2(n_297),
.B1(n_177),
.B2(n_316),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_361),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_325),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_350),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_327),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_372),
.B(n_310),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_327),
.Y(n_423)
);

INVx6_ASAP7_75t_L g424 ( 
.A(n_348),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_372),
.B(n_213),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_348),
.B(n_273),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_334),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_350),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_328),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_362),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_364),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_351),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_353),
.A2(n_251),
.B1(n_295),
.B2(n_235),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_374),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_378),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_328),
.B(n_204),
.Y(n_437)
);

INVxp33_ASAP7_75t_SL g438 ( 
.A(n_382),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_324),
.A2(n_264),
.B1(n_192),
.B2(n_233),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_329),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_354),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_329),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_L g444 ( 
.A(n_390),
.B(n_179),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_191),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_355),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_358),
.B(n_191),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_375),
.B(n_213),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_398),
.A2(n_180),
.B1(n_186),
.B2(n_239),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g450 ( 
.A(n_355),
.B(n_163),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_330),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_365),
.B(n_173),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_343),
.A2(n_251),
.B1(n_268),
.B2(n_265),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_388),
.B(n_230),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_337),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_330),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_332),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_356),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_339),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_332),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_375),
.B(n_269),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_335),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_358),
.B(n_189),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_356),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_357),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_357),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_326),
.B(n_205),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_335),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_352),
.B(n_178),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_336),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_336),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_367),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_367),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_379),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_383),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_472),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_410),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_472),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_376),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_405),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_475),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_338),
.C(n_391),
.Y(n_482)
);

NAND2x1p5_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_222),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_468),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_454),
.B(n_204),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_406),
.B(n_302),
.Y(n_486)
);

AO21x2_ASAP7_75t_L g487 ( 
.A1(n_445),
.A2(n_211),
.B(n_208),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_472),
.Y(n_488)
);

BUFx10_ASAP7_75t_L g489 ( 
.A(n_403),
.Y(n_489)
);

AO22x2_ASAP7_75t_L g490 ( 
.A1(n_417),
.A2(n_272),
.B1(n_269),
.B2(n_252),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_406),
.B(n_463),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_473),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_473),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_468),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_228),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_473),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_438),
.B(n_373),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_463),
.B(n_204),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_408),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_408),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_463),
.B(n_376),
.Y(n_502)
);

AO22x2_ASAP7_75t_L g503 ( 
.A1(n_449),
.A2(n_272),
.B1(n_313),
.B2(n_281),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_422),
.A2(n_257),
.B1(n_259),
.B2(n_274),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_419),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_419),
.Y(n_506)
);

OAI22xp33_ASAP7_75t_L g507 ( 
.A1(n_433),
.A2(n_293),
.B1(n_262),
.B2(n_185),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_471),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_421),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_427),
.B(n_399),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_444),
.A2(n_344),
.B1(n_349),
.B2(n_360),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_421),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_421),
.B(n_231),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_443),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_422),
.A2(n_326),
.B1(n_384),
.B2(n_385),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_453),
.B(n_204),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_419),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_443),
.B(n_236),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_405),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_450),
.B(n_204),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_423),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_443),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_423),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_423),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_429),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_443),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_430),
.B(n_369),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_467),
.A2(n_431),
.B1(n_434),
.B2(n_436),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_418),
.B(n_377),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_412),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_457),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_447),
.B(n_218),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_425),
.B(n_359),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_457),
.B(n_470),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_429),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_452),
.B(n_167),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_457),
.B(n_243),
.Y(n_538)
);

AND3x2_ASAP7_75t_L g539 ( 
.A(n_425),
.B(n_254),
.C(n_229),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_448),
.B(n_167),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_457),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_470),
.B(n_248),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_470),
.Y(n_543)
);

BUFx4f_ASAP7_75t_L g544 ( 
.A(n_437),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_470),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_437),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_429),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_405),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_405),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_459),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_440),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_440),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_440),
.Y(n_553)
);

OA22x2_ASAP7_75t_L g554 ( 
.A1(n_448),
.A2(n_461),
.B1(n_439),
.B2(n_401),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_451),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_412),
.B(n_253),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_451),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_451),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_447),
.B(n_224),
.Y(n_559)
);

OAI21xp33_ASAP7_75t_SL g560 ( 
.A1(n_461),
.A2(n_366),
.B(n_359),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_439),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_404),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_405),
.Y(n_563)
);

INVxp67_ASAP7_75t_SL g564 ( 
.A(n_456),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_412),
.B(n_256),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_456),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_412),
.A2(n_182),
.B1(n_238),
.B2(n_322),
.Y(n_567)
);

OAI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_416),
.A2(n_186),
.B1(n_180),
.B2(n_239),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_416),
.B(n_260),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_456),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_460),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_416),
.A2(n_183),
.B1(n_182),
.B2(n_322),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_416),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_426),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_405),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_426),
.A2(n_183),
.B1(n_175),
.B2(n_171),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_426),
.B(n_261),
.Y(n_577)
);

NOR2x1p5_ASAP7_75t_L g578 ( 
.A(n_474),
.B(n_307),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_428),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_426),
.A2(n_238),
.B1(n_175),
.B2(n_171),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_424),
.Y(n_581)
);

OAI22xp33_ASAP7_75t_L g582 ( 
.A1(n_474),
.A2(n_164),
.B1(n_234),
.B2(n_282),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_460),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_428),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_424),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_447),
.B(n_386),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_460),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_462),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_L g589 ( 
.A1(n_424),
.A2(n_232),
.B1(n_194),
.B2(n_206),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_462),
.Y(n_590)
);

NAND3xp33_ASAP7_75t_L g591 ( 
.A(n_447),
.B(n_244),
.C(n_223),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_462),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_402),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_424),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_424),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_402),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_407),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_407),
.B(n_366),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_409),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_409),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_411),
.B(n_379),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_411),
.B(n_380),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_413),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_437),
.A2(n_169),
.B1(n_170),
.B2(n_320),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_413),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_414),
.B(n_266),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_414),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_466),
.B(n_380),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_437),
.B(n_209),
.Y(n_609)
);

OAI22xp33_ASAP7_75t_L g610 ( 
.A1(n_415),
.A2(n_225),
.B1(n_215),
.B2(n_258),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_415),
.B(n_267),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_420),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_420),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_437),
.A2(n_169),
.B1(n_170),
.B2(n_315),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_466),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_428),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_432),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_432),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_442),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_465),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_465),
.B(n_246),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_442),
.B(n_270),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_458),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_L g624 ( 
.A(n_437),
.B(n_209),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_458),
.B(n_271),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_544),
.B(n_209),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_620),
.B(n_428),
.Y(n_627)
);

O2A1O1Ixp33_ASAP7_75t_L g628 ( 
.A1(n_516),
.A2(n_392),
.B(n_387),
.C(n_401),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_593),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_562),
.Y(n_630)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_540),
.B(n_286),
.C(n_289),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_573),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_573),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_531),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_507),
.B(n_393),
.C(n_400),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_593),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_477),
.B(n_315),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_561),
.B(n_387),
.Y(n_638)
);

NOR2xp67_ASAP7_75t_SL g639 ( 
.A(n_546),
.B(n_247),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_544),
.B(n_209),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_620),
.B(n_428),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_L g642 ( 
.A(n_485),
.B(n_394),
.C(n_400),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_477),
.B(n_318),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_597),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_598),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_597),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_598),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_SL g648 ( 
.A(n_546),
.B(n_291),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_L g649 ( 
.A(n_515),
.B(n_287),
.C(n_280),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_484),
.B(n_428),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_494),
.B(n_435),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_508),
.B(n_435),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_599),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_537),
.B(n_435),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_543),
.B(n_435),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_544),
.B(n_483),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_534),
.B(n_389),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_550),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_601),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_479),
.B(n_435),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_483),
.B(n_299),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_479),
.B(n_435),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_535),
.A2(n_437),
.B(n_321),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_516),
.A2(n_395),
.B(n_394),
.C(n_393),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_574),
.B(n_277),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_578),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_600),
.B(n_318),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_502),
.B(n_441),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_554),
.A2(n_172),
.B1(n_276),
.B2(n_278),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_600),
.B(n_605),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_601),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_605),
.B(n_279),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_510),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_599),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_602),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_602),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_574),
.B(n_320),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_502),
.B(n_441),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_482),
.B(n_301),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_586),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_554),
.A2(n_311),
.B1(n_305),
.B2(n_437),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_564),
.B(n_596),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_612),
.B(n_441),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_615),
.B(n_307),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_L g685 ( 
.A(n_504),
.B(n_314),
.C(n_308),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_586),
.Y(n_686)
);

BUFx2_ASAP7_75t_SL g687 ( 
.A(n_489),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_613),
.B(n_441),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_603),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_617),
.B(n_441),
.Y(n_690)
);

NOR2xp67_ASAP7_75t_L g691 ( 
.A(n_497),
.B(n_283),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_511),
.B(n_481),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_603),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_486),
.B(n_308),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_581),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_585),
.B(n_389),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_618),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_495),
.B(n_441),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_525),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_607),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_607),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_560),
.A2(n_395),
.B(n_392),
.C(n_370),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_619),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_487),
.B(n_446),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_546),
.B(n_509),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_619),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_487),
.B(n_446),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_487),
.B(n_446),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_623),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_623),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_595),
.B(n_284),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_546),
.B(n_285),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_476),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_534),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_485),
.B(n_312),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_585),
.B(n_368),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_608),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_608),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_567),
.B(n_312),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_546),
.B(n_512),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_476),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_550),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_478),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_529),
.B(n_292),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_608),
.B(n_370),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_608),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_539),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_556),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_514),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_478),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_530),
.B(n_294),
.Y(n_731)
);

NOR2xp67_ASAP7_75t_L g732 ( 
.A(n_528),
.B(n_298),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_522),
.Y(n_733)
);

O2A1O1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_621),
.A2(n_368),
.B(n_381),
.C(n_371),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_527),
.B(n_464),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_532),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_541),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_545),
.B(n_464),
.Y(n_738)
);

INVxp33_ASAP7_75t_L g739 ( 
.A(n_562),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_491),
.B(n_464),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_591),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_572),
.B(n_314),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_565),
.A2(n_306),
.B1(n_303),
.B2(n_304),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_491),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_488),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_513),
.B(n_518),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_488),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_538),
.B(n_464),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_492),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_492),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_569),
.A2(n_230),
.B1(n_464),
.B2(n_446),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_576),
.B(n_580),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_581),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_489),
.B(n_316),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_493),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_493),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_496),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_496),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_542),
.B(n_464),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_606),
.B(n_317),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_577),
.A2(n_625),
.B1(n_622),
.B2(n_611),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_551),
.B(n_446),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_568),
.B(n_230),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_553),
.B(n_396),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_555),
.B(n_396),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_489),
.Y(n_766)
);

NOR3xp33_ASAP7_75t_L g767 ( 
.A(n_582),
.B(n_317),
.C(n_381),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_557),
.B(n_371),
.Y(n_768)
);

AND2x2_ASAP7_75t_SL g769 ( 
.A(n_624),
.B(n_68),
.Y(n_769)
);

OA21x2_ASAP7_75t_L g770 ( 
.A1(n_498),
.A2(n_69),
.B(n_143),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_566),
.B(n_66),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_499),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_L g773 ( 
.A(n_604),
.B(n_60),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_610),
.B(n_1),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_499),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_570),
.B(n_78),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_480),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_571),
.B(n_59),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_589),
.B(n_1),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_533),
.B(n_2),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_500),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_533),
.B(n_559),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_559),
.B(n_4),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_500),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_501),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_501),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_621),
.B(n_4),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_588),
.B(n_84),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_505),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_592),
.B(n_86),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_505),
.B(n_79),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_506),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_614),
.B(n_583),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_506),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_517),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_517),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_629),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_629),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_673),
.B(n_547),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_744),
.B(n_521),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_636),
.Y(n_801)
);

BUFx8_ASAP7_75t_L g802 ( 
.A(n_630),
.Y(n_802)
);

AO22x2_ASAP7_75t_L g803 ( 
.A1(n_752),
.A2(n_490),
.B1(n_503),
.B2(n_520),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_716),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_716),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_636),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_728),
.A2(n_594),
.B1(n_490),
.B2(n_498),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_777),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_638),
.B(n_520),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_694),
.B(n_523),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_644),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_658),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_644),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_670),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_646),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_670),
.B(n_490),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_646),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_653),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_717),
.B(n_519),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_761),
.A2(n_490),
.B1(n_503),
.B2(n_523),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_741),
.A2(n_503),
.B1(n_624),
.B2(n_609),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_779),
.A2(n_609),
.B(n_558),
.C(n_590),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_696),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_653),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_779),
.A2(n_503),
.B1(n_14),
.B2(n_17),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_793),
.A2(n_552),
.B(n_590),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_637),
.B(n_587),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_746),
.B(n_769),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_674),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_SL g830 ( 
.A(n_656),
.B(n_616),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_718),
.B(n_549),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_689),
.Y(n_832)
);

INVx5_ASAP7_75t_L g833 ( 
.A(n_777),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_637),
.B(n_667),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_722),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_748),
.A2(n_549),
.B(n_548),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_777),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_760),
.A2(n_549),
.B1(n_548),
.B2(n_584),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_689),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_760),
.B(n_524),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_645),
.B(n_647),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_687),
.B(n_521),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_696),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_657),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_693),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_700),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_659),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_700),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_SL g849 ( 
.A1(n_774),
.A2(n_769),
.B1(n_719),
.B2(n_742),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_701),
.Y(n_850)
);

INVxp67_ASAP7_75t_SL g851 ( 
.A(n_777),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_697),
.B(n_552),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_793),
.A2(n_548),
.B1(n_563),
.B2(n_584),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_725),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_701),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_699),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_706),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_706),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_782),
.B(n_536),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_695),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_710),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_726),
.B(n_563),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_695),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_R g864 ( 
.A(n_766),
.B(n_112),
.Y(n_864)
);

OAI22xp33_ASAP7_75t_L g865 ( 
.A1(n_787),
.A2(n_526),
.B1(n_587),
.B2(n_536),
.Y(n_865)
);

AOI221xp5_ASAP7_75t_L g866 ( 
.A1(n_719),
.A2(n_524),
.B1(n_526),
.B2(n_547),
.C(n_583),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_774),
.A2(n_584),
.B1(n_563),
.B2(n_519),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_695),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_725),
.B(n_519),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_710),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_634),
.B(n_579),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_666),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_682),
.B(n_579),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_731),
.B(n_714),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_780),
.A2(n_616),
.B1(n_575),
.B2(n_480),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_698),
.A2(n_616),
.B(n_575),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_671),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_632),
.A2(n_616),
.B1(n_575),
.B2(n_480),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_680),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_739),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_667),
.B(n_575),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_713),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_686),
.Y(n_883)
);

AND2x6_ASAP7_75t_SL g884 ( 
.A(n_742),
.B(n_11),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_675),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_703),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_676),
.B(n_480),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_713),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_721),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_681),
.B(n_90),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_709),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_721),
.Y(n_892)
);

OR2x6_ASAP7_75t_L g893 ( 
.A(n_727),
.B(n_11),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_681),
.B(n_94),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_660),
.B(n_57),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_SL g896 ( 
.A1(n_669),
.A2(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_684),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_729),
.B(n_24),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_723),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_733),
.B(n_736),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_L g901 ( 
.A(n_631),
.B(n_98),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_780),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_723),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_730),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_684),
.B(n_25),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_737),
.B(n_35),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_753),
.B(n_35),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_775),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_753),
.B(n_691),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_695),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_633),
.B(n_108),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_775),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_784),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_662),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_668),
.B(n_38),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_783),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_730),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_678),
.B(n_41),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_732),
.B(n_715),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_656),
.B(n_116),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_633),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_754),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_747),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_643),
.B(n_45),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_SL g925 ( 
.A(n_679),
.B(n_46),
.C(n_48),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_627),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_641),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_740),
.B(n_692),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_747),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_669),
.B(n_53),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_759),
.A2(n_95),
.B(n_97),
.Y(n_931)
);

BUFx12f_ASAP7_75t_L g932 ( 
.A(n_635),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_784),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_785),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_715),
.B(n_101),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_724),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_785),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_679),
.B(n_113),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_677),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_786),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_672),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_654),
.A2(n_124),
.B(n_125),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_749),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_770),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_786),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_665),
.B(n_131),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_665),
.B(n_132),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_792),
.B(n_134),
.Y(n_948)
);

BUFx8_ASAP7_75t_L g949 ( 
.A(n_772),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_770),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_649),
.B(n_661),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_749),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_704),
.B(n_135),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_792),
.B(n_153),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_783),
.A2(n_773),
.B1(n_767),
.B2(n_794),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_707),
.B(n_708),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_661),
.A2(n_712),
.B1(n_743),
.B2(n_711),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_763),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_770),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_642),
.B(n_705),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_794),
.Y(n_961)
);

AND2x2_ASAP7_75t_SL g962 ( 
.A(n_771),
.B(n_790),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_750),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_750),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_781),
.B(n_796),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_745),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_789),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_795),
.A2(n_685),
.B1(n_755),
.B2(n_758),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_650),
.B(n_651),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_626),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_756),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_705),
.B(n_720),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_757),
.B(n_655),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_652),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_628),
.B(n_664),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_712),
.A2(n_751),
.B1(n_720),
.B2(n_690),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_683),
.B(n_688),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_764),
.B(n_768),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_626),
.A2(n_640),
.B1(n_735),
.B2(n_738),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_791),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_762),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_776),
.Y(n_982)
);

NOR2x1_ASAP7_75t_R g983 ( 
.A(n_640),
.B(n_788),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_765),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_849),
.A2(n_663),
.B(n_702),
.C(n_734),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_SL g986 ( 
.A1(n_896),
.A2(n_778),
.B1(n_639),
.B2(n_648),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_808),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_834),
.B(n_916),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_814),
.B(n_897),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_880),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_912),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_913),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_849),
.A2(n_828),
.B1(n_955),
.B2(n_916),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_814),
.B(n_897),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_856),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_844),
.B(n_941),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_799),
.B(n_914),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_799),
.B(n_914),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_863),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_L g1000 ( 
.A(n_812),
.B(n_872),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_938),
.A2(n_905),
.B(n_951),
.C(n_924),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_905),
.B(n_809),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_R g1003 ( 
.A(n_856),
.B(n_922),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_956),
.A2(n_873),
.B(n_833),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_SL g1005 ( 
.A1(n_825),
.A2(n_902),
.B1(n_932),
.B2(n_893),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_854),
.B(n_879),
.Y(n_1006)
);

NOR2xp67_ASAP7_75t_L g1007 ( 
.A(n_939),
.B(n_835),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_938),
.B(n_936),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_835),
.Y(n_1009)
);

INVx3_ASAP7_75t_SL g1010 ( 
.A(n_893),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_808),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_827),
.B(n_810),
.Y(n_1012)
);

INVx4_ASAP7_75t_L g1013 ( 
.A(n_863),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_SL g1014 ( 
.A(n_925),
.B(n_924),
.C(n_820),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_913),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_841),
.B(n_840),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_SL g1017 ( 
.A1(n_951),
.A2(n_955),
.B(n_919),
.C(n_969),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_SL g1018 ( 
.A1(n_890),
.A2(n_894),
.B(n_935),
.C(n_828),
.Y(n_1018)
);

CKINVDCx10_ASAP7_75t_R g1019 ( 
.A(n_893),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_930),
.B(n_874),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_879),
.B(n_883),
.Y(n_1021)
);

AND3x1_ASAP7_75t_L g1022 ( 
.A(n_816),
.B(n_902),
.C(n_805),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_925),
.A2(n_894),
.B(n_890),
.C(n_906),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_802),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_798),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_945),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_883),
.B(n_804),
.Y(n_1027)
);

BUFx4f_ASAP7_75t_L g1028 ( 
.A(n_946),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_982),
.B(n_981),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_833),
.A2(n_978),
.B(n_909),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_802),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_946),
.B(n_947),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_984),
.B(n_881),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_869),
.B(n_819),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_945),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_833),
.A2(n_973),
.B(n_830),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_970),
.A2(n_875),
.B1(n_821),
.B2(n_976),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_898),
.A2(n_928),
.B(n_847),
.C(n_877),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_984),
.B(n_926),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_804),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_R g1041 ( 
.A(n_921),
.B(n_830),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_957),
.A2(n_807),
.B(n_947),
.C(n_928),
.Y(n_1042)
);

OAI22x1_ASAP7_75t_L g1043 ( 
.A1(n_823),
.A2(n_843),
.B1(n_847),
.B2(n_958),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_823),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_SL g1045 ( 
.A1(n_980),
.A2(n_826),
.B(n_921),
.C(n_875),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_885),
.B(n_869),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_843),
.B(n_900),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_833),
.B(n_911),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_983),
.A2(n_876),
.B(n_977),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_977),
.A2(n_953),
.B(n_871),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_846),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_842),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_846),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_822),
.A2(n_887),
.B(n_918),
.C(n_915),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_R g1055 ( 
.A(n_863),
.B(n_868),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_851),
.A2(n_859),
.B(n_920),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_859),
.A2(n_920),
.B(n_980),
.Y(n_1057)
);

CKINVDCx16_ASAP7_75t_R g1058 ( 
.A(n_864),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_822),
.A2(n_907),
.B(n_895),
.C(n_891),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_864),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_962),
.A2(n_979),
.B(n_800),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_842),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_960),
.A2(n_886),
.B(n_974),
.C(n_972),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_911),
.B(n_960),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_808),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_926),
.B(n_927),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_863),
.B(n_868),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_927),
.B(n_974),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_868),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_808),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_803),
.B(n_967),
.Y(n_1071)
);

CKINVDCx6p67_ASAP7_75t_R g1072 ( 
.A(n_842),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_949),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_971),
.B(n_966),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_803),
.B(n_806),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_868),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_803),
.B(n_815),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_825),
.A2(n_901),
.B1(n_857),
.B2(n_850),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_SL g1079 ( 
.A(n_837),
.B(n_910),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_882),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_972),
.A2(n_975),
.B(n_895),
.C(n_852),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_819),
.B(n_831),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_865),
.A2(n_965),
.B(n_855),
.C(n_848),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_837),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_831),
.B(n_862),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_837),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_888),
.Y(n_1087)
);

NAND3xp33_ASAP7_75t_SL g1088 ( 
.A(n_942),
.B(n_931),
.C(n_968),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_862),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_SL g1090 ( 
.A(n_865),
.B(n_884),
.C(n_866),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_962),
.A2(n_954),
.B(n_948),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_889),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_892),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_860),
.B(n_910),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_949),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_968),
.B(n_797),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_SL g1097 ( 
.A(n_818),
.B(n_839),
.C(n_870),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_950),
.A2(n_837),
.B(n_860),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_950),
.A2(n_944),
.B(n_959),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_824),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_899),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_910),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_903),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_829),
.B(n_845),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_SL g1105 ( 
.A1(n_867),
.A2(n_838),
.B(n_853),
.C(n_878),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_944),
.A2(n_959),
.B(n_867),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_904),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_SL g1108 ( 
.A1(n_801),
.A2(n_811),
.B(n_813),
.C(n_817),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_944),
.A2(n_959),
.B1(n_963),
.B2(n_910),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_SL g1110 ( 
.A1(n_908),
.A2(n_934),
.B(n_961),
.C(n_940),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_944),
.A2(n_959),
.B(n_963),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_917),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_963),
.A2(n_836),
.B(n_832),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_963),
.A2(n_858),
.B(n_861),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_933),
.A2(n_937),
.B(n_929),
.C(n_923),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_943),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_952),
.A2(n_905),
.B(n_897),
.C(n_916),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_964),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_905),
.A2(n_897),
.B(n_916),
.C(n_834),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_956),
.A2(n_873),
.B(n_833),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_912),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_834),
.B(n_849),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_905),
.A2(n_897),
.B(n_916),
.C(n_834),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_814),
.B(n_897),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_834),
.B(n_916),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_834),
.B(n_916),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_834),
.B(n_916),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_956),
.A2(n_873),
.B(n_833),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_905),
.A2(n_897),
.B(n_916),
.C(n_834),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_863),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_856),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_956),
.A2(n_873),
.B(n_833),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_804),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_912),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1113),
.A2(n_1111),
.B(n_1049),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1001),
.A2(n_1023),
.B(n_1042),
.C(n_1002),
.Y(n_1136)
);

AOI221x1_ASAP7_75t_L g1137 ( 
.A1(n_993),
.A2(n_1088),
.B1(n_1037),
.B2(n_985),
.C(n_1061),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_SL g1138 ( 
.A1(n_1071),
.A2(n_1077),
.B(n_1075),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_SL g1139 ( 
.A1(n_1017),
.A2(n_1063),
.B(n_1032),
.C(n_1081),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_987),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1018),
.A2(n_1091),
.B(n_1017),
.Y(n_1141)
);

BUFx10_ASAP7_75t_L g1142 ( 
.A(n_1060),
.Y(n_1142)
);

BUFx10_ASAP7_75t_L g1143 ( 
.A(n_1031),
.Y(n_1143)
);

BUFx10_ASAP7_75t_L g1144 ( 
.A(n_1006),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1059),
.A2(n_1054),
.B(n_1050),
.Y(n_1145)
);

NOR2x1_ASAP7_75t_SL g1146 ( 
.A(n_1064),
.B(n_1020),
.Y(n_1146)
);

OAI22x1_ASAP7_75t_L g1147 ( 
.A1(n_1008),
.A2(n_1122),
.B1(n_1002),
.B2(n_1010),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1029),
.B(n_1021),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1057),
.A2(n_1099),
.B(n_1056),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1016),
.B(n_997),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_1021),
.B(n_1028),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1131),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1025),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_990),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1078),
.A2(n_1123),
.B(n_1119),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_988),
.B(n_1125),
.Y(n_1156)
);

OAI21xp33_ASAP7_75t_L g1157 ( 
.A1(n_1014),
.A2(n_1047),
.B(n_1124),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_998),
.B(n_1126),
.Y(n_1158)
);

OR2x6_ASAP7_75t_L g1159 ( 
.A(n_1048),
.B(n_1007),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1100),
.Y(n_1160)
);

AO21x1_ASAP7_75t_L g1161 ( 
.A1(n_1129),
.A2(n_1117),
.B(n_1038),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1034),
.B(n_1006),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1106),
.A2(n_1014),
.B(n_1012),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1004),
.A2(n_1128),
.B(n_1132),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1033),
.A2(n_1109),
.B(n_1083),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1003),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_1009),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1127),
.B(n_989),
.Y(n_1168)
);

NOR2xp67_ASAP7_75t_L g1169 ( 
.A(n_1000),
.B(n_1044),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1030),
.A2(n_1120),
.B(n_1045),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1114),
.A2(n_1098),
.B(n_1036),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_989),
.B(n_1124),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1027),
.B(n_1040),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1039),
.B(n_1074),
.Y(n_1174)
);

AO32x2_ASAP7_75t_L g1175 ( 
.A1(n_1005),
.A2(n_1022),
.A3(n_1076),
.B1(n_1013),
.B2(n_1090),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1034),
.B(n_1089),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1024),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1074),
.B(n_1118),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1094),
.A2(n_1115),
.B(n_1102),
.Y(n_1179)
);

AOI21xp33_ASAP7_75t_L g1180 ( 
.A1(n_1078),
.A2(n_1105),
.B(n_1028),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_995),
.B(n_1133),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1104),
.A2(n_1068),
.B(n_1067),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_1043),
.A2(n_1134),
.A3(n_1121),
.B(n_992),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1015),
.A2(n_1026),
.B(n_1035),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_SL g1185 ( 
.A(n_1058),
.B(n_1079),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1027),
.B(n_1003),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1051),
.A2(n_1053),
.A3(n_1066),
.B(n_1112),
.Y(n_1187)
);

NOR2x1_ASAP7_75t_SL g1188 ( 
.A(n_987),
.B(n_1086),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_1097),
.A2(n_1096),
.B(n_1116),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_999),
.A2(n_1069),
.B(n_1130),
.Y(n_1190)
);

NOR4xp25_ASAP7_75t_L g1191 ( 
.A(n_994),
.B(n_1110),
.C(n_996),
.D(n_1044),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1040),
.Y(n_1192)
);

AOI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1065),
.A2(n_1070),
.B(n_1084),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_987),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1105),
.A2(n_1090),
.B(n_1108),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1108),
.A2(n_1094),
.B(n_1046),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_987),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1082),
.A2(n_1085),
.B1(n_1062),
.B2(n_1052),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_999),
.A2(n_1069),
.B(n_1130),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1133),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1097),
.A2(n_986),
.B(n_1080),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_SL g1202 ( 
.A1(n_1011),
.A2(n_1086),
.B(n_1076),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1082),
.B(n_1085),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1087),
.A2(n_1107),
.A3(n_1103),
.B(n_1101),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1065),
.A2(n_1070),
.B(n_1084),
.Y(n_1205)
);

INVx3_ASAP7_75t_SL g1206 ( 
.A(n_1073),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_986),
.A2(n_1093),
.B(n_1092),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1072),
.B(n_1010),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1041),
.A2(n_1055),
.B(n_1013),
.Y(n_1209)
);

OAI21xp33_ASAP7_75t_L g1210 ( 
.A1(n_1095),
.A2(n_1041),
.B(n_1055),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1011),
.B(n_1086),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1011),
.A2(n_454),
.B1(n_1028),
.B2(n_1029),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1086),
.A2(n_1011),
.B(n_1019),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1113),
.A2(n_836),
.B(n_1111),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1002),
.B(n_670),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1001),
.A2(n_938),
.B(n_849),
.C(n_1023),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1002),
.B(n_834),
.Y(n_1217)
);

OR2x6_ASAP7_75t_L g1218 ( 
.A(n_1064),
.B(n_687),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1001),
.A2(n_1061),
.B(n_1042),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_990),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1018),
.A2(n_1091),
.B(n_1061),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1025),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1018),
.A2(n_1091),
.B(n_1061),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1018),
.A2(n_1091),
.B(n_1061),
.Y(n_1224)
);

OR2x6_ASAP7_75t_L g1225 ( 
.A(n_1064),
.B(n_687),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1001),
.A2(n_849),
.B1(n_1028),
.B2(n_1032),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1002),
.B(n_834),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1001),
.A2(n_849),
.B1(n_1028),
.B2(n_1032),
.Y(n_1228)
);

NAND3xp33_ASAP7_75t_L g1229 ( 
.A(n_1001),
.B(n_849),
.C(n_834),
.Y(n_1229)
);

OAI22x1_ASAP7_75t_L g1230 ( 
.A1(n_1008),
.A2(n_1032),
.B1(n_905),
.B2(n_1122),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1029),
.B(n_670),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1018),
.A2(n_1091),
.B(n_1061),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1001),
.A2(n_849),
.B1(n_1028),
.B2(n_1032),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1094),
.Y(n_1234)
);

O2A1O1Ixp5_ASAP7_75t_SL g1235 ( 
.A1(n_1122),
.A2(n_1008),
.B(n_993),
.C(n_1020),
.Y(n_1235)
);

AOI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1113),
.A2(n_1061),
.B(n_1020),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1025),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1001),
.A2(n_938),
.B(n_849),
.C(n_1023),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1002),
.B(n_834),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_995),
.B(n_562),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1131),
.Y(n_1241)
);

AOI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1113),
.A2(n_1061),
.B(n_1020),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1003),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1018),
.A2(n_1091),
.B(n_1061),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_991),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1002),
.B(n_670),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1008),
.A2(n_849),
.B1(n_670),
.B2(n_528),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1002),
.B(n_834),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1008),
.A2(n_849),
.B1(n_670),
.B2(n_528),
.Y(n_1249)
);

AO21x2_ASAP7_75t_L g1250 ( 
.A1(n_1001),
.A2(n_1088),
.B(n_1017),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1094),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1034),
.B(n_1006),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_SL g1253 ( 
.A1(n_1002),
.A2(n_905),
.B1(n_834),
.B2(n_670),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1001),
.A2(n_1061),
.B(n_1042),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1018),
.A2(n_1091),
.B(n_1061),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1018),
.A2(n_1091),
.B(n_1061),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_995),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1029),
.B(n_670),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1113),
.A2(n_836),
.B(n_1111),
.Y(n_1259)
);

NOR2x1_ASAP7_75t_R g1260 ( 
.A(n_1031),
.B(n_658),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1094),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1001),
.A2(n_1061),
.B(n_1042),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1025),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1018),
.A2(n_1091),
.B(n_1061),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_995),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1025),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1131),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1018),
.A2(n_1091),
.B(n_1061),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1008),
.A2(n_849),
.B1(n_670),
.B2(n_528),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1002),
.B(n_834),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1018),
.A2(n_1091),
.B(n_1061),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1034),
.B(n_1006),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1002),
.B(n_834),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1002),
.B(n_670),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1002),
.B(n_834),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1001),
.A2(n_1088),
.B(n_1017),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1131),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1001),
.A2(n_1061),
.B(n_1042),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1002),
.B(n_834),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1113),
.A2(n_836),
.B(n_1111),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1131),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1009),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1001),
.A2(n_938),
.B(n_849),
.C(n_1023),
.Y(n_1283)
);

OAI21xp33_ASAP7_75t_SL g1284 ( 
.A1(n_1180),
.A2(n_1235),
.B(n_1247),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1153),
.Y(n_1285)
);

BUFx5_ASAP7_75t_L g1286 ( 
.A(n_1160),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1200),
.Y(n_1287)
);

NAND2x1p5_ASAP7_75t_L g1288 ( 
.A(n_1151),
.B(n_1209),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1156),
.B(n_1217),
.Y(n_1289)
);

INVx3_ASAP7_75t_SL g1290 ( 
.A(n_1166),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1249),
.A2(n_1269),
.B1(n_1238),
.B2(n_1283),
.Y(n_1291)
);

AO21x2_ASAP7_75t_L g1292 ( 
.A1(n_1141),
.A2(n_1216),
.B(n_1170),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1137),
.A2(n_1264),
.A3(n_1221),
.B(n_1232),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1280),
.A2(n_1135),
.B(n_1149),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1227),
.B(n_1239),
.Y(n_1295)
);

BUFx12f_ASAP7_75t_L g1296 ( 
.A(n_1143),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1145),
.A2(n_1223),
.B(n_1255),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1257),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1215),
.B(n_1246),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1171),
.A2(n_1236),
.B(n_1242),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1164),
.A2(n_1244),
.B(n_1224),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1136),
.A2(n_1229),
.B(n_1231),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_1167),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1256),
.A2(n_1268),
.B(n_1271),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1145),
.A2(n_1196),
.B(n_1182),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1161),
.A2(n_1228),
.A3(n_1226),
.B(n_1233),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1229),
.A2(n_1278),
.B(n_1262),
.C(n_1254),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1226),
.A2(n_1228),
.A3(n_1233),
.B(n_1230),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1219),
.A2(n_1278),
.B(n_1262),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1178),
.A2(n_1274),
.B1(n_1275),
.B2(n_1279),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1195),
.A2(n_1163),
.B(n_1199),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1248),
.B(n_1270),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1273),
.A2(n_1253),
.B1(n_1172),
.B2(n_1150),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1222),
.Y(n_1314)
);

CKINVDCx6p67_ASAP7_75t_R g1315 ( 
.A(n_1206),
.Y(n_1315)
);

AOI221xp5_ASAP7_75t_L g1316 ( 
.A1(n_1155),
.A2(n_1258),
.B1(n_1157),
.B2(n_1180),
.C(n_1139),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1245),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1163),
.A2(n_1193),
.B(n_1207),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1234),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1250),
.A2(n_1276),
.B1(n_1147),
.B2(n_1148),
.Y(n_1320)
);

NAND3xp33_ASAP7_75t_L g1321 ( 
.A(n_1253),
.B(n_1155),
.C(n_1201),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1237),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1263),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1165),
.A2(n_1276),
.B(n_1250),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1201),
.A2(n_1158),
.B(n_1174),
.C(n_1207),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1168),
.A2(n_1266),
.B(n_1185),
.C(n_1210),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1243),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1203),
.B(n_1173),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1138),
.A2(n_1205),
.B(n_1190),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1187),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1177),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1187),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1251),
.B(n_1261),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1211),
.A2(n_1213),
.B(n_1179),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1187),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1143),
.Y(n_1336)
);

BUFx2_ASAP7_75t_SL g1337 ( 
.A(n_1169),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1189),
.A2(n_1197),
.B(n_1202),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1189),
.A2(n_1197),
.B(n_1251),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1185),
.A2(n_1198),
.B1(n_1212),
.B2(n_1218),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1218),
.A2(n_1225),
.B1(n_1186),
.B2(n_1241),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1208),
.A2(n_1146),
.B(n_1181),
.Y(n_1342)
);

INVx6_ASAP7_75t_L g1343 ( 
.A(n_1144),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1183),
.A2(n_1191),
.B(n_1188),
.Y(n_1344)
);

NOR2x1_ASAP7_75t_SL g1345 ( 
.A(n_1218),
.B(n_1225),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1282),
.Y(n_1346)
);

AO21x2_ASAP7_75t_L g1347 ( 
.A1(n_1191),
.A2(n_1183),
.B(n_1175),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1183),
.A2(n_1225),
.B(n_1204),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1204),
.A2(n_1175),
.B(n_1240),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1204),
.A2(n_1175),
.B(n_1159),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1159),
.A2(n_1140),
.B(n_1194),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1192),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1159),
.A2(n_1265),
.B1(n_1257),
.B2(n_1267),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1152),
.A2(n_1281),
.B1(n_1277),
.B2(n_1265),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1140),
.A2(n_1194),
.B(n_1144),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1142),
.Y(n_1356)
);

NAND3xp33_ASAP7_75t_L g1357 ( 
.A(n_1154),
.B(n_1220),
.C(n_1162),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1194),
.A2(n_1162),
.B(n_1252),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_SL g1359 ( 
.A1(n_1260),
.A2(n_1272),
.B(n_1176),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1272),
.A2(n_1259),
.B(n_1214),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1215),
.B(n_1246),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1152),
.Y(n_1362)
);

AO22x2_ASAP7_75t_L g1363 ( 
.A1(n_1226),
.A2(n_1233),
.B1(n_1228),
.B2(n_1137),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1216),
.A2(n_1001),
.B(n_1238),
.C(n_1283),
.Y(n_1364)
);

OR2x6_ASAP7_75t_L g1365 ( 
.A(n_1179),
.B(n_1218),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1153),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1234),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1216),
.A2(n_1001),
.B(n_1283),
.C(n_1238),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1229),
.A2(n_849),
.B1(n_1005),
.B2(n_896),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1153),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1156),
.B(n_1217),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_SL g1372 ( 
.A1(n_1146),
.A2(n_1161),
.B(n_1201),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1229),
.A2(n_849),
.B1(n_1005),
.B2(n_896),
.Y(n_1373)
);

AOI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1247),
.A2(n_849),
.B1(n_922),
.B2(n_331),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1200),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1247),
.A2(n_849),
.B1(n_1001),
.B2(n_1249),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1141),
.A2(n_1137),
.B(n_1221),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1184),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1167),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1257),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1153),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1234),
.B(n_1251),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1153),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1234),
.B(n_1251),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1229),
.A2(n_849),
.B1(n_1005),
.B2(n_896),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1184),
.Y(n_1386)
);

INVx6_ASAP7_75t_L g1387 ( 
.A(n_1144),
.Y(n_1387)
);

INVxp67_ASAP7_75t_SL g1388 ( 
.A(n_1200),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1152),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1234),
.B(n_1251),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1156),
.B(n_1217),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1216),
.A2(n_1001),
.B(n_834),
.Y(n_1392)
);

NAND2xp33_ASAP7_75t_SL g1393 ( 
.A(n_1226),
.B(n_1032),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1153),
.Y(n_1394)
);

NOR2xp67_ASAP7_75t_SL g1395 ( 
.A(n_1179),
.B(n_687),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1257),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1153),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1229),
.A2(n_849),
.B1(n_1005),
.B2(n_896),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1253),
.A2(n_1005),
.B1(n_896),
.B2(n_454),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1184),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1282),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1216),
.A2(n_1001),
.B(n_834),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1152),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1184),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1153),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1234),
.B(n_1251),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1153),
.Y(n_1407)
);

NOR3xp33_ASAP7_75t_L g1408 ( 
.A(n_1216),
.B(n_1001),
.C(n_849),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1399),
.A2(n_1398),
.B1(n_1385),
.B2(n_1373),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1399),
.A2(n_1398),
.B1(n_1385),
.B2(n_1373),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1287),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1299),
.B(n_1361),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1376),
.A2(n_1402),
.B(n_1392),
.C(n_1291),
.Y(n_1413)
);

O2A1O1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1368),
.A2(n_1408),
.B(n_1364),
.C(n_1307),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1297),
.A2(n_1304),
.B(n_1368),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1369),
.A2(n_1374),
.B1(n_1321),
.B2(n_1371),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1328),
.B(n_1352),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1408),
.A2(n_1393),
.B(n_1302),
.C(n_1316),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1289),
.B(n_1391),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1312),
.B(n_1295),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1285),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1369),
.A2(n_1341),
.B1(n_1354),
.B2(n_1312),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1310),
.B(n_1298),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1324),
.A2(n_1305),
.B(n_1301),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1313),
.B(n_1325),
.Y(n_1425)
);

A2O1A1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1393),
.A2(n_1284),
.B(n_1326),
.C(n_1395),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1287),
.B(n_1388),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1325),
.B(n_1380),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1326),
.A2(n_1372),
.B(n_1340),
.C(n_1353),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1396),
.B(n_1388),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1341),
.A2(n_1354),
.B1(n_1357),
.B2(n_1363),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1303),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1382),
.B(n_1384),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1390),
.B(n_1406),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1340),
.A2(n_1346),
.B1(n_1401),
.B2(n_1331),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1375),
.B(n_1362),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1390),
.B(n_1406),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1363),
.A2(n_1337),
.B1(n_1320),
.B2(n_1403),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1375),
.B(n_1389),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1318),
.A2(n_1300),
.B(n_1344),
.Y(n_1440)
);

BUFx12f_ASAP7_75t_L g1441 ( 
.A(n_1336),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1365),
.A2(n_1345),
.B(n_1377),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1317),
.B(n_1358),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1317),
.B(n_1342),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1314),
.A2(n_1407),
.B(n_1405),
.C(n_1322),
.Y(n_1445)
);

AOI21x1_ASAP7_75t_SL g1446 ( 
.A1(n_1363),
.A2(n_1306),
.B(n_1292),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1323),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1366),
.B(n_1370),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1381),
.A2(n_1394),
.B(n_1383),
.C(n_1397),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1379),
.B(n_1367),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1379),
.B(n_1367),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1300),
.A2(n_1311),
.B(n_1309),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1319),
.B(n_1308),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1319),
.B(n_1308),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1349),
.B(n_1350),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1346),
.B(n_1303),
.Y(n_1456)
);

AOI211xp5_ASAP7_75t_L g1457 ( 
.A1(n_1290),
.A2(n_1334),
.B(n_1336),
.C(n_1327),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1356),
.A2(n_1343),
.B1(n_1387),
.B2(n_1288),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1356),
.A2(n_1343),
.B1(n_1387),
.B2(n_1288),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1387),
.A2(n_1290),
.B1(n_1331),
.B2(n_1333),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1338),
.A2(n_1351),
.B(n_1348),
.C(n_1339),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1355),
.B(n_1286),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1348),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1327),
.A2(n_1329),
.B(n_1347),
.Y(n_1464)
);

O2A1O1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1359),
.A2(n_1335),
.B(n_1332),
.C(n_1330),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1315),
.A2(n_1296),
.B1(n_1329),
.B2(n_1404),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1286),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1286),
.B(n_1293),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1347),
.B(n_1293),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1296),
.A2(n_1378),
.B1(n_1400),
.B2(n_1386),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1293),
.B(n_1360),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1294),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1297),
.A2(n_1238),
.B(n_1216),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1289),
.B(n_1371),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_SL g1475 ( 
.A1(n_1368),
.A2(n_1001),
.B(n_1216),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1364),
.A2(n_1001),
.B(n_849),
.C(n_1216),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1362),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1328),
.B(n_1352),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1287),
.Y(n_1479)
);

OAI31xp33_ASAP7_75t_L g1480 ( 
.A1(n_1376),
.A2(n_1001),
.A3(n_1238),
.B(n_1216),
.Y(n_1480)
);

BUFx4f_ASAP7_75t_SL g1481 ( 
.A(n_1303),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1289),
.B(n_1371),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1469),
.B(n_1471),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1420),
.B(n_1479),
.Y(n_1484)
);

OR2x6_ASAP7_75t_L g1485 ( 
.A(n_1415),
.B(n_1442),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1455),
.B(n_1468),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1453),
.B(n_1454),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1452),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1432),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1472),
.B(n_1461),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1447),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1409),
.A2(n_1410),
.B1(n_1416),
.B2(n_1480),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1462),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1463),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1444),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1422),
.A2(n_1473),
.B1(n_1425),
.B2(n_1435),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1411),
.B(n_1427),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1411),
.B(n_1421),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1440),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1467),
.B(n_1443),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1470),
.Y(n_1501)
);

INVxp67_ASAP7_75t_SL g1502 ( 
.A(n_1445),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1430),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1424),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1445),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1449),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1473),
.B(n_1418),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1475),
.B(n_1423),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1466),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1448),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1449),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1464),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1428),
.B(n_1438),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1465),
.Y(n_1514)
);

AO31x2_ASAP7_75t_L g1515 ( 
.A1(n_1476),
.A2(n_1426),
.A3(n_1446),
.B(n_1431),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1494),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1492),
.A2(n_1413),
.B1(n_1482),
.B2(n_1419),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1483),
.B(n_1465),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_SL g1519 ( 
.A(n_1507),
.B(n_1413),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1488),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1483),
.B(n_1414),
.Y(n_1521)
);

INVxp67_ASAP7_75t_SL g1522 ( 
.A(n_1502),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1483),
.B(n_1414),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1490),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1503),
.B(n_1417),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1495),
.B(n_1437),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1499),
.B(n_1495),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1495),
.B(n_1433),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1503),
.B(n_1478),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1490),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1492),
.A2(n_1507),
.B1(n_1496),
.B2(n_1513),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1499),
.B(n_1439),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1499),
.B(n_1436),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1495),
.B(n_1434),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1504),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1486),
.B(n_1412),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1531),
.A2(n_1496),
.B1(n_1507),
.B2(n_1513),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1519),
.A2(n_1508),
.B1(n_1513),
.B2(n_1509),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1524),
.B(n_1530),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_R g1540 ( 
.A(n_1519),
.B(n_1489),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1536),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1516),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1532),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1519),
.B(n_1501),
.C(n_1508),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1531),
.A2(n_1508),
.B1(n_1509),
.B2(n_1485),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1520),
.Y(n_1546)
);

NAND2xp33_ASAP7_75t_SL g1547 ( 
.A(n_1517),
.B(n_1509),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1517),
.A2(n_1429),
.B1(n_1457),
.B2(n_1485),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1532),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1536),
.B(n_1526),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1526),
.B(n_1493),
.Y(n_1551)
);

AOI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1522),
.A2(n_1502),
.B1(n_1429),
.B2(n_1491),
.C(n_1484),
.Y(n_1552)
);

OR2x6_ASAP7_75t_L g1553 ( 
.A(n_1524),
.B(n_1485),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1516),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_L g1555 ( 
.A(n_1524),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1532),
.Y(n_1556)
);

OAI31xp33_ASAP7_75t_L g1557 ( 
.A1(n_1522),
.A2(n_1460),
.A3(n_1458),
.B(n_1459),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1521),
.A2(n_1512),
.B(n_1501),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1526),
.B(n_1493),
.Y(n_1559)
);

OAI31xp33_ASAP7_75t_L g1560 ( 
.A1(n_1521),
.A2(n_1512),
.A3(n_1505),
.B(n_1506),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1521),
.A2(n_1485),
.B1(n_1511),
.B2(n_1505),
.Y(n_1561)
);

NAND4xp25_ASAP7_75t_L g1562 ( 
.A(n_1533),
.B(n_1474),
.C(n_1484),
.D(n_1506),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1533),
.B(n_1511),
.C(n_1506),
.Y(n_1563)
);

INVx5_ASAP7_75t_L g1564 ( 
.A(n_1535),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1528),
.B(n_1534),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_SL g1566 ( 
.A1(n_1524),
.A2(n_1489),
.B1(n_1481),
.B2(n_1441),
.Y(n_1566)
);

OAI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1525),
.A2(n_1485),
.B1(n_1451),
.B2(n_1450),
.C(n_1491),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1525),
.B(n_1477),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1523),
.A2(n_1510),
.B1(n_1498),
.B2(n_1497),
.C(n_1487),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1529),
.Y(n_1570)
);

A2O1A1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1523),
.A2(n_1512),
.B(n_1514),
.C(n_1515),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1530),
.B(n_1500),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1564),
.B(n_1530),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1546),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1569),
.B(n_1533),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1549),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1556),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1540),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1542),
.Y(n_1579)
);

INVx4_ASAP7_75t_SL g1580 ( 
.A(n_1566),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1554),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1564),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1543),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1563),
.B(n_1527),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1564),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1562),
.B(n_1533),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1543),
.Y(n_1587)
);

INVxp67_ASAP7_75t_SL g1588 ( 
.A(n_1555),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1564),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1564),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1565),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1548),
.A2(n_1512),
.B(n_1518),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1555),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1555),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1555),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1553),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1553),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1550),
.B(n_1551),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1539),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1573),
.B(n_1539),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1578),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1574),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1599),
.B(n_1539),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1578),
.B(n_1570),
.Y(n_1604)
);

AND2x2_ASAP7_75t_SL g1605 ( 
.A(n_1590),
.B(n_1538),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1579),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1586),
.B(n_1570),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1574),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1579),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1586),
.B(n_1552),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1573),
.B(n_1553),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1579),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1596),
.A2(n_1547),
.B1(n_1537),
.B2(n_1544),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1573),
.B(n_1553),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1581),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1573),
.B(n_1591),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1583),
.Y(n_1617)
);

OAI31xp33_ASAP7_75t_SL g1618 ( 
.A1(n_1588),
.A2(n_1567),
.A3(n_1547),
.B(n_1568),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1573),
.B(n_1572),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1573),
.B(n_1572),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1581),
.Y(n_1621)
);

NOR2xp67_ASAP7_75t_L g1622 ( 
.A(n_1585),
.B(n_1558),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1575),
.B(n_1560),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1574),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1581),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1580),
.B(n_1557),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1598),
.B(n_1559),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1583),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1575),
.B(n_1518),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1588),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1592),
.B(n_1571),
.C(n_1545),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1577),
.B(n_1518),
.Y(n_1632)
);

INVx2_ASAP7_75t_SL g1633 ( 
.A(n_1590),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1576),
.A2(n_1518),
.B1(n_1541),
.B2(n_1571),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1622),
.B(n_1580),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1617),
.B(n_1584),
.Y(n_1636)
);

INVxp67_ASAP7_75t_SL g1637 ( 
.A(n_1622),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1601),
.B(n_1592),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1601),
.B(n_1587),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1606),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1617),
.B(n_1584),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1633),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1600),
.B(n_1603),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1616),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1606),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1609),
.Y(n_1646)
);

NAND2x1p5_ASAP7_75t_L g1647 ( 
.A(n_1633),
.B(n_1590),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1609),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1616),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1610),
.B(n_1587),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1612),
.Y(n_1651)
);

AOI21xp33_ASAP7_75t_L g1652 ( 
.A1(n_1605),
.A2(n_1585),
.B(n_1590),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1605),
.A2(n_1580),
.B1(n_1597),
.B2(n_1596),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1610),
.B(n_1587),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1600),
.B(n_1593),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1600),
.B(n_1603),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1627),
.B(n_1593),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1612),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1615),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1615),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1621),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1623),
.B(n_1598),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1604),
.B(n_1597),
.Y(n_1663)
);

OAI21xp33_ASAP7_75t_L g1664 ( 
.A1(n_1618),
.A2(n_1596),
.B(n_1561),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1616),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1633),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1628),
.B(n_1632),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1626),
.B(n_1597),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1602),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1628),
.B(n_1580),
.Y(n_1670)
);

CKINVDCx14_ASAP7_75t_R g1671 ( 
.A(n_1663),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1664),
.A2(n_1605),
.B1(n_1631),
.B2(n_1634),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1640),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1650),
.B(n_1618),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1640),
.Y(n_1675)
);

INVx4_ASAP7_75t_L g1676 ( 
.A(n_1670),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1637),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1668),
.B(n_1607),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1645),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1642),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1654),
.B(n_1607),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1647),
.Y(n_1683)
);

AOI222xp33_ASAP7_75t_L g1684 ( 
.A1(n_1638),
.A2(n_1623),
.B1(n_1631),
.B2(n_1613),
.C1(n_1629),
.C2(n_1580),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1636),
.B(n_1630),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1642),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1645),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1639),
.B(n_1629),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1646),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1662),
.B(n_1670),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1646),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1647),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1670),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1648),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1647),
.A2(n_1582),
.B(n_1589),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1677),
.B(n_1643),
.Y(n_1698)
);

AOI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1686),
.A2(n_1666),
.B(n_1641),
.Y(n_1699)
);

NOR2x1_ASAP7_75t_L g1700 ( 
.A(n_1676),
.B(n_1666),
.Y(n_1700)
);

CKINVDCx14_ASAP7_75t_R g1701 ( 
.A(n_1671),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1672),
.A2(n_1653),
.B(n_1652),
.Y(n_1702)
);

INVx4_ASAP7_75t_L g1703 ( 
.A(n_1676),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1676),
.Y(n_1704)
);

INVxp67_ASAP7_75t_SL g1705 ( 
.A(n_1685),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1673),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1674),
.A2(n_1634),
.B1(n_1636),
.B2(n_1641),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1673),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1681),
.A2(n_1630),
.B1(n_1667),
.B2(n_1643),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1695),
.Y(n_1710)
);

NAND2xp33_ASAP7_75t_R g1711 ( 
.A(n_1685),
.B(n_1667),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1684),
.B(n_1656),
.Y(n_1712)
);

NAND2x1_ASAP7_75t_L g1713 ( 
.A(n_1676),
.B(n_1656),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1678),
.A2(n_1580),
.B1(n_1655),
.B2(n_1657),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1690),
.B(n_1655),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1675),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1707),
.A2(n_1682),
.B1(n_1694),
.B2(n_1691),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1701),
.B(n_1682),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1705),
.B(n_1691),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1710),
.B(n_1694),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1700),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1698),
.B(n_1688),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1702),
.A2(n_1680),
.B1(n_1597),
.B2(n_1596),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1704),
.B(n_1680),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1706),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1708),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1723),
.A2(n_1702),
.B1(n_1709),
.B2(n_1712),
.C(n_1715),
.Y(n_1727)
);

OAI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1717),
.A2(n_1711),
.B1(n_1714),
.B2(n_1713),
.C(n_1703),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1718),
.B(n_1703),
.Y(n_1729)
);

AO22x1_ASAP7_75t_L g1730 ( 
.A1(n_1721),
.A2(n_1680),
.B1(n_1693),
.B2(n_1683),
.Y(n_1730)
);

OAI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1719),
.A2(n_1699),
.B1(n_1716),
.B2(n_1696),
.C(n_1683),
.Y(n_1731)
);

NAND3xp33_ASAP7_75t_SL g1732 ( 
.A(n_1720),
.B(n_1722),
.C(n_1724),
.Y(n_1732)
);

OAI211xp5_ASAP7_75t_SL g1733 ( 
.A1(n_1725),
.A2(n_1696),
.B(n_1679),
.C(n_1692),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1726),
.B(n_1580),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1718),
.A2(n_1693),
.B(n_1697),
.Y(n_1735)
);

XNOR2xp5_ASAP7_75t_L g1736 ( 
.A(n_1727),
.B(n_1693),
.Y(n_1736)
);

XNOR2xp5_ASAP7_75t_L g1737 ( 
.A(n_1728),
.B(n_1456),
.Y(n_1737)
);

O2A1O1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1731),
.A2(n_1732),
.B(n_1734),
.C(n_1733),
.Y(n_1738)
);

AOI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1730),
.A2(n_1675),
.B1(n_1692),
.B2(n_1689),
.C(n_1687),
.Y(n_1739)
);

AOI322xp5_ASAP7_75t_L g1740 ( 
.A1(n_1729),
.A2(n_1689),
.A3(n_1687),
.B1(n_1679),
.B2(n_1644),
.C1(n_1649),
.C2(n_1665),
.Y(n_1740)
);

NOR2xp67_ASAP7_75t_L g1741 ( 
.A(n_1736),
.B(n_1735),
.Y(n_1741)
);

NOR3xp33_ASAP7_75t_L g1742 ( 
.A(n_1738),
.B(n_1697),
.C(n_1649),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1737),
.B(n_1657),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1739),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1740),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1736),
.B(n_1644),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1743),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1741),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1746),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1744),
.Y(n_1750)
);

OAI221xp5_ASAP7_75t_SL g1751 ( 
.A1(n_1745),
.A2(n_1665),
.B1(n_1659),
.B2(n_1661),
.C(n_1660),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1748),
.Y(n_1752)
);

NAND4xp75_ASAP7_75t_L g1753 ( 
.A(n_1749),
.B(n_1742),
.C(n_1658),
.D(n_1651),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1747),
.B(n_1620),
.Y(n_1754)
);

NOR4xp25_ASAP7_75t_L g1755 ( 
.A(n_1754),
.B(n_1751),
.C(n_1750),
.D(n_1669),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1755),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1756),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1756),
.B(n_1752),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1757),
.A2(n_1751),
.B(n_1753),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1758),
.A2(n_1669),
.B1(n_1621),
.B2(n_1625),
.Y(n_1760)
);

XNOR2xp5_ASAP7_75t_L g1761 ( 
.A(n_1759),
.B(n_1758),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1760),
.A2(n_1590),
.B1(n_1594),
.B2(n_1589),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1761),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1762),
.A2(n_1590),
.B1(n_1594),
.B2(n_1589),
.Y(n_1764)
);

NOR4xp25_ASAP7_75t_L g1765 ( 
.A(n_1763),
.B(n_1625),
.C(n_1608),
.D(n_1602),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1764),
.B(n_1608),
.Y(n_1766)
);

OAI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1766),
.A2(n_1624),
.B1(n_1608),
.B2(n_1602),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1767),
.A2(n_1611),
.B1(n_1614),
.B2(n_1595),
.Y(n_1768)
);

AOI211xp5_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1590),
.B(n_1589),
.C(n_1624),
.Y(n_1769)
);


endmodule