module fake_jpeg_275_n_689 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_689);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_689;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_441;
wire n_161;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_61),
.Y(n_159)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_64),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_67),
.Y(n_202)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_73),
.Y(n_214)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_22),
.B(n_15),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_87),
.Y(n_138)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g189 ( 
.A(n_76),
.Y(n_189)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_79),
.Y(n_167)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_22),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_81),
.B(n_83),
.Y(n_197)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_1),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_84),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_23),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_30),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_88),
.B(n_91),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_89),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_28),
.Y(n_90)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_38),
.B(n_40),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_92),
.Y(n_196)
);

BUFx4f_ASAP7_75t_SL g93 ( 
.A(n_28),
.Y(n_93)
);

BUFx24_ASAP7_75t_L g178 ( 
.A(n_93),
.Y(n_178)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_95),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_96),
.B(n_100),
.Y(n_171)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_37),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_23),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_38),
.B(n_2),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_101),
.B(n_21),
.Y(n_154)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_51),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_107),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_106),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_36),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_111),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_51),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_112),
.B(n_118),
.Y(n_182)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_29),
.Y(n_113)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_29),
.Y(n_115)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_116),
.Y(n_219)
);

BUFx4f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_117),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_47),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_119),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_40),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_125),
.B(n_126),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_35),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_34),
.Y(n_127)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_127),
.Y(n_225)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_34),
.Y(n_128)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_48),
.Y(n_130)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_64),
.B(n_48),
.C(n_39),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_134),
.B(n_189),
.C(n_156),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_135),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_93),
.B(n_42),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_142),
.B(n_187),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_58),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_151),
.B(n_72),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_154),
.B(n_168),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_84),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_157),
.B(n_170),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_117),
.B(n_21),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_89),
.Y(n_170)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_92),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g235 ( 
.A(n_176),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_104),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_177),
.B(n_181),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_111),
.Y(n_181)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_73),
.Y(n_184)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_184),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_119),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_185),
.B(n_206),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_73),
.A2(n_26),
.B1(n_58),
.B2(n_42),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g301 ( 
.A1(n_186),
.A2(n_205),
.B1(n_9),
.B2(n_10),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_93),
.B(n_50),
.Y(n_187)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_188),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_77),
.B(n_50),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_193),
.B(n_201),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_71),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_195),
.Y(n_270)
);

BUFx16f_ASAP7_75t_L g199 ( 
.A(n_90),
.Y(n_199)
);

BUFx8_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_94),
.B(n_43),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_110),
.B(n_43),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_204),
.B(n_211),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_122),
.A2(n_26),
.B1(n_41),
.B2(n_25),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_120),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_210),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_106),
.B(n_41),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_98),
.B(n_25),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_216),
.B(n_221),
.Y(n_291)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_70),
.B(n_24),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_61),
.Y(n_222)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_132),
.Y(n_226)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_226),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_131),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_227),
.B(n_252),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_140),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_228),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_218),
.A2(n_129),
.B1(n_123),
.B2(n_103),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_229),
.A2(n_251),
.B1(n_262),
.B2(n_271),
.Y(n_321)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_140),
.Y(n_230)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_230),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx3_ASAP7_75t_SL g325 ( 
.A(n_231),
.Y(n_325)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_232),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_138),
.A2(n_63),
.B1(n_65),
.B2(n_69),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_233),
.A2(n_283),
.B1(n_289),
.B2(n_292),
.Y(n_310)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_236),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_238),
.Y(n_363)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_165),
.Y(n_239)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_239),
.Y(n_337)
);

NAND2x1_ASAP7_75t_SL g331 ( 
.A(n_242),
.B(n_257),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_190),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_243),
.B(n_268),
.Y(n_335)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_244),
.Y(n_342)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_159),
.Y(n_246)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_246),
.Y(n_329)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_248),
.Y(n_361)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_179),
.Y(n_249)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_249),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_218),
.A2(n_99),
.B1(n_95),
.B2(n_86),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_24),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_143),
.Y(n_253)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_139),
.Y(n_254)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_254),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_151),
.B(n_85),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_147),
.Y(n_258)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_147),
.Y(n_260)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_260),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_261),
.B(n_180),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_171),
.A2(n_202),
.B1(n_189),
.B2(n_163),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_173),
.B(n_207),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_264),
.B(n_265),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_172),
.B(n_2),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_205),
.A2(n_54),
.B(n_55),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_266),
.A2(n_286),
.B(n_271),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_182),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_203),
.Y(n_269)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_202),
.A2(n_55),
.B1(n_36),
.B2(n_4),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_133),
.B(n_2),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_272),
.B(n_273),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_167),
.B(n_3),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_156),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_274),
.B(n_287),
.Y(n_350)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_194),
.Y(n_275)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_203),
.Y(n_276)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_276),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_192),
.Y(n_277)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_277),
.Y(n_369)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_139),
.Y(n_278)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_192),
.Y(n_279)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_279),
.Y(n_318)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_158),
.Y(n_282)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_208),
.A2(n_225),
.B1(n_212),
.B2(n_150),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_155),
.Y(n_284)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_178),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_136),
.B(n_7),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_178),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_288),
.B(n_293),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_137),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_183),
.Y(n_290)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_290),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_186),
.A2(n_149),
.B1(n_146),
.B2(n_145),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_183),
.B(n_8),
.Y(n_293)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_143),
.Y(n_294)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_163),
.B(n_8),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_302),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_153),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_296),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_196),
.Y(n_297)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_141),
.B(n_8),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_298),
.Y(n_354)
);

BUFx12_ASAP7_75t_L g299 ( 
.A(n_178),
.Y(n_299)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_175),
.Y(n_300)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_301),
.A2(n_166),
.B1(n_169),
.B2(n_219),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_200),
.B(n_9),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_180),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_303),
.A2(n_196),
.B1(n_215),
.B2(n_217),
.Y(n_315)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_200),
.Y(n_304)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_209),
.Y(n_305)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_141),
.B(n_11),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_12),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_152),
.B(n_14),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_184),
.C(n_166),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_308),
.B(n_322),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_315),
.A2(n_310),
.B1(n_359),
.B2(n_369),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_316),
.B(n_12),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_237),
.C(n_227),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_291),
.A2(n_266),
.B1(n_245),
.B2(n_298),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_323),
.A2(n_334),
.B1(n_360),
.B2(n_235),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_326),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_152),
.C(n_169),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_332),
.B(n_344),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_252),
.A2(n_176),
.B1(n_191),
.B2(n_164),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_L g370 ( 
.A1(n_341),
.A2(n_251),
.B1(n_229),
.B2(n_267),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_242),
.B(n_158),
.C(n_223),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_345),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_257),
.B(n_219),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_346),
.B(n_362),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_267),
.A2(n_166),
.B1(n_188),
.B2(n_144),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_347),
.A2(n_270),
.B1(n_263),
.B2(n_241),
.Y(n_389)
);

O2A1O1Ixp33_ASAP7_75t_SL g349 ( 
.A1(n_301),
.A2(n_144),
.B(n_148),
.C(n_210),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_349),
.A2(n_247),
.B(n_270),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_234),
.B(n_164),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_286),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_280),
.B(n_223),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_355),
.B(n_303),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_283),
.A2(n_191),
.B1(n_174),
.B2(n_160),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_256),
.B(n_160),
.C(n_174),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_301),
.B(n_209),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_365),
.A2(n_367),
.B(n_263),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_262),
.A2(n_148),
.B(n_210),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_370),
.B(n_374),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_371),
.B(n_376),
.Y(n_420)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_363),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_372),
.Y(n_452)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_230),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_307),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_377),
.B(n_365),
.Y(n_437)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_329),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_325),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_379),
.Y(n_451)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_363),
.Y(n_380)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_380),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_308),
.B(n_255),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_381),
.B(n_396),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_336),
.B(n_240),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_383),
.B(n_392),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_326),
.B(n_282),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_384),
.A2(n_365),
.B(n_321),
.Y(n_434)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_319),
.Y(n_385)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_385),
.Y(n_445)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_386),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_365),
.A2(n_253),
.B1(n_294),
.B2(n_269),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_387),
.A2(n_389),
.B(n_399),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_388),
.A2(n_397),
.B1(n_402),
.B2(n_412),
.Y(n_439)
);

INVx13_ASAP7_75t_L g390 ( 
.A(n_357),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_390),
.Y(n_426)
);

OAI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_391),
.A2(n_314),
.B1(n_369),
.B2(n_318),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_351),
.B(n_232),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_339),
.B(n_322),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_393),
.B(n_403),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_367),
.A2(n_250),
.B(n_285),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_394),
.A2(n_416),
.B(n_241),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_324),
.B(n_278),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_345),
.A2(n_289),
.B1(n_159),
.B2(n_217),
.Y(n_397)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_400),
.Y(n_450)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_333),
.Y(n_401)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_401),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_315),
.A2(n_215),
.B1(n_246),
.B2(n_235),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_364),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_332),
.B(n_276),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_407),
.Y(n_432)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_405),
.Y(n_459)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_406),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_350),
.B(n_260),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_410),
.Y(n_435)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_352),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_414),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_328),
.A2(n_277),
.B1(n_297),
.B2(n_279),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_356),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_312),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_309),
.Y(n_444)
);

O2A1O1Ixp33_ASAP7_75t_L g416 ( 
.A1(n_349),
.A2(n_241),
.B(n_305),
.C(n_299),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_331),
.B(n_346),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_417),
.A2(n_309),
.B(n_364),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_313),
.B(n_258),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_325),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_395),
.A2(n_377),
.B1(n_398),
.B2(n_384),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_419),
.A2(n_442),
.B1(n_454),
.B2(n_397),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_388),
.A2(n_362),
.B1(n_328),
.B2(n_344),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_425),
.A2(n_430),
.B1(n_376),
.B2(n_381),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_313),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_429),
.B(n_430),
.C(n_408),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_331),
.C(n_353),
.Y(n_430)
);

AO21x1_ASAP7_75t_L g460 ( 
.A1(n_434),
.A2(n_458),
.B(n_399),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_437),
.B(n_330),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_396),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_440),
.B(n_443),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_441),
.A2(n_449),
.B(n_394),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_395),
.A2(n_354),
.B1(n_316),
.B2(n_360),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_406),
.Y(n_443)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_446),
.A2(n_412),
.B1(n_402),
.B2(n_401),
.Y(n_471)
);

FAx1_ASAP7_75t_SL g448 ( 
.A(n_382),
.B(n_366),
.CI(n_311),
.CON(n_448),
.SN(n_448)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_448),
.B(n_455),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_384),
.A2(n_340),
.B(n_320),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_398),
.A2(n_338),
.B1(n_153),
.B2(n_161),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_385),
.B(n_348),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_403),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_460),
.A2(n_463),
.B(n_469),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_440),
.B(n_418),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_461),
.B(n_470),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_387),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_462),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_428),
.A2(n_374),
.B(n_416),
.Y(n_463)
);

BUFx24_ASAP7_75t_SL g465 ( 
.A(n_423),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_465),
.B(n_483),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_423),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_466),
.B(n_474),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_439),
.A2(n_391),
.B1(n_398),
.B2(n_408),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_467),
.A2(n_486),
.B1(n_487),
.B2(n_492),
.Y(n_503)
);

INVx13_ASAP7_75t_L g468 ( 
.A(n_453),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_468),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_429),
.B(n_358),
.Y(n_470)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_471),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_472),
.B(n_495),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_428),
.A2(n_417),
.B(n_408),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_473),
.A2(n_458),
.B(n_424),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_438),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_475),
.B(n_493),
.Y(n_508)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_438),
.Y(n_476)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_476),
.Y(n_499)
);

INVx13_ASAP7_75t_L g478 ( 
.A(n_453),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_478),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_434),
.B(n_417),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_479),
.B(n_436),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_447),
.B(n_371),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_481),
.B(n_485),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_482),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_444),
.Y(n_484)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_484),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_433),
.B(n_414),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_439),
.A2(n_400),
.B1(n_411),
.B2(n_405),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_428),
.A2(n_378),
.B1(n_373),
.B2(n_372),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_447),
.B(n_409),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_488),
.B(n_489),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_457),
.B(n_415),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_490),
.B(n_419),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_435),
.B(n_410),
.Y(n_491)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_491),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_431),
.A2(n_380),
.B1(n_379),
.B2(n_343),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_431),
.B(n_368),
.C(n_337),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_435),
.B(n_432),
.Y(n_494)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_494),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_448),
.B(n_386),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_SL g496 ( 
.A(n_449),
.B(n_379),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_496),
.A2(n_426),
.B(n_456),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_420),
.A2(n_343),
.B1(n_368),
.B2(n_337),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_497),
.A2(n_450),
.B1(n_445),
.B2(n_421),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_SL g550 ( 
.A(n_501),
.B(n_473),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_482),
.A2(n_425),
.B1(n_420),
.B2(n_432),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_505),
.A2(n_530),
.B1(n_452),
.B2(n_478),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_474),
.B(n_454),
.Y(n_509)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_509),
.Y(n_555)
);

NOR3xp33_ASAP7_75t_L g512 ( 
.A(n_480),
.B(n_424),
.C(n_448),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_512),
.B(n_529),
.Y(n_540)
);

AO21x1_ASAP7_75t_L g559 ( 
.A1(n_514),
.A2(n_531),
.B(n_478),
.Y(n_559)
);

NOR4xp25_ASAP7_75t_L g517 ( 
.A(n_483),
.B(n_448),
.C(n_437),
.D(n_450),
.Y(n_517)
);

NOR3xp33_ASAP7_75t_SL g563 ( 
.A(n_517),
.B(n_534),
.C(n_468),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_464),
.B(n_456),
.Y(n_518)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_518),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_480),
.B(n_442),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_519),
.B(n_528),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_464),
.B(n_459),
.Y(n_520)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_520),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_523),
.A2(n_531),
.B(n_500),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_463),
.A2(n_443),
.B1(n_436),
.B2(n_459),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_524),
.A2(n_486),
.B1(n_487),
.B2(n_489),
.Y(n_539)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_477),
.Y(n_525)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_525),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_494),
.B(n_455),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_472),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_469),
.A2(n_426),
.B(n_421),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_477),
.Y(n_532)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_532),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_533),
.B(n_462),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_488),
.B(n_445),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_527),
.A2(n_461),
.B1(n_481),
.B2(n_476),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_535),
.A2(n_546),
.B1(n_554),
.B2(n_557),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_510),
.A2(n_462),
.B(n_460),
.Y(n_536)
);

AO21x1_ASAP7_75t_L g579 ( 
.A1(n_536),
.A2(n_543),
.B(n_548),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_513),
.B(n_484),
.Y(n_537)
);

CKINVDCx14_ASAP7_75t_R g588 ( 
.A(n_537),
.Y(n_588)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_538),
.Y(n_569)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_539),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_508),
.B(n_475),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_541),
.B(n_559),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_513),
.B(n_493),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_542),
.B(n_549),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_508),
.B(n_501),
.C(n_505),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_544),
.B(n_551),
.C(n_553),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_529),
.A2(n_467),
.B1(n_479),
.B2(n_490),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_510),
.A2(n_460),
.B(n_496),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_534),
.B(n_492),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g571 ( 
.A(n_550),
.B(n_516),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_533),
.B(n_479),
.C(n_491),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_515),
.B(n_497),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_552),
.B(n_518),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_533),
.B(n_427),
.C(n_422),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_503),
.A2(n_495),
.B1(n_452),
.B2(n_422),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_503),
.A2(n_452),
.B1(n_427),
.B2(n_451),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_560),
.A2(n_526),
.B1(n_507),
.B2(n_506),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_511),
.B(n_522),
.C(n_525),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_561),
.B(n_562),
.C(n_500),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_522),
.B(n_285),
.C(n_342),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_563),
.B(n_565),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g565 ( 
.A(n_516),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_514),
.B(n_532),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_566),
.B(n_520),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_523),
.A2(n_468),
.B(n_451),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_567),
.B(n_526),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_498),
.A2(n_451),
.B1(n_342),
.B2(n_312),
.Y(n_568)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_568),
.Y(n_580)
);

FAx1_ASAP7_75t_SL g570 ( 
.A(n_548),
.B(n_517),
.CI(n_515),
.CON(n_570),
.SN(n_570)
);

A2O1A1O1Ixp25_ASAP7_75t_L g609 ( 
.A1(n_570),
.A2(n_550),
.B(n_563),
.C(n_556),
.D(n_564),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_571),
.B(n_585),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_561),
.Y(n_572)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_572),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_567),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_573),
.B(n_576),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_545),
.B(n_504),
.Y(n_576)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_547),
.Y(n_582)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_582),
.Y(n_601)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_584),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_541),
.B(n_502),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_586),
.B(n_591),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_587),
.B(n_562),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_540),
.B(n_504),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_589),
.B(n_595),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_590),
.A2(n_555),
.B(n_554),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_544),
.B(n_502),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_558),
.Y(n_592)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_592),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_593),
.A2(n_557),
.B1(n_539),
.B2(n_556),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_565),
.B(n_507),
.Y(n_594)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_594),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_566),
.B(n_524),
.C(n_499),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_594),
.B(n_499),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_597),
.B(n_600),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_577),
.B(n_553),
.C(n_551),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_598),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_577),
.B(n_543),
.C(n_558),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_599),
.B(n_602),
.C(n_613),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_592),
.B(n_564),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_587),
.B(n_546),
.C(n_536),
.Y(n_602)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_605),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_578),
.Y(n_608)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_608),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_L g623 ( 
.A1(n_609),
.A2(n_574),
.B(n_585),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_610),
.B(n_580),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_575),
.B(n_586),
.C(n_595),
.Y(n_613)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_614),
.Y(n_625)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_593),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_615),
.B(n_569),
.Y(n_630)
);

AOI321xp33_ASAP7_75t_L g616 ( 
.A1(n_570),
.A2(n_559),
.A3(n_555),
.B1(n_506),
.B2(n_538),
.C(n_521),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_616),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_574),
.A2(n_538),
.B(n_535),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_618),
.A2(n_590),
.B(n_579),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_597),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_620),
.B(n_624),
.Y(n_643)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_613),
.B(n_575),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_621),
.B(n_628),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_623),
.B(n_626),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_618),
.A2(n_581),
.B1(n_578),
.B2(n_588),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_599),
.B(n_591),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_605),
.A2(n_581),
.B1(n_569),
.B2(n_498),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_629),
.B(n_632),
.Y(n_651)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_630),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_616),
.A2(n_579),
.B(n_583),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_631),
.A2(n_604),
.B(n_570),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_603),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_633),
.B(n_638),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_598),
.B(n_571),
.C(n_509),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_635),
.B(n_610),
.C(n_602),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_600),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_637),
.A2(n_608),
.B1(n_611),
.B2(n_614),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_641),
.B(n_644),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_634),
.B(n_596),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_642),
.B(n_645),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_SL g644 ( 
.A1(n_623),
.A2(n_612),
.B(n_609),
.Y(n_644)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_648),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_627),
.B(n_601),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_649),
.B(n_650),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_627),
.B(n_617),
.C(n_607),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_628),
.B(n_617),
.C(n_607),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_652),
.B(n_624),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_SL g653 ( 
.A1(n_637),
.A2(n_606),
.B1(n_521),
.B2(n_530),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_653),
.B(n_654),
.Y(n_665)
);

XNOR2xp5_ASAP7_75t_L g654 ( 
.A(n_635),
.B(n_390),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_645),
.B(n_621),
.C(n_631),
.Y(n_657)
);

XNOR2xp5_ASAP7_75t_L g671 ( 
.A(n_657),
.B(n_661),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_640),
.A2(n_636),
.B1(n_625),
.B2(n_619),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_658),
.A2(n_636),
.B1(n_625),
.B2(n_648),
.Y(n_670)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_641),
.Y(n_660)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_660),
.Y(n_669)
);

XNOR2xp5_ASAP7_75t_L g663 ( 
.A(n_650),
.B(n_630),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_663),
.B(n_647),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_647),
.B(n_619),
.Y(n_664)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_664),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_639),
.B(n_622),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_666),
.A2(n_646),
.B(n_626),
.Y(n_673)
);

INVxp67_ASAP7_75t_SL g678 ( 
.A(n_667),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_655),
.B(n_652),
.C(n_654),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_668),
.A2(n_670),
.B(n_675),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_SL g672 ( 
.A1(n_659),
.A2(n_643),
.B1(n_651),
.B2(n_622),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_SL g676 ( 
.A1(n_672),
.A2(n_666),
.B(n_662),
.C(n_656),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_SL g679 ( 
.A(n_673),
.B(n_665),
.C(n_386),
.Y(n_679)
);

AOI21x1_ASAP7_75t_L g675 ( 
.A1(n_656),
.A2(n_646),
.B(n_629),
.Y(n_675)
);

AOI322xp5_ASAP7_75t_L g683 ( 
.A1(n_676),
.A2(n_680),
.A3(n_299),
.B1(n_161),
.B2(n_238),
.C1(n_259),
.C2(n_250),
.Y(n_683)
);

AOI21x1_ASAP7_75t_L g677 ( 
.A1(n_669),
.A2(n_665),
.B(n_390),
.Y(n_677)
);

A2O1A1O1Ixp25_ASAP7_75t_L g681 ( 
.A1(n_677),
.A2(n_679),
.B(n_674),
.C(n_668),
.D(n_667),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_681),
.A2(n_682),
.B(n_327),
.Y(n_685)
);

MAJIxp5_ASAP7_75t_L g682 ( 
.A(n_678),
.B(n_671),
.C(n_231),
.Y(n_682)
);

AO21x1_ASAP7_75t_L g684 ( 
.A1(n_683),
.A2(n_259),
.B(n_361),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_684),
.B(n_685),
.C(n_327),
.Y(n_686)
);

O2A1O1Ixp33_ASAP7_75t_SL g687 ( 
.A1(n_686),
.A2(n_13),
.B(n_14),
.C(n_361),
.Y(n_687)
);

XNOR2xp5_ASAP7_75t_L g688 ( 
.A(n_687),
.B(n_13),
.Y(n_688)
);

MAJIxp5_ASAP7_75t_L g689 ( 
.A(n_688),
.B(n_13),
.C(n_14),
.Y(n_689)
);


endmodule