module fake_jpeg_11734_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_11),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_6),
.B(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_25),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_10),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_1),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_89),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_57),
.B1(n_61),
.B2(n_48),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_54),
.B1(n_59),
.B2(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_63),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_68),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_48),
.B1(n_54),
.B2(n_59),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_60),
.C(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_53),
.Y(n_108)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_103),
.Y(n_126)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_114),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_56),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_58),
.B1(n_52),
.B2(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_112),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_116),
.C(n_2),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_6),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_51),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_113),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_60),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_83),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_29),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_60),
.B1(n_3),
.B2(n_4),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_66),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_9),
.C(n_10),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_138),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_33),
.C(n_46),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_4),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_5),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_5),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_136),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_34),
.C(n_45),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_7),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_132),
.B(n_137),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_7),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_135),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_8),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_35),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_8),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_144),
.C(n_145),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_36),
.C(n_44),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_16),
.B1(n_18),
.B2(n_21),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_149),
.C(n_152),
.Y(n_156)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_119),
.B(n_22),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_24),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_37),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_121),
.B1(n_136),
.B2(n_134),
.C(n_42),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_153),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_163),
.B(n_156),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_143),
.C(n_155),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_164),
.A2(n_139),
.B1(n_142),
.B2(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_166),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_159),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_168),
.B(n_147),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_139),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_161),
.B(n_150),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_38),
.Y(n_172)
);


endmodule