module fake_jpeg_30903_n_445 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_445);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_445;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_52),
.Y(n_133)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_54),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_21),
.B(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_86),
.Y(n_101)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_85),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_30),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_8),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_44),
.Y(n_130)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_29),
.B(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_29),
.B(n_8),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_90),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_43),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_19),
.B1(n_43),
.B2(n_27),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_93),
.A2(n_106),
.B1(n_115),
.B2(n_116),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_105),
.B(n_117),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_48),
.A2(n_27),
.B1(n_43),
.B2(n_30),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_57),
.A2(n_44),
.B1(n_42),
.B2(n_38),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_49),
.A2(n_27),
.B1(n_43),
.B2(n_20),
.Y(n_116)
);

BUFx2_ASAP7_75t_R g121 ( 
.A(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_36),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_50),
.A2(n_27),
.B1(n_43),
.B2(n_20),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_129),
.A2(n_87),
.B1(n_54),
.B2(n_64),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_37),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_33),
.C(n_25),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_89),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_52),
.A2(n_60),
.B1(n_81),
.B2(n_78),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_56),
.B1(n_55),
.B2(n_76),
.Y(n_170)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_140),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_158),
.Y(n_195)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_148),
.Y(n_194)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_169),
.B1(n_116),
.B2(n_129),
.Y(n_191)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_101),
.B(n_34),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_25),
.B1(n_15),
.B2(n_28),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_105),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_162),
.Y(n_201)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_174),
.Y(n_215)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_167),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_102),
.B(n_42),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_172),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_113),
.A2(n_28),
.B1(n_33),
.B2(n_27),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_170),
.A2(n_175),
.B1(n_185),
.B2(n_37),
.Y(n_222)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_130),
.B(n_38),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_114),
.A2(n_66),
.B1(n_63),
.B2(n_91),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_106),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_179),
.Y(n_217)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_177),
.Y(n_213)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_94),
.Y(n_179)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_95),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_182),
.Y(n_212)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_103),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_183),
.B(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_107),
.A2(n_135),
.B1(n_126),
.B2(n_100),
.Y(n_185)
);

XNOR2x1_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_99),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_191),
.A2(n_208),
.B1(n_186),
.B2(n_177),
.Y(n_237)
);

AOI22x1_ASAP7_75t_L g192 ( 
.A1(n_143),
.A2(n_128),
.B1(n_122),
.B2(n_120),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_192),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_139),
.B1(n_93),
.B2(n_133),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_183),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_145),
.A2(n_137),
.B1(n_133),
.B2(n_100),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_180),
.A2(n_137),
.B1(n_109),
.B2(n_110),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_154),
.A2(n_110),
.B1(n_109),
.B2(n_125),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_220),
.A2(n_183),
.B1(n_165),
.B2(n_160),
.Y(n_229)
);

OAI22x1_ASAP7_75t_SL g221 ( 
.A1(n_180),
.A2(n_120),
.B1(n_99),
.B2(n_16),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_222),
.B1(n_186),
.B2(n_144),
.Y(n_232)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_225),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_226),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_193),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_240),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_221),
.A2(n_150),
.B1(n_184),
.B2(n_181),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_228),
.A2(n_236),
.B(n_190),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_232),
.B1(n_238),
.B2(n_255),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_252),
.B1(n_230),
.B2(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_171),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_239),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_191),
.A2(n_178),
.B1(n_157),
.B2(n_173),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_242),
.B(n_249),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_204),
.A2(n_222),
.B1(n_192),
.B2(n_208),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_152),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_223),
.Y(n_240)
);

INVx4_ASAP7_75t_SL g241 ( 
.A(n_200),
.Y(n_241)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

NOR2x1_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_168),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_212),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_248),
.Y(n_258)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_244),
.Y(n_263)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_245),
.Y(n_284)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_247),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_195),
.B(n_155),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_204),
.A2(n_151),
.B(n_34),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_217),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_254),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_195),
.B(n_149),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_253),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_192),
.A2(n_147),
.B1(n_182),
.B2(n_166),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_210),
.A2(n_202),
.B1(n_194),
.B2(n_201),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_271),
.B1(n_242),
.B2(n_243),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_215),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_266),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_201),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_267),
.B(n_268),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_207),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_197),
.B(n_194),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_269),
.A2(n_257),
.B(n_275),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_230),
.A2(n_205),
.B1(n_218),
.B2(n_199),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_238),
.A2(n_197),
.B1(n_218),
.B2(n_199),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_262),
.B1(n_231),
.B2(n_284),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_200),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_276),
.B(n_278),
.Y(n_289)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_232),
.A2(n_213),
.A3(n_163),
.B1(n_189),
.B2(n_187),
.Y(n_277)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_190),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_216),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_280),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_251),
.B(n_211),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_211),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_224),
.C(n_225),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_285),
.A2(n_7),
.B(n_14),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_286),
.A2(n_280),
.B1(n_269),
.B2(n_270),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_242),
.B(n_252),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_287),
.A2(n_7),
.B(n_13),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_265),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_290),
.A2(n_302),
.B1(n_303),
.B2(n_283),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_234),
.Y(n_291)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_291),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_SL g340 ( 
.A1(n_292),
.A2(n_297),
.B(n_308),
.C(n_313),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_233),
.C(n_246),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_265),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_260),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_294),
.B(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_254),
.C(n_213),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_306),
.C(n_307),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_SL g297 ( 
.A1(n_271),
.A2(n_229),
.B(n_241),
.C(n_226),
.Y(n_297)
);

AND2x2_ASAP7_75t_SL g298 ( 
.A(n_275),
.B(n_241),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_298),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_274),
.B(n_240),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_211),
.Y(n_300)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_300),
.Y(n_337)
);

OAI32xp33_ASAP7_75t_L g301 ( 
.A1(n_274),
.A2(n_244),
.A3(n_187),
.B1(n_214),
.B2(n_189),
.Y(n_301)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_262),
.A2(n_205),
.B1(n_248),
.B2(n_219),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_273),
.A2(n_248),
.B1(n_188),
.B2(n_214),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_188),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_179),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_261),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_264),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_314),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_258),
.A2(n_9),
.B(n_14),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_316),
.B(n_318),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_290),
.A2(n_284),
.B1(n_277),
.B2(n_285),
.Y(n_318)
);

AOI21xp33_ASAP7_75t_L g319 ( 
.A1(n_308),
.A2(n_269),
.B(n_272),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_319),
.B(n_331),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_312),
.Y(n_320)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_320),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_304),
.A2(n_261),
.B1(n_272),
.B2(n_270),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_322),
.A2(n_324),
.B1(n_303),
.B2(n_298),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_304),
.Y(n_325)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_325),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_328),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_263),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_336),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_298),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_305),
.B(n_263),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_332),
.B(n_335),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_16),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_307),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_291),
.B(n_7),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_16),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_338),
.A2(n_287),
.B(n_297),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_286),
.A2(n_5),
.B1(n_12),
.B2(n_2),
.Y(n_339)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_339),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_345),
.Y(n_374)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_363),
.Y(n_381)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_289),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_351),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_296),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_352),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_353),
.A2(n_359),
.B1(n_364),
.B2(n_340),
.Y(n_379)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_354),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_288),
.C(n_311),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_328),
.C(n_336),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_314),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_357),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_321),
.A2(n_302),
.B1(n_313),
.B2(n_297),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_315),
.B(n_292),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_360),
.B(n_362),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_311),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_338),
.Y(n_364)
);

MAJx2_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_329),
.C(n_326),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_370),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_375),
.C(n_383),
.Y(n_384)
);

OAI21xp33_ASAP7_75t_L g370 ( 
.A1(n_348),
.A2(n_349),
.B(n_357),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_333),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_372),
.B(n_378),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_354),
.B1(n_358),
.B2(n_356),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_373),
.A2(n_353),
.B1(n_359),
.B2(n_350),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_293),
.C(n_318),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_316),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_362),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_345),
.Y(n_382)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_382),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_330),
.C(n_340),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_392),
.Y(n_401)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_388),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_381),
.C(n_367),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_389),
.B(n_390),
.C(n_391),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_343),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_343),
.C(n_350),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_371),
.A2(n_346),
.B(n_340),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_372),
.B(n_347),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_395),
.C(n_396),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_330),
.C(n_340),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_365),
.B(n_344),
.C(n_361),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_382),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_397),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_366),
.A2(n_297),
.B1(n_301),
.B2(n_2),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_398),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_4),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_3),
.C(n_10),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_399),
.Y(n_403)
);

INVx11_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

OAI21x1_ASAP7_75t_L g404 ( 
.A1(n_385),
.A2(n_376),
.B(n_369),
.Y(n_404)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_404),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_395),
.A2(n_368),
.B(n_380),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_384),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_388),
.A2(n_368),
.B(n_396),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_408),
.A2(n_412),
.B(n_11),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_394),
.A2(n_377),
.B1(n_374),
.B2(n_2),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_411),
.Y(n_419)
);

MAJx2_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_3),
.C(n_4),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_410),
.B(n_0),
.Y(n_422)
);

OAI21x1_ASAP7_75t_SL g412 ( 
.A1(n_385),
.A2(n_3),
.B(n_11),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_384),
.C(n_389),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_414),
.B(n_415),
.Y(n_426)
);

OAI21xp33_ASAP7_75t_L g416 ( 
.A1(n_401),
.A2(n_387),
.B(n_393),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_416),
.A2(n_400),
.B(n_407),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_390),
.C(n_16),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_423),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_422),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_406),
.B(n_0),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_0),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_411),
.C(n_410),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_415),
.A2(n_405),
.B(n_408),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_425),
.A2(n_417),
.B(n_424),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_429),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_401),
.C(n_400),
.Y(n_429)
);

BUFx24_ASAP7_75t_SL g431 ( 
.A(n_420),
.Y(n_431)
);

A2O1A1O1Ixp25_ASAP7_75t_L g436 ( 
.A1(n_431),
.A2(n_432),
.B(n_416),
.C(n_421),
.D(n_403),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_434),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_427),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_435),
.A2(n_436),
.B1(n_421),
.B2(n_432),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_426),
.B(n_413),
.C(n_419),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_437),
.A2(n_433),
.B(n_430),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_439),
.A2(n_440),
.B(n_422),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_441),
.A2(n_438),
.B(n_1),
.Y(n_442)
);

BUFx24_ASAP7_75t_SL g443 ( 
.A(n_442),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_443),
.A2(n_1),
.B(n_426),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_444),
.A2(n_1),
.B(n_57),
.Y(n_445)
);


endmodule