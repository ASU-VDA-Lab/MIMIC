module fake_jpeg_15482_n_386 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_386);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_386;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_39),
.Y(n_102)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_43),
.B(n_55),
.Y(n_98)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

NAND2x1_ASAP7_75t_SL g46 ( 
.A(n_14),
.B(n_0),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_46),
.B(n_52),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_62),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_1),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_36),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_69),
.B(n_71),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_36),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_72),
.B(n_80),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_36),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_73),
.B(n_87),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_19),
.B1(n_16),
.B2(n_24),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_74),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_76),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_39),
.Y(n_77)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_19),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_84),
.B(n_86),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_30),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_26),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_94),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_28),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

BUFx10_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_44),
.B(n_26),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_42),
.B(n_18),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_30),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_22),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_47),
.B(n_28),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_28),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_22),
.B1(n_30),
.B2(n_34),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_67),
.B1(n_60),
.B2(n_38),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_64),
.A2(n_18),
.B1(n_34),
.B2(n_27),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_28),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_121),
.B(n_125),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_24),
.B1(n_20),
.B2(n_18),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_122),
.A2(n_127),
.B1(n_162),
.B2(n_113),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_123),
.B(n_10),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_22),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_97),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_126),
.B(n_153),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_91),
.A2(n_25),
.B1(n_20),
.B2(n_34),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_52),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_53),
.B1(n_41),
.B2(n_24),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_132),
.A2(n_133),
.B1(n_146),
.B2(n_148),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_70),
.A2(n_20),
.B1(n_25),
.B2(n_27),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_138),
.A2(n_141),
.B1(n_163),
.B2(n_108),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_87),
.A2(n_38),
.B1(n_31),
.B2(n_57),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_118),
.B1(n_82),
.B2(n_81),
.Y(n_182)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_70),
.A2(n_67),
.B1(n_60),
.B2(n_31),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_31),
.B1(n_32),
.B2(n_17),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_31),
.B1(n_32),
.B2(n_17),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_150),
.A2(n_159),
.B1(n_170),
.B2(n_93),
.Y(n_193)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_187)
);

AOI32xp33_ASAP7_75t_L g153 ( 
.A1(n_75),
.A2(n_32),
.A3(n_17),
.B1(n_15),
.B2(n_28),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_156),
.Y(n_179)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_158),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_89),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_2),
.C(n_7),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_105),
.C(n_76),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_102),
.A2(n_2),
.B1(n_8),
.B2(n_9),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_103),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_167),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_111),
.B(n_8),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_10),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_100),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_79),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_181),
.B(n_183),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_182),
.A2(n_165),
.B1(n_168),
.B2(n_126),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_134),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_123),
.B(n_98),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_190),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_200),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_187),
.A2(n_99),
.B1(n_154),
.B2(n_13),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_188),
.A2(n_201),
.B1(n_152),
.B2(n_141),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_147),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_189),
.B(n_192),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_95),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_135),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_193),
.A2(n_204),
.B1(n_213),
.B2(n_88),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_161),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_151),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_216),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_124),
.B(n_130),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_198),
.B(n_199),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_78),
.B1(n_93),
.B2(n_108),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_128),
.B(n_120),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_202),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_148),
.B(n_150),
.C(n_169),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_203),
.B(n_185),
.Y(n_258)
);

OAI22x1_ASAP7_75t_SL g204 ( 
.A1(n_143),
.A2(n_88),
.B1(n_116),
.B2(n_102),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_208),
.Y(n_250)
);

NOR2x1_ASAP7_75t_R g206 ( 
.A(n_131),
.B(n_77),
.Y(n_206)
);

OR2x4_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_199),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_135),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_120),
.Y(n_215)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_143),
.B(n_116),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_144),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_144),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_218),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_129),
.A2(n_113),
.B1(n_12),
.B2(n_13),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_125),
.B1(n_121),
.B2(n_149),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_173),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_221),
.B(n_254),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_222),
.A2(n_226),
.B1(n_230),
.B2(n_236),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_225),
.A2(n_235),
.B(n_244),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_131),
.C(n_136),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_183),
.C(n_208),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_204),
.A2(n_131),
.B1(n_142),
.B2(n_137),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_229),
.A2(n_178),
.B(n_179),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_137),
.B1(n_159),
.B2(n_172),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_232),
.A2(n_234),
.B1(n_241),
.B2(n_242),
.Y(n_280)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_196),
.A2(n_172),
.B1(n_134),
.B2(n_158),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_196),
.A2(n_11),
.B(n_12),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_255),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_191),
.A2(n_99),
.B1(n_100),
.B2(n_154),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_239),
.A2(n_243),
.B1(n_247),
.B2(n_256),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_177),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_191),
.A2(n_11),
.B1(n_12),
.B2(n_216),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_202),
.A2(n_176),
.B(n_215),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_177),
.A2(n_209),
.B1(n_182),
.B2(n_193),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_245),
.A2(n_226),
.B1(n_232),
.B2(n_252),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_187),
.A2(n_195),
.B1(n_176),
.B2(n_209),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_181),
.B(n_199),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_253),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_249),
.A2(n_244),
.B(n_248),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_184),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_207),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_194),
.A2(n_185),
.B1(n_201),
.B2(n_198),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_175),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_189),
.B(n_192),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_197),
.Y(n_282)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_263),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_267),
.C(n_271),
.Y(n_296)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

AO22x1_ASAP7_75t_SL g266 ( 
.A1(n_245),
.A2(n_174),
.B1(n_175),
.B2(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

NAND2x1_ASAP7_75t_SL g269 ( 
.A(n_249),
.B(n_174),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_269),
.A2(n_273),
.B(n_275),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_180),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_282),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_240),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_227),
.B(n_180),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_272),
.B(n_276),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_238),
.A2(n_178),
.B(n_179),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_260),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_214),
.C(n_174),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_293),
.C(n_243),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_225),
.A2(n_212),
.B1(n_197),
.B2(n_200),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_279),
.A2(n_289),
.B(n_291),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_283),
.A2(n_286),
.B1(n_280),
.B2(n_277),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_250),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_287),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_225),
.A2(n_256),
.B1(n_230),
.B2(n_255),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_259),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_224),
.B(n_257),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

OAI21xp33_ASAP7_75t_L g289 ( 
.A1(n_223),
.A2(n_253),
.B(n_231),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_233),
.Y(n_290)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_246),
.Y(n_292)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_223),
.B(n_247),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_286),
.A2(n_229),
.B1(n_241),
.B2(n_246),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_294),
.A2(n_301),
.B1(n_303),
.B2(n_317),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_297),
.B(n_298),
.C(n_308),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_228),
.C(n_239),
.Y(n_298)
);

OA22x2_ASAP7_75t_L g300 ( 
.A1(n_266),
.A2(n_221),
.B1(n_237),
.B2(n_234),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_300),
.A2(n_315),
.B1(n_299),
.B2(n_309),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_269),
.A2(n_292),
.B1(n_273),
.B2(n_284),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_283),
.A2(n_220),
.B1(n_242),
.B2(n_259),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_265),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_263),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_271),
.B(n_293),
.C(n_262),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_265),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_311),
.B(n_304),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_235),
.C(n_281),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_314),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_269),
.A2(n_268),
.B(n_276),
.Y(n_314)
);

XNOR2x1_ASAP7_75t_L g316 ( 
.A(n_268),
.B(n_279),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_314),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_266),
.A2(n_280),
.B1(n_264),
.B2(n_281),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_264),
.A2(n_275),
.B1(n_274),
.B2(n_278),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_319),
.A2(n_303),
.B1(n_313),
.B2(n_300),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_270),
.Y(n_321)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_321),
.Y(n_344)
);

FAx1_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_290),
.CI(n_261),
.CON(n_322),
.SN(n_322)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_333),
.Y(n_343)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_324),
.A2(n_330),
.B1(n_331),
.B2(n_340),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_306),
.Y(n_325)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_325),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_306),
.Y(n_327)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_327),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_318),
.B(n_320),
.Y(n_329)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_329),
.Y(n_356)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_301),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_300),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_299),
.A2(n_317),
.B1(n_294),
.B2(n_319),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_334),
.A2(n_324),
.B1(n_327),
.B2(n_332),
.Y(n_353)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_335),
.B(n_337),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_302),
.Y(n_346)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_300),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_332),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_302),
.Y(n_340)
);

XNOR2x1_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_310),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_341),
.B(n_346),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_308),
.C(n_296),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_348),
.C(n_328),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_296),
.C(n_297),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_337),
.A2(n_333),
.B1(n_340),
.B2(n_326),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_351),
.B1(n_322),
.B2(n_339),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_326),
.A2(n_298),
.B1(n_318),
.B2(n_325),
.Y(n_351)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_353),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_355),
.B(n_334),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_358),
.Y(n_372)
);

NAND3xp33_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_322),
.C(n_330),
.Y(n_359)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_359),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_SL g361 ( 
.A(n_344),
.B(n_328),
.C(n_335),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_362),
.Y(n_371)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_350),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_366),
.C(n_348),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_350),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_364),
.B(n_365),
.C(n_345),
.Y(n_369)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_354),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_343),
.A2(n_356),
.B(n_345),
.Y(n_366)
);

FAx1_ASAP7_75t_SL g368 ( 
.A(n_357),
.B(n_343),
.CI(n_346),
.CON(n_368),
.SN(n_368)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_368),
.B(n_369),
.Y(n_375)
);

MAJx2_ASAP7_75t_L g377 ( 
.A(n_373),
.B(n_363),
.C(n_347),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_370),
.A2(n_360),
.B1(n_355),
.B2(n_351),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_374),
.B(n_376),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_369),
.A2(n_349),
.B1(n_342),
.B2(n_359),
.Y(n_376)
);

AO21x1_ASAP7_75t_L g378 ( 
.A1(n_377),
.A2(n_373),
.B(n_371),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_378),
.A2(n_377),
.B(n_368),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_379),
.A2(n_352),
.B1(n_375),
.B2(n_353),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_380),
.B(n_381),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_382),
.B(n_368),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_372),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_384),
.A2(n_372),
.B(n_367),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_367),
.Y(n_386)
);


endmodule