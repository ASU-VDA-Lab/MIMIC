module fake_jpeg_27673_n_102 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx24_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVxp33_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_26),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_28),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_35),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_23),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_15),
.B1(n_13),
.B2(n_3),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_21),
.C(n_14),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_35),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_15),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_31),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_46),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_19),
.B1(n_11),
.B2(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_44),
.B1(n_13),
.B2(n_4),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_11),
.B1(n_22),
.B2(n_16),
.Y(n_44)
);

NOR3xp33_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_13),
.C(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_1),
.Y(n_60)
);

AND2x6_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_58),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_55),
.Y(n_68)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_59),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_33),
.C(n_37),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_49),
.C(n_45),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_41),
.Y(n_62)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_41),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_48),
.B(n_44),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_53),
.B(n_5),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_5),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_4),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_75),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_65),
.B1(n_70),
.B2(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_76),
.Y(n_83)
);

AOI322xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_50),
.A3(n_54),
.B1(n_55),
.B2(n_51),
.C1(n_58),
.C2(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_4),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_66),
.C(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_82),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_63),
.C(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_85),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_86),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_78),
.C(n_80),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_76),
.B(n_72),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_72),
.B(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_95),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_89),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_70),
.B(n_79),
.C(n_7),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_98),
.C(n_95),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_5),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_100),
.B(n_8),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_9),
.Y(n_102)
);


endmodule