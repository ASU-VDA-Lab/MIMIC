module fake_jpeg_30934_n_82 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_82);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_82;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_13),
.B1(n_24),
.B2(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_0),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_35),
.B1(n_29),
.B2(n_30),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_2),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_28),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_36),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_30),
.C(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_5),
.Y(n_56)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_54),
.B1(n_9),
.B2(n_11),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_3),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_65),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_47),
.B(n_10),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_68),
.B1(n_69),
.B2(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_14),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_72),
.C(n_62),
.Y(n_75)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_67),
.B(n_20),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_72),
.C(n_76),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_67),
.B(n_74),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_73),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_19),
.B(n_22),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_25),
.Y(n_82)
);


endmodule