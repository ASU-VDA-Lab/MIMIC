module fake_jpeg_30789_n_194 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_194);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_5),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_23),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_24),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_3),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_54),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_33),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_28),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_67),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_34),
.A2(n_26),
.B1(n_30),
.B2(n_17),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_24),
.B1(n_28),
.B2(n_19),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_16),
.B1(n_28),
.B2(n_19),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_26),
.B1(n_30),
.B2(n_27),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_28),
.B1(n_19),
.B2(n_16),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_0),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_9),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_39),
.B(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_9),
.Y(n_87)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_91),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_86),
.B1(n_74),
.B2(n_72),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_84),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_97),
.B1(n_50),
.B2(n_56),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_19),
.Y(n_84)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_31),
.CI(n_46),
.CON(n_85),
.SN(n_85)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_31),
.B1(n_3),
.B2(n_0),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_31),
.C(n_3),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_5),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_78),
.Y(n_111)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_10),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_56),
.B(n_4),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_113),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_72),
.B1(n_59),
.B2(n_75),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_80),
.B1(n_86),
.B2(n_82),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_112),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_53),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_53),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_114),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_59),
.B1(n_75),
.B2(n_74),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_100),
.B1(n_98),
.B2(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_130),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_97),
.B(n_99),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_140),
.B1(n_116),
.B2(n_119),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_85),
.B(n_84),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_85),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_135),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_88),
.B1(n_93),
.B2(n_77),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_136),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_76),
.B1(n_12),
.B2(n_14),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_138),
.A2(n_141),
.B1(n_121),
.B2(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_6),
.B1(n_12),
.B2(n_15),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_15),
.B1(n_107),
.B2(n_102),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_137),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_151),
.B1(n_152),
.B2(n_126),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_104),
.C(n_106),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_154),
.C(n_141),
.Y(n_159)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_121),
.B1(n_106),
.B2(n_104),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_129),
.C(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_137),
.B(n_131),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_153),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_160),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_164),
.C(n_166),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_137),
.B1(n_138),
.B2(n_125),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_163),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_146),
.C(n_143),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_153),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_150),
.C(n_155),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_169),
.C(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_177),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_143),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_179),
.Y(n_183)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_180),
.A2(n_161),
.B1(n_163),
.B2(n_142),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_157),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_167),
.C(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_144),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_186),
.A2(n_185),
.B(n_182),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_184),
.A2(n_174),
.B1(n_160),
.B2(n_152),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_183),
.B1(n_181),
.B2(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_191),
.B(n_190),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_192),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_165),
.Y(n_194)
);


endmodule