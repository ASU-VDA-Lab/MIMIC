module fake_jpeg_18382_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_26),
.Y(n_44)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_53),
.Y(n_66)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_20),
.B1(n_26),
.B2(n_22),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_52),
.B1(n_39),
.B2(n_37),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_24),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_20),
.B1(n_26),
.B2(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_15),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_77),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_59),
.A2(n_60),
.B1(n_68),
.B2(n_45),
.Y(n_106)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_65),
.B(n_66),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_39),
.B(n_29),
.C(n_37),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_32),
.B1(n_37),
.B2(n_34),
.Y(n_95)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_16),
.B(n_31),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_20),
.B1(n_30),
.B2(n_22),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_34),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_76),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_75),
.B(n_24),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_34),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_24),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_39),
.C(n_35),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_37),
.B1(n_34),
.B2(n_42),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_35),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_101),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_108),
.B1(n_111),
.B2(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_103),
.B1(n_79),
.B2(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_65),
.B(n_51),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_15),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_34),
.B1(n_37),
.B2(n_42),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_72),
.B(n_15),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_23),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_42),
.B1(n_38),
.B2(n_36),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_42),
.B1(n_38),
.B2(n_36),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_67),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_116),
.B(n_136),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_69),
.C(n_80),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_111),
.B1(n_108),
.B2(n_93),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_76),
.B1(n_71),
.B2(n_70),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_119),
.A2(n_129),
.B1(n_93),
.B2(n_99),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_64),
.C(n_62),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_135),
.C(n_103),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_35),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_128),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_137),
.B1(n_100),
.B2(n_109),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_88),
.Y(n_126)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_35),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_84),
.A2(n_57),
.B1(n_55),
.B2(n_60),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_138),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_35),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_134),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_87),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_98),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_84),
.A2(n_81),
.B(n_22),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_21),
.B(n_18),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_95),
.A2(n_28),
.B1(n_23),
.B2(n_61),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_158),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_29),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_156),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_149),
.A2(n_29),
.B1(n_8),
.B2(n_10),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_85),
.Y(n_150)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_168),
.B1(n_152),
.B2(n_153),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_98),
.B(n_91),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_157),
.A2(n_16),
.B(n_31),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_119),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_38),
.B1(n_36),
.B2(n_30),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_118),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_164),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_169),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_163),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_165),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_91),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_113),
.A2(n_90),
.B1(n_88),
.B2(n_57),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_90),
.B1(n_55),
.B2(n_59),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_170),
.A2(n_38),
.B1(n_36),
.B2(n_30),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_155),
.A2(n_124),
.B1(n_115),
.B2(n_138),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_171),
.A2(n_193),
.B1(n_196),
.B2(n_141),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_113),
.A3(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_175),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_134),
.C(n_38),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_27),
.C(n_19),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_178),
.A2(n_191),
.B1(n_200),
.B2(n_170),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_28),
.B(n_23),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_179),
.A2(n_180),
.B(n_145),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_189),
.B1(n_168),
.B2(n_142),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_24),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_194),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_16),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_36),
.B1(n_28),
.B2(n_31),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_151),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_192),
.B(n_144),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_143),
.A2(n_146),
.B1(n_142),
.B2(n_141),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_29),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_143),
.A2(n_21),
.B1(n_18),
.B2(n_29),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_21),
.B1(n_18),
.B2(n_17),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_177),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_203),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_206),
.A2(n_207),
.B1(n_213),
.B2(n_215),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_175),
.A2(n_140),
.B1(n_169),
.B2(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_216),
.Y(n_225)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_212),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_190),
.A2(n_167),
.B1(n_164),
.B2(n_17),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_167),
.B1(n_164),
.B2(n_2),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_172),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_182),
.B(n_19),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_222),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_178),
.C(n_181),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_174),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_188),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_176),
.A2(n_27),
.B1(n_19),
.B2(n_2),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_171),
.A2(n_27),
.B1(n_19),
.B2(n_2),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_27),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_199),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_223),
.A2(n_238),
.B(n_201),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_229),
.C(n_232),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_183),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_231),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_183),
.C(n_187),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_173),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_195),
.C(n_185),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_179),
.Y(n_251)
);

XOR2x1_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_180),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_184),
.B1(n_200),
.B2(n_186),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_209),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_246),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_201),
.B(n_195),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_247),
.B(n_249),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_209),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_225),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_238),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_191),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_224),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_204),
.B1(n_220),
.B2(n_221),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_254),
.B1(n_213),
.B2(n_231),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_235),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_237),
.A2(n_215),
.B(n_207),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_227),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_253),
.C(n_241),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_260),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_236),
.C(n_253),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_196),
.C(n_7),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_229),
.C(n_228),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_262),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_242),
.C(n_224),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_267),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_218),
.C(n_232),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_254),
.B1(n_211),
.B2(n_252),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_268),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_270),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_264),
.A2(n_263),
.B(n_256),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_258),
.B(n_7),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_14),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_7),
.B(n_12),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_277),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_14),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_283),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_277),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_14),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_273),
.B(n_1),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_12),
.C(n_10),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_8),
.C(n_12),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_287),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_276),
.B1(n_1),
.B2(n_3),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_279),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_293),
.B(n_290),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_279),
.C(n_1),
.Y(n_293)
);

NAND3xp33_ASAP7_75t_SL g296 ( 
.A(n_294),
.B(n_295),
.C(n_0),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_288),
.B(n_4),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_296),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_0),
.C(n_4),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_5),
.B(n_294),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_5),
.Y(n_300)
);


endmodule