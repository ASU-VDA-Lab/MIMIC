module real_jpeg_33286_n_5 (n_4, n_0, n_21, n_1, n_2, n_22, n_3, n_5);

input n_4;
input n_0;
input n_21;
input n_1;
input n_2;
input n_22;
input n_3;

output n_5;

wire n_17;
wire n_8;
wire n_10;
wire n_9;
wire n_12;
wire n_6;
wire n_11;
wire n_14;
wire n_7;
wire n_18;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_0),
.B(n_21),
.Y(n_9)
);

AOI22xp33_ASAP7_75t_L g5 ( 
.A1(n_1),
.A2(n_6),
.B1(n_7),
.B2(n_19),
.Y(n_5)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

AOI221xp5_ASAP7_75t_L g7 ( 
.A1(n_3),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_7)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.C(n_11),
.Y(n_8)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_22),
.Y(n_10)
);


endmodule