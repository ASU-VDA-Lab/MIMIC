module fake_jpeg_12475_n_227 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_5),
.B(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_19),
.Y(n_56)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_73),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_26),
.B1(n_24),
.B2(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_60),
.A2(n_62),
.B1(n_70),
.B2(n_69),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_24),
.B1(n_31),
.B2(n_26),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_74),
.B1(n_34),
.B2(n_18),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_26),
.B1(n_17),
.B2(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_40),
.B(n_21),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_17),
.B1(n_33),
.B2(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_76),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_36),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_34),
.B(n_43),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_52),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_79),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_68),
.B(n_78),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_99),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_92),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_98),
.Y(n_127)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_94),
.Y(n_113)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_100),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_25),
.B1(n_21),
.B2(n_70),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_0),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_104),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_58),
.A2(n_18),
.B1(n_34),
.B2(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_103),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_0),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_124),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_15),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_57),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_72),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_86),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_18),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_67),
.C(n_64),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_90),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_83),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_131),
.B(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_81),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_132),
.B(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_125),
.A2(n_95),
.B(n_102),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_138),
.B(n_121),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_125),
.A2(n_87),
.B1(n_65),
.B2(n_94),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_140),
.B1(n_122),
.B2(n_108),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_113),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_139),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_79),
.B(n_96),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_89),
.B1(n_54),
.B2(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_100),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_146),
.B(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_54),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_150),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_67),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_64),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_8),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_15),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_120),
.B(n_1),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_159),
.B(n_143),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_107),
.B1(n_108),
.B2(n_117),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_136),
.B1(n_140),
.B2(n_146),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_110),
.B(n_126),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_119),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_169),
.C(n_148),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_141),
.B1(n_133),
.B2(n_137),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_165),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_109),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_168),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_123),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_174),
.B1(n_158),
.B2(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_161),
.A2(n_139),
.B1(n_117),
.B2(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_179),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_150),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_177),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_172),
.B(n_174),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_142),
.B1(n_128),
.B2(n_122),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_113),
.B1(n_114),
.B2(n_105),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_180),
.A2(n_181),
.B(n_154),
.Y(n_189)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_114),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_153),
.C(n_163),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_153),
.C(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_105),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_8),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_11),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_179),
.B1(n_180),
.B2(n_175),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_176),
.C(n_185),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_191),
.B(n_184),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_196),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_162),
.C(n_155),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_170),
.B(n_3),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_198),
.B(n_181),
.Y(n_200)
);

NOR3xp33_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_203),
.C(n_205),
.Y(n_212)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_202),
.B(n_204),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_170),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_207),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_11),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_196),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_213),
.B(n_214),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_193),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_193),
.C(n_198),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_211),
.A2(n_194),
.B1(n_206),
.B2(n_190),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_217),
.C(n_1),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_197),
.B(n_14),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_67),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_14),
.B1(n_5),
.B2(n_6),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_210),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_218),
.A2(n_1),
.B(n_6),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_221),
.C(n_222),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_219),
.B(n_59),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_223),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_218),
.C(n_59),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_224),
.Y(n_227)
);


endmodule