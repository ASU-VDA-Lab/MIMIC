module fake_jpeg_12721_n_579 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_579);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_579;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_60),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_61),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_62),
.B(n_76),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_20),
.A2(n_8),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_63),
.B(n_77),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_64),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_65),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_11),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_66),
.B(n_69),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_67),
.Y(n_183)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_11),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_71),
.Y(n_190)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_74),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_75),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_22),
.B(n_11),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_78),
.Y(n_202)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_24),
.B(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_96),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx16f_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_12),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_15),
.Y(n_133)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_84),
.Y(n_215)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_86),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_25),
.B(n_12),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_88),
.B(n_89),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_12),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_90),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_93),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_94),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_95),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_26),
.B(n_12),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g205 ( 
.A(n_97),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g148 ( 
.A(n_105),
.Y(n_148)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_106),
.Y(n_210)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

BUFx4f_ASAP7_75t_SL g196 ( 
.A(n_110),
.Y(n_196)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_115),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g147 ( 
.A(n_114),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_49),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g156 ( 
.A(n_116),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_28),
.B(n_6),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_117),
.B(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_119),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_57),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_28),
.B(n_6),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx6_ASAP7_75t_SL g165 ( 
.A(n_121),
.Y(n_165)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_122),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_124),
.Y(n_180)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_31),
.B(n_6),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_125),
.B(n_16),
.Y(n_175)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_33),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_126),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_128),
.Y(n_181)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_54),
.B1(n_56),
.B2(n_53),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_131),
.A2(n_134),
.B1(n_144),
.B2(n_172),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_133),
.A2(n_162),
.B(n_4),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_78),
.A2(n_56),
.B1(n_53),
.B2(n_47),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_62),
.B(n_52),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_136),
.B(n_143),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_52),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_59),
.A2(n_47),
.B1(n_44),
.B2(n_40),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_119),
.A2(n_21),
.B1(n_49),
.B2(n_37),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_150),
.A2(n_151),
.B1(n_160),
.B2(n_161),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_110),
.A2(n_21),
.B1(n_49),
.B2(n_33),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_113),
.A2(n_21),
.B1(n_49),
.B2(n_37),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_74),
.A2(n_21),
.B1(n_49),
.B2(n_37),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_104),
.A2(n_49),
.B(n_50),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_84),
.A2(n_42),
.B1(n_48),
.B2(n_23),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_164),
.A2(n_178),
.B1(n_197),
.B2(n_200),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_64),
.A2(n_42),
.B1(n_48),
.B2(n_23),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_171),
.A2(n_191),
.B1(n_137),
.B2(n_156),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_67),
.A2(n_40),
.B1(n_44),
.B2(n_50),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_175),
.B(n_192),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_97),
.A2(n_19),
.B1(n_48),
.B2(n_30),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_68),
.B(n_46),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_189),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_75),
.A2(n_30),
.B1(n_27),
.B2(n_23),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_184),
.A2(n_122),
.B1(n_126),
.B2(n_112),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_72),
.B(n_0),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_61),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_87),
.A2(n_30),
.B1(n_27),
.B2(n_19),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_188),
.A2(n_208),
.B1(n_214),
.B2(n_18),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_86),
.B(n_46),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_93),
.A2(n_27),
.B1(n_19),
.B2(n_13),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_82),
.B(n_5),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_106),
.A2(n_13),
.B1(n_17),
.B2(n_15),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_65),
.A2(n_13),
.B1(n_17),
.B2(n_15),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_114),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_204),
.A2(n_208),
.B(n_210),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_L g208 ( 
.A1(n_94),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_121),
.B(n_1),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_61),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_82),
.B(n_4),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_207),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_98),
.A2(n_99),
.B1(n_109),
.B2(n_116),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_219),
.B(n_223),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_220),
.A2(n_242),
.B1(n_244),
.B2(n_250),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_162),
.A2(n_124),
.B1(n_101),
.B2(n_102),
.Y(n_221)
);

OAI32xp33_ASAP7_75t_L g312 ( 
.A1(n_221),
.A2(n_235),
.A3(n_206),
.B1(n_196),
.B2(n_216),
.Y(n_312)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_222),
.Y(n_309)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_224),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_226),
.B(n_267),
.Y(n_320)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_227),
.Y(n_323)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_132),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_228),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_230),
.B(n_239),
.Y(n_317)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_143),
.Y(n_231)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_231),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_133),
.B(n_123),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_232),
.B(n_237),
.Y(n_302)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_156),
.Y(n_233)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_233),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_95),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_234),
.B(n_238),
.C(n_255),
.Y(n_298)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_184),
.A2(n_105),
.B1(n_14),
.B2(n_18),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_152),
.B1(n_154),
.B2(n_153),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_236),
.A2(n_278),
.B1(n_206),
.B2(n_216),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_4),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_18),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_168),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g240 ( 
.A(n_182),
.B(n_189),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_240),
.B(n_253),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_136),
.B(n_193),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_243),
.B(n_261),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_130),
.A2(n_155),
.B1(n_166),
.B2(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_245),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_246),
.Y(n_339)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_135),
.Y(n_248)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_248),
.Y(n_329)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_249),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_141),
.A2(n_140),
.B1(n_177),
.B2(n_152),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_252),
.B(n_254),
.Y(n_318)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_135),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_157),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_167),
.B(n_157),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_165),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_256),
.B(n_259),
.Y(n_324)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_145),
.B(n_129),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_284),
.C(n_196),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_165),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_260),
.A2(n_282),
.B1(n_224),
.B2(n_222),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_147),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_138),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_262),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_191),
.A2(n_195),
.B1(n_209),
.B2(n_137),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_263),
.A2(n_187),
.B1(n_215),
.B2(n_210),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_129),
.B(n_142),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_264),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_153),
.A2(n_145),
.B1(n_163),
.B2(n_146),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_268),
.B(n_282),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_147),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_270),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_142),
.B(n_159),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_207),
.A2(n_205),
.B1(n_209),
.B2(n_163),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_269),
.A2(n_280),
.B1(n_285),
.B2(n_286),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_169),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_159),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_271),
.Y(n_301)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_272),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_176),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_273),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_169),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_274),
.B(n_275),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_185),
.B(n_198),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_174),
.A2(n_146),
.B1(n_139),
.B2(n_183),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_201),
.B1(n_183),
.B2(n_202),
.Y(n_294)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_277),
.B(n_279),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_176),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_169),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_205),
.A2(n_138),
.B1(n_190),
.B2(n_149),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_210),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_281),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_149),
.B(n_179),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_174),
.B(n_179),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_287),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_190),
.B(n_170),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_190),
.A2(n_195),
.B1(n_170),
.B2(n_215),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_139),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_187),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_173),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_288),
.A2(n_290),
.B1(n_233),
.B2(n_271),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_173),
.B(n_201),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_237),
.Y(n_337)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_159),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_294),
.A2(n_305),
.B1(n_314),
.B2(n_316),
.Y(n_348)
);

AND2x2_ASAP7_75t_SL g295 ( 
.A(n_225),
.B(n_170),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_295),
.B(n_297),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_275),
.A2(n_210),
.B(n_206),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_300),
.A2(n_270),
.B(n_274),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_231),
.A2(n_196),
.B1(n_158),
.B2(n_216),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_306),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_311),
.Y(n_350)
);

OA21x2_ASAP7_75t_L g352 ( 
.A1(n_312),
.A2(n_344),
.B(n_284),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_241),
.A2(n_158),
.B1(n_240),
.B2(n_225),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_240),
.A2(n_158),
.B1(n_220),
.B2(n_255),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_321),
.Y(n_388)
);

O2A1O1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_223),
.A2(n_221),
.B(n_234),
.C(n_268),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_SL g364 ( 
.A1(n_326),
.A2(n_258),
.B(n_284),
.C(n_266),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_218),
.B(n_232),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_342),
.C(n_298),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_260),
.A2(n_226),
.B1(n_218),
.B2(n_247),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_342),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_276),
.A2(n_239),
.B1(n_230),
.B2(n_235),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_334),
.A2(n_335),
.B1(n_346),
.B2(n_316),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_223),
.A2(n_234),
.B1(n_235),
.B2(n_238),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_217),
.A2(n_221),
.B1(n_287),
.B2(n_249),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_336),
.A2(n_345),
.B1(n_344),
.B2(n_340),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_337),
.B(n_261),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_243),
.B(n_238),
.C(n_221),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_235),
.A2(n_289),
.B1(n_283),
.B2(n_265),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_227),
.A2(n_228),
.B1(n_254),
.B2(n_253),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_355),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_351),
.A2(n_352),
.B(n_368),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_310),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_353),
.B(n_358),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_354),
.B(n_338),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_308),
.B(n_229),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_313),
.Y(n_356)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_356),
.Y(n_391)
);

AO22x1_ASAP7_75t_SL g357 ( 
.A1(n_307),
.A2(n_277),
.B1(n_251),
.B2(n_257),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_357),
.B(n_361),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_310),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_258),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_371),
.C(n_380),
.Y(n_406)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_323),
.Y(n_360)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_302),
.B(n_256),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_313),
.Y(n_362)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_362),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_302),
.B(n_259),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_363),
.B(n_367),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_303),
.Y(n_365)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_365),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_314),
.A2(n_288),
.B1(n_286),
.B2(n_245),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_366),
.A2(n_379),
.B1(n_383),
.B2(n_311),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_308),
.B(n_248),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_322),
.B(n_279),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_369),
.B(n_376),
.Y(n_408)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_331),
.Y(n_370)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_298),
.B(n_290),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_372),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_326),
.A2(n_293),
.B(n_300),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_373),
.A2(n_291),
.B(n_304),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_296),
.A2(n_262),
.B(n_272),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_374),
.A2(n_377),
.B(n_299),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_322),
.B(n_246),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_296),
.A2(n_335),
.B(n_328),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_328),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_389),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_307),
.B(n_327),
.C(n_320),
.Y(n_380)
);

INVx11_ASAP7_75t_L g381 ( 
.A(n_301),
.Y(n_381)
);

BUFx5_ASAP7_75t_L g393 ( 
.A(n_381),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_317),
.B(n_341),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_382),
.B(n_387),
.Y(n_416)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_330),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_384),
.B(n_324),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_327),
.B(n_320),
.C(n_295),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_386),
.C(n_329),
.Y(n_415)
);

MAJx2_ASAP7_75t_L g386 ( 
.A(n_327),
.B(n_296),
.C(n_295),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_341),
.B(n_318),
.Y(n_387)
);

A2O1A1Ixp33_ASAP7_75t_L g389 ( 
.A1(n_295),
.A2(n_333),
.B(n_340),
.C(n_343),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_382),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_392),
.B(n_421),
.Y(n_441)
);

AND2x4_ASAP7_75t_SL g396 ( 
.A(n_364),
.B(n_330),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_396),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_398),
.A2(n_347),
.B1(n_350),
.B2(n_368),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_353),
.A2(n_292),
.B1(n_343),
.B2(n_293),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_400),
.A2(n_401),
.B1(n_405),
.B2(n_414),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_384),
.A2(n_292),
.B1(n_306),
.B2(n_312),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_404),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_403),
.A2(n_409),
.B(n_390),
.Y(n_431)
);

AND2x6_ASAP7_75t_L g404 ( 
.A(n_351),
.B(n_305),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_358),
.A2(n_294),
.B1(n_297),
.B2(n_339),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_373),
.A2(n_299),
.B(n_304),
.Y(n_409)
);

INVx8_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_411),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_399),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_361),
.A2(n_339),
.B1(n_346),
.B2(n_303),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_423),
.C(n_371),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_355),
.B(n_301),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_419),
.B(n_369),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g421 ( 
.A(n_387),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_363),
.A2(n_315),
.B1(n_329),
.B2(n_325),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_422),
.A2(n_366),
.B1(n_348),
.B2(n_375),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_367),
.B(n_315),
.Y(n_425)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_425),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_418),
.Y(n_427)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_428),
.A2(n_436),
.B1(n_445),
.B2(n_452),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_432),
.C(n_435),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_431),
.A2(n_443),
.B(n_409),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_354),
.C(n_385),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_433),
.A2(n_426),
.B1(n_439),
.B2(n_440),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_380),
.C(n_386),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_398),
.A2(n_347),
.B1(n_389),
.B2(n_352),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_437),
.B(n_448),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_438),
.B(n_395),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_401),
.A2(n_352),
.B1(n_383),
.B2(n_348),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_439),
.A2(n_440),
.B1(n_447),
.B2(n_394),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_400),
.A2(n_352),
.B1(n_375),
.B2(n_378),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_403),
.A2(n_377),
.B(n_364),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_406),
.B(n_386),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_450),
.C(n_451),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_398),
.A2(n_375),
.B1(n_349),
.B2(n_388),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_405),
.A2(n_356),
.B1(n_372),
.B2(n_370),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_416),
.B(n_359),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_392),
.A2(n_376),
.B1(n_362),
.B2(n_357),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_449),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_406),
.B(n_374),
.C(n_357),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_406),
.B(n_415),
.C(n_417),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_417),
.A2(n_357),
.B1(n_365),
.B2(n_360),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_413),
.A2(n_309),
.B1(n_325),
.B2(n_323),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_414),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_319),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_455),
.C(n_412),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_395),
.B(n_402),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_456),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_457),
.B(n_444),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_399),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_459),
.B(n_435),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_441),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_463),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_453),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_455),
.B(n_394),
.Y(n_464)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_464),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_416),
.Y(n_466)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_466),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_430),
.B(n_419),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_467),
.B(n_472),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_469),
.A2(n_473),
.B1(n_475),
.B2(n_446),
.Y(n_507)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_470),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_430),
.B(n_408),
.Y(n_471)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_471),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_408),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_434),
.B(n_422),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_480),
.Y(n_493)
);

OAI22xp33_ASAP7_75t_L g475 ( 
.A1(n_426),
.A2(n_410),
.B1(n_403),
.B2(n_425),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_476),
.A2(n_478),
.B(n_482),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_443),
.A2(n_409),
.B(n_396),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_434),
.B(n_404),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_396),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_431),
.A2(n_410),
.B(n_396),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_447),
.Y(n_483)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_483),
.Y(n_498)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_433),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_484),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_483),
.Y(n_486)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_486),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_432),
.C(n_451),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_487),
.B(n_499),
.C(n_500),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_413),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g526 ( 
.A(n_488),
.B(n_424),
.C(n_391),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_494),
.B(n_495),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_484),
.A2(n_442),
.B1(n_450),
.B2(n_404),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_496),
.A2(n_465),
.B1(n_482),
.B2(n_477),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_454),
.C(n_438),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_436),
.C(n_445),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_472),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_501),
.B(n_460),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_462),
.B(n_396),
.C(n_442),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_504),
.C(n_476),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_505),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_459),
.B(n_446),
.C(n_407),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_407),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_507),
.A2(n_474),
.B1(n_478),
.B2(n_470),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_492),
.A2(n_473),
.B1(n_465),
.B2(n_469),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_509),
.A2(n_513),
.B1(n_497),
.B2(n_489),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_510),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_507),
.A2(n_465),
.B1(n_477),
.B2(n_466),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_512),
.B(n_514),
.Y(n_528)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_491),
.Y(n_516)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_516),
.Y(n_530)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_491),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_519),
.Y(n_537)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_506),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_SL g539 ( 
.A(n_520),
.B(n_523),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_493),
.A2(n_471),
.B(n_480),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_522),
.A2(n_500),
.B(n_490),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_493),
.A2(n_467),
.B1(n_461),
.B2(n_464),
.Y(n_523)
);

OAI21xp33_ASAP7_75t_SL g524 ( 
.A1(n_498),
.A2(n_457),
.B(n_468),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_496),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_487),
.B(n_458),
.C(n_468),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_504),
.C(n_502),
.Y(n_531)
);

AOI31xp67_ASAP7_75t_SL g532 ( 
.A1(n_526),
.A2(n_485),
.A3(n_411),
.B(n_393),
.Y(n_532)
);

MAJx2_ASAP7_75t_L g542 ( 
.A(n_527),
.B(n_538),
.C(n_514),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_531),
.B(n_534),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_519),
.Y(n_545)
);

AO21x1_ASAP7_75t_L g533 ( 
.A1(n_516),
.A2(n_517),
.B(n_515),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_533),
.A2(n_486),
.B(n_497),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_525),
.B(n_499),
.C(n_505),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_509),
.A2(n_497),
.B1(n_489),
.B2(n_498),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_535),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_518),
.B(n_520),
.C(n_495),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_536),
.B(n_541),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_540),
.A2(n_513),
.B(n_490),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_518),
.B(n_503),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_542),
.B(n_546),
.C(n_531),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_545),
.B(n_549),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_521),
.C(n_511),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_529),
.B(n_523),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_548),
.B(n_551),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_539),
.A2(n_522),
.B(n_515),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_550),
.A2(n_552),
.B1(n_553),
.B2(n_533),
.Y(n_554)
);

NAND2x1_ASAP7_75t_SL g551 ( 
.A(n_530),
.B(n_521),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_540),
.A2(n_511),
.B(n_486),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_554),
.Y(n_567)
);

AOI322xp5_ASAP7_75t_L g556 ( 
.A1(n_547),
.A2(n_512),
.A3(n_527),
.B1(n_535),
.B2(n_537),
.C1(n_528),
.C2(n_458),
.Y(n_556)
);

AOI21xp33_ASAP7_75t_L g569 ( 
.A1(n_556),
.A2(n_562),
.B(n_555),
.Y(n_569)
);

CKINVDCx14_ASAP7_75t_R g557 ( 
.A(n_543),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_557),
.B(n_560),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_558),
.B(n_546),
.C(n_542),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_544),
.B(n_534),
.C(n_541),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_545),
.B(n_528),
.Y(n_561)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_561),
.Y(n_568)
);

AOI322xp5_ASAP7_75t_L g562 ( 
.A1(n_547),
.A2(n_508),
.A3(n_538),
.B1(n_424),
.B2(n_420),
.C1(n_494),
.C2(n_397),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_563),
.B(n_565),
.C(n_566),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_560),
.B(n_552),
.C(n_551),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_558),
.B(n_418),
.C(n_397),
.Y(n_566)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_569),
.Y(n_573)
);

AOI31xp33_ASAP7_75t_L g570 ( 
.A1(n_568),
.A2(n_559),
.A3(n_555),
.B(n_554),
.Y(n_570)
);

OAI321xp33_ASAP7_75t_L g575 ( 
.A1(n_570),
.A2(n_573),
.A3(n_567),
.B1(n_571),
.B2(n_420),
.C(n_411),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_564),
.Y(n_572)
);

AOI21x1_ASAP7_75t_L g574 ( 
.A1(n_572),
.A2(n_559),
.B(n_567),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_574),
.B(n_575),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_575),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_577),
.A2(n_576),
.B1(n_393),
.B2(n_309),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_393),
.Y(n_579)
);


endmodule