module fake_jpeg_15819_n_388 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_388);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_388;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_45),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g102 ( 
.A(n_46),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_67),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_63),
.B1(n_55),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_72),
.A2(n_84),
.B1(n_114),
.B2(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_14),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_77),
.B(n_80),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_90),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_37),
.B(n_35),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_101),
.Y(n_136)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_82),
.B(n_83),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_38),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_25),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_14),
.B1(n_19),
.B2(n_32),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_93),
.A2(n_117),
.B1(n_12),
.B2(n_13),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_35),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_96),
.A2(n_98),
.B(n_15),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_27),
.B(n_60),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_26),
.Y(n_99)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_45),
.A2(n_37),
.B(n_34),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_61),
.A2(n_34),
.B1(n_29),
.B2(n_24),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_30),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_29),
.B1(n_24),
.B2(n_16),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_24),
.B1(n_16),
.B2(n_32),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_20),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_113),
.Y(n_148)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_112),
.B(n_115),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_20),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_49),
.A2(n_26),
.B1(n_30),
.B2(n_15),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_39),
.A2(n_30),
.B1(n_15),
.B2(n_27),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_120),
.A2(n_135),
.B1(n_166),
.B2(n_131),
.Y(n_189)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_129),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_125),
.A2(n_87),
.B1(n_97),
.B2(n_91),
.Y(n_182)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_130),
.B(n_139),
.Y(n_188)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_88),
.Y(n_132)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_164),
.B(n_88),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_27),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_89),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_71),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_137),
.A2(n_138),
.B1(n_154),
.B2(n_167),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_71),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_2),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_140),
.A2(n_160),
.B(n_162),
.Y(n_181)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_145),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_27),
.B1(n_15),
.B2(n_7),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_103),
.B1(n_109),
.B2(n_104),
.Y(n_172)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_85),
.A2(n_15),
.B(n_27),
.C(n_7),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_146),
.B(n_91),
.Y(n_183)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_147),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_70),
.B(n_5),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_161),
.C(n_164),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_106),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_156),
.B1(n_112),
.B2(n_115),
.Y(n_178)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

BUFx4f_ASAP7_75t_SL g213 ( 
.A(n_153),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_157),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_95),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_96),
.B(n_10),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_107),
.B(n_13),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_13),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_163),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_76),
.A2(n_11),
.B(n_12),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_165),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_79),
.A2(n_13),
.B1(n_103),
.B2(n_102),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_168),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_169),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_172),
.A2(n_189),
.B1(n_171),
.B2(n_183),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_102),
.B(n_109),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_176),
.A2(n_183),
.B(n_186),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_177),
.A2(n_185),
.B(n_197),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_178),
.A2(n_208),
.B1(n_209),
.B2(n_212),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_182),
.A2(n_184),
.B1(n_207),
.B2(n_194),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_135),
.A2(n_87),
.B1(n_97),
.B2(n_73),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_122),
.B(n_89),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g187 ( 
.A(n_136),
.B(n_89),
.CI(n_148),
.CON(n_187),
.SN(n_187)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_187),
.B(n_201),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_192),
.B(n_186),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_136),
.A2(n_133),
.B(n_146),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_140),
.B(n_160),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_203),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_140),
.B(n_160),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_181),
.B(n_200),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_130),
.B(n_152),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_143),
.B(n_162),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_211),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_196),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_144),
.A2(n_120),
.B1(n_166),
.B2(n_147),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_121),
.A2(n_128),
.B1(n_123),
.B2(n_126),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_162),
.B(n_168),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_159),
.B(n_127),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_151),
.A2(n_141),
.B1(n_132),
.B2(n_153),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_163),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_213),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_219),
.A2(n_222),
.B1(n_245),
.B2(n_252),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_205),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_231),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_197),
.B1(n_172),
.B2(n_176),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_SL g264 ( 
.A(n_223),
.B(n_226),
.C(n_228),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_173),
.B(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_224),
.B(n_225),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_247),
.C(n_256),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_190),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_230),
.B(n_236),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_211),
.Y(n_231)
);

NAND2xp33_ASAP7_75t_SL g233 ( 
.A(n_177),
.B(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_233),
.Y(n_290)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_203),
.B(n_206),
.Y(n_236)
);

NOR2xp67_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_213),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_209),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_240),
.Y(n_262)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_188),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_186),
.B(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_178),
.B(n_199),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_246),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_179),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_193),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_180),
.B(n_216),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_180),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_249),
.A2(n_254),
.B(n_256),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_194),
.Y(n_250)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_216),
.B(n_204),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_207),
.A2(n_174),
.B1(n_202),
.B2(n_204),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_253),
.A2(n_239),
.B1(n_230),
.B2(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_175),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_251),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_258),
.B(n_272),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_261),
.B(n_287),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_175),
.B1(n_202),
.B2(n_174),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_266),
.A2(n_275),
.B1(n_279),
.B2(n_280),
.Y(n_301)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_242),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_227),
.Y(n_273)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_234),
.A2(n_243),
.B1(n_241),
.B2(n_219),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_222),
.A2(n_232),
.B1(n_220),
.B2(n_218),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_282),
.B1(n_231),
.B2(n_237),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_232),
.A2(n_220),
.B1(n_218),
.B2(n_254),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_285),
.A2(n_249),
.B(n_231),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_235),
.Y(n_287)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_244),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_225),
.B1(n_277),
.B2(n_284),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_226),
.C(n_247),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_292),
.C(n_302),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_229),
.C(n_233),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_221),
.Y(n_293)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_293),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_249),
.B1(n_245),
.B2(n_221),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_295),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_309),
.Y(n_325)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_297),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_298),
.B(n_312),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_299),
.A2(n_314),
.B(n_316),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_300),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_301),
.A2(n_277),
.B1(n_270),
.B2(n_268),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_282),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_273),
.Y(n_303)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_303),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_269),
.A2(n_263),
.B1(n_280),
.B2(n_279),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_306),
.A2(n_317),
.B1(n_293),
.B2(n_303),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_274),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_313),
.Y(n_331)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_285),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_264),
.B(n_259),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_310),
.B(n_291),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_278),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_263),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_290),
.A2(n_266),
.B(n_262),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_284),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_297),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_290),
.A2(n_260),
.B1(n_288),
.B2(n_276),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_307),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_332),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_260),
.B(n_283),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_319),
.A2(n_324),
.B(n_305),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_320),
.A2(n_321),
.B1(n_334),
.B2(n_323),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_306),
.A2(n_270),
.B1(n_268),
.B2(n_286),
.Y(n_321)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_314),
.A2(n_294),
.B(n_296),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_330),
.A2(n_338),
.B(n_309),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_308),
.Y(n_332)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_310),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_305),
.A2(n_292),
.B(n_317),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_302),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_347),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_340),
.A2(n_323),
.B(n_332),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_333),
.B(n_311),
.Y(n_342)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_344),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_348),
.C(n_350),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_313),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_304),
.C(n_311),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_324),
.B(n_304),
.Y(n_349)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_349),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_325),
.C(n_338),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_351),
.A2(n_327),
.B1(n_341),
.B2(n_355),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_334),
.C(n_319),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_352),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_322),
.C(n_326),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_353),
.B(n_354),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_321),
.C(n_329),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_320),
.B(n_318),
.C(n_335),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_355),
.B(n_339),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_353),
.Y(n_372)
);

MAJx2_ASAP7_75t_L g360 ( 
.A(n_347),
.B(n_335),
.C(n_327),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_360),
.A2(n_354),
.B(n_344),
.Y(n_371)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_363),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_365),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_366),
.B(n_350),
.C(n_348),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_358),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_368),
.B(n_372),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_369),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_371),
.B(n_373),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_359),
.A2(n_352),
.B(n_345),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_374),
.A2(n_365),
.B1(n_360),
.B2(n_361),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_377),
.B(n_361),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_368),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_380),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_378),
.A2(n_364),
.B(n_356),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_381),
.B(n_366),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_383),
.A2(n_375),
.B(n_370),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_384),
.A2(n_382),
.B(n_377),
.Y(n_385)
);

AO21x1_ASAP7_75t_L g386 ( 
.A1(n_385),
.A2(n_372),
.B(n_367),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_364),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_387),
.B(n_362),
.Y(n_388)
);


endmodule