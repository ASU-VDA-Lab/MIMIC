module fake_jpeg_19994_n_86 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_0),
.Y(n_57)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_40),
.B(n_37),
.C(n_42),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_38),
.B1(n_39),
.B2(n_2),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_59),
.B1(n_12),
.B2(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_3),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_15),
.B1(n_29),
.B2(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_1),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_14),
.C(n_24),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_13),
.B1(n_22),
.B2(n_4),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_77),
.B1(n_73),
.B2(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_78),
.A2(n_79),
.B1(n_54),
.B2(n_58),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_69),
.C(n_74),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_72),
.B(n_7),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_6),
.C(n_8),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_16),
.C(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_18),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_20),
.Y(n_86)
);


endmodule