module real_jpeg_384_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_206;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_30),
.B1(n_33),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_2),
.A2(n_39),
.B1(n_49),
.B2(n_50),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_2),
.B(n_24),
.C(n_26),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_2),
.B(n_22),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_2),
.A2(n_39),
.B1(n_63),
.B2(n_70),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_26),
.B1(n_28),
.B2(n_39),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_2),
.B(n_46),
.C(n_50),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_2),
.B(n_63),
.C(n_68),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_2),
.B(n_56),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_2),
.B(n_79),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_2),
.B(n_61),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_5),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_26),
.B1(n_28),
.B2(n_32),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_5),
.A2(n_32),
.B1(n_49),
.B2(n_50),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_5),
.A2(n_32),
.B1(n_63),
.B2(n_70),
.Y(n_174)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_8),
.A2(n_63),
.B1(n_70),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_10),
.A2(n_26),
.B1(n_28),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_10),
.A2(n_53),
.B1(n_63),
.B2(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_10),
.A2(n_30),
.B1(n_33),
.B2(n_53),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_125),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_124),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_102),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_16),
.B(n_102),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_76),
.C(n_89),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_17),
.A2(n_18),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_40),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_19),
.B(n_42),
.C(n_58),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_34),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_29),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_22),
.B(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_24),
.B1(n_30),
.B2(n_33),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_28),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_26),
.B(n_135),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_29),
.B(n_36),
.Y(n_113)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_30),
.B(n_86),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_58),
.B2(n_59),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_54),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_52),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_44),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_44),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_46),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_52),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_50),
.B1(n_67),
.B2(n_68),
.Y(n_73)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_50),
.B(n_166),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_55),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_56),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21x1_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_71),
.B(n_74),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_61),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_61),
.B(n_75),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_61),
.B(n_141),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_62)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_63),
.B(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_75),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_72),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_72),
.B(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_76),
.B(n_89),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_88),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B(n_82),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_84),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_78),
.A2(n_83),
.B(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_78),
.B(n_174),
.Y(n_188)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_79),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_80),
.A2(n_83),
.B(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_82),
.B(n_187),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_83),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.C(n_95),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_98),
.B(n_188),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_101),
.B(n_173),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_116),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_115),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_110),
.B2(n_114),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_108),
.B(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_110),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_153),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_140),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_145),
.B(n_206),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_142),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_127),
.B(n_142),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.C(n_137),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_129),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_137),
.B1(n_138),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21x1_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_160),
.B(n_205),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_158),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_203),
.Y(n_202)
);

OAI21x1_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_200),
.B(n_204),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_182),
.B(n_199),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_168),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_175),
.B1(n_176),
.B2(n_181),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_179),
.C(n_181),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_189),
.B(n_198),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_186),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_194),
.B(n_197),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_196),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_202),
.Y(n_204)
);


endmodule