module fake_netlist_6_3120_n_1239 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1239);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1239;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_1094;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_177;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_169;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_218;
wire n_1213;
wire n_172;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_653;
wire n_236;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_709;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_192;
wire n_649;

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_87),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_154),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_53),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_117),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_107),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_54),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_3),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_98),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_25),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_147),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_36),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_43),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_35),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_19),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_155),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_80),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_27),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_113),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_5),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_82),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_7),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_146),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_29),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_81),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_47),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_76),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_57),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_3),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_16),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_60),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_130),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_129),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_55),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_145),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_69),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_8),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_102),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_29),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_137),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_148),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_139),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_84),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_122),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_138),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_86),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_14),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_77),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_35),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_136),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_158),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_79),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_25),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_134),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_12),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_50),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_118),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_151),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_165),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_162),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_157),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_125),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_18),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_109),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_18),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_88),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_63),
.Y(n_242)
);

BUFx2_ASAP7_75t_SL g243 ( 
.A(n_92),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_160),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_78),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_64),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_140),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_164),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_142),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_75),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_32),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_23),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_114),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_52),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_141),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_166),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_156),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_135),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_89),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_39),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_2),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_10),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_58),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_15),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_93),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_143),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_74),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_62),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_42),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_149),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_41),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_133),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_132),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_1),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_12),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_23),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_38),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_11),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_16),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_150),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_13),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_101),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_33),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_52),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_59),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_27),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_163),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_20),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_2),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_152),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_214),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_176),
.B(n_0),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_178),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_229),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_180),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_224),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_229),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_249),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_228),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_252),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_249),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_268),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_268),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_175),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_181),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_190),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_276),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_213),
.B(n_0),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_176),
.B(n_1),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_216),
.B(n_4),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_193),
.Y(n_320)
);

INVxp33_ASAP7_75t_SL g321 ( 
.A(n_181),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_197),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_231),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_265),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_238),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_219),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_264),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_199),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_202),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_170),
.B(n_4),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_201),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_182),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_203),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_211),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_289),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_230),
.Y(n_340)
);

NOR2xp67_ASAP7_75t_L g341 ( 
.A(n_278),
.B(n_5),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_251),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_254),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_170),
.B(n_6),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_201),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_271),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_276),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_207),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_217),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_206),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_206),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_227),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_225),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_227),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_171),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_278),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_182),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_187),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_196),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_279),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_218),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_220),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_232),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_183),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_183),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_200),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_237),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_177),
.B(n_6),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_186),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_239),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_186),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_169),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_173),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_242),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_247),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_281),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_281),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_189),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_177),
.B(n_7),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_194),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_223),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_312),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

CKINVDCx11_ASAP7_75t_R g384 ( 
.A(n_296),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_312),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_314),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_168),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_319),
.B(n_174),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_381),
.Y(n_389)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_314),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_294),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_295),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_381),
.A2(n_285),
.B(n_223),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_303),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_306),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_308),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_310),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_317),
.B(n_200),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_358),
.B(n_168),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_350),
.B(n_285),
.Y(n_403)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_366),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_323),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_351),
.B(n_270),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_325),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_304),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_327),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_359),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_372),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_362),
.B(n_184),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_367),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_324),
.B(n_357),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_184),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_374),
.B(n_185),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_330),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_337),
.Y(n_421)
);

CKINVDCx8_ASAP7_75t_R g422 ( 
.A(n_365),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_352),
.B(n_272),
.Y(n_423)
);

BUFx8_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_339),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_354),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_368),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_356),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_356),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_364),
.B(n_179),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_333),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_373),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_345),
.B(n_185),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_344),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_379),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_291),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_301),
.Y(n_438)
);

AND2x2_ASAP7_75t_R g439 ( 
.A(n_321),
.B(n_222),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_369),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_315),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_292),
.B(n_280),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_347),
.B(n_282),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_318),
.Y(n_444)
);

INVx6_ASAP7_75t_L g445 ( 
.A(n_326),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_315),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_313),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_335),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_371),
.B(n_290),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_341),
.B(n_188),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_320),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_389),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_432),
.A2(n_435),
.B1(n_436),
.B2(n_427),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_419),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_388),
.B(n_321),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_388),
.B(n_378),
.Y(n_456)
);

OAI22xp33_ASAP7_75t_L g457 ( 
.A1(n_445),
.A2(n_261),
.B1(n_284),
.B2(n_286),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_426),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_322),
.C(n_320),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_426),
.Y(n_461)
);

BUFx8_ASAP7_75t_SL g462 ( 
.A(n_412),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_385),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_385),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_322),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_331),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_426),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_432),
.B(n_188),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_404),
.B(n_348),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_419),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_172),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_406),
.B(n_331),
.Y(n_473)
);

INVx4_ASAP7_75t_SL g474 ( 
.A(n_432),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_391),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_401),
.B(n_380),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_419),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_406),
.B(n_332),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_430),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_445),
.B(n_243),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_399),
.Y(n_483)
);

AO22x2_ASAP7_75t_L g484 ( 
.A1(n_401),
.A2(n_235),
.B1(n_198),
.B2(n_192),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_382),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_404),
.B(n_353),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_419),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_435),
.B(n_432),
.Y(n_488)
);

NOR2x1p5_ASAP7_75t_L g489 ( 
.A(n_441),
.B(n_293),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_406),
.B(n_423),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_389),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_419),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_411),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_432),
.A2(n_188),
.B1(n_191),
.B2(n_215),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_404),
.B(n_332),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_423),
.B(n_188),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_419),
.Y(n_499)
);

NOR2x1p5_ASAP7_75t_L g500 ( 
.A(n_441),
.B(n_293),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_435),
.B(n_336),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_411),
.Y(n_502)
);

BUFx10_ASAP7_75t_L g503 ( 
.A(n_431),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_389),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_404),
.B(n_336),
.Y(n_505)
);

BUFx6f_ASAP7_75t_SL g506 ( 
.A(n_446),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_389),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_435),
.B(n_338),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_389),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_411),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_445),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_445),
.B(n_338),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_435),
.B(n_340),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_435),
.B(n_340),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_414),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_414),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_404),
.B(n_342),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_435),
.B(n_342),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_389),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_432),
.B(n_343),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_432),
.B(n_343),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_445),
.Y(n_522)
);

NAND3xp33_ASAP7_75t_L g523 ( 
.A(n_455),
.B(n_416),
.C(n_451),
.Y(n_523)
);

INVxp33_ASAP7_75t_L g524 ( 
.A(n_465),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_478),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_503),
.B(n_441),
.Y(n_526)
);

NOR3xp33_ASAP7_75t_L g527 ( 
.A(n_456),
.B(n_441),
.C(n_451),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_503),
.B(n_441),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_466),
.B(n_408),
.Y(n_529)
);

AO221x1_ASAP7_75t_L g530 ( 
.A1(n_484),
.A2(n_446),
.B1(n_436),
.B2(n_444),
.C(n_215),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_483),
.Y(n_531)
);

INVx8_ASAP7_75t_L g532 ( 
.A(n_482),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_453),
.B(n_446),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_478),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_503),
.B(n_446),
.Y(n_535)
);

OAI22xp33_ASAP7_75t_L g536 ( 
.A1(n_501),
.A2(n_446),
.B1(n_445),
.B2(n_440),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_485),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_483),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_495),
.Y(n_539)
);

NOR3xp33_ASAP7_75t_L g540 ( 
.A(n_476),
.B(n_416),
.C(n_384),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_473),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_511),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_488),
.B(n_446),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_495),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_502),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_460),
.B(n_446),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_511),
.B(n_430),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_484),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_485),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_520),
.B(n_446),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_521),
.B(n_404),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_508),
.B(n_434),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_474),
.B(n_404),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_502),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_473),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_510),
.Y(n_556)
);

BUFx8_ASAP7_75t_L g557 ( 
.A(n_480),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_474),
.B(n_404),
.Y(n_558)
);

AOI221x1_ASAP7_75t_L g559 ( 
.A1(n_484),
.A2(n_442),
.B1(n_449),
.B2(n_402),
.C(n_413),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_474),
.B(n_440),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_490),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_522),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_474),
.B(n_440),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_513),
.B(n_434),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_462),
.B(n_422),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_510),
.Y(n_566)
);

NAND2x1_ASAP7_75t_L g567 ( 
.A(n_468),
.B(n_454),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_515),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_480),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_514),
.B(n_450),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_518),
.B(n_450),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_515),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_522),
.A2(n_387),
.B(n_402),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_490),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_516),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_491),
.B(n_450),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_489),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_512),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_516),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_491),
.B(n_390),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_481),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_491),
.B(n_447),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_491),
.B(n_311),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_498),
.B(n_387),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_484),
.A2(n_449),
.B1(n_448),
.B2(n_447),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_459),
.Y(n_586)
);

AND2x2_ASAP7_75t_SL g587 ( 
.A(n_472),
.B(n_191),
.Y(n_587)
);

NOR2x1p5_ASAP7_75t_L g588 ( 
.A(n_457),
.B(n_297),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_493),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_498),
.B(n_390),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_459),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_498),
.B(n_493),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_L g593 ( 
.A(n_472),
.B(n_448),
.C(n_360),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_463),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_498),
.B(n_390),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_496),
.B(n_442),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_458),
.B(n_390),
.Y(n_597)
);

O2A1O1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_497),
.A2(n_417),
.B(n_413),
.C(n_418),
.Y(n_598)
);

AO221x1_ASAP7_75t_L g599 ( 
.A1(n_452),
.A2(n_444),
.B1(n_191),
.B2(n_215),
.C(n_439),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_458),
.B(n_442),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_469),
.B(n_328),
.Y(n_601)
);

INVx8_ASAP7_75t_L g602 ( 
.A(n_482),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_461),
.B(n_390),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_L g604 ( 
.A1(n_482),
.A2(n_422),
.B1(n_418),
.B2(n_417),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_461),
.B(n_442),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_467),
.B(n_390),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_467),
.B(n_442),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_482),
.B(n_390),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_489),
.B(n_423),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_500),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_468),
.A2(n_410),
.B1(n_394),
.B2(n_383),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_468),
.A2(n_410),
.B1(n_394),
.B2(n_383),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_500),
.B(n_437),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_468),
.B(n_390),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_477),
.B(n_422),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_486),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_468),
.B(n_410),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_463),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_464),
.Y(n_619)
);

AO22x2_ASAP7_75t_L g620 ( 
.A1(n_505),
.A2(n_439),
.B1(n_273),
.B2(n_443),
.Y(n_620)
);

BUFx6f_ASAP7_75t_SL g621 ( 
.A(n_468),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_524),
.B(n_346),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_543),
.A2(n_470),
.B(n_454),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_582),
.B(n_517),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_529),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_550),
.A2(n_470),
.B(n_454),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_551),
.A2(n_471),
.B(n_464),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_539),
.Y(n_628)
);

NOR2x1_ASAP7_75t_R g629 ( 
.A(n_541),
.B(n_384),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_552),
.B(n_443),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_564),
.B(n_443),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_555),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_570),
.A2(n_487),
.B(n_470),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_533),
.A2(n_468),
.B(n_452),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_571),
.A2(n_612),
.B(n_611),
.Y(n_635)
);

AOI21x1_ASAP7_75t_L g636 ( 
.A1(n_551),
.A2(n_580),
.B(n_563),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_569),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_539),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_578),
.B(n_410),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_557),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_585),
.A2(n_403),
.B(n_438),
.C(n_437),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_576),
.A2(n_584),
.B(n_573),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_524),
.B(n_346),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_544),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_546),
.A2(n_305),
.B1(n_307),
.B2(n_309),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_557),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_544),
.Y(n_647)
);

AOI21x1_ASAP7_75t_L g648 ( 
.A1(n_580),
.A2(n_475),
.B(n_471),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_592),
.A2(n_492),
.B(n_452),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_598),
.A2(n_504),
.B(n_492),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_581),
.B(n_410),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_600),
.A2(n_487),
.B(n_477),
.Y(n_652)
);

AOI21x1_ASAP7_75t_L g653 ( 
.A1(n_560),
.A2(n_479),
.B(n_475),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_613),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_536),
.B(n_424),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_605),
.A2(n_504),
.B(n_492),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_547),
.B(n_383),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_532),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_547),
.B(n_383),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_607),
.A2(n_487),
.B(n_477),
.Y(n_660)
);

A2O1A1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_523),
.A2(n_403),
.B(n_438),
.C(n_437),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_590),
.A2(n_494),
.B(n_477),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_604),
.B(n_424),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_616),
.A2(n_506),
.B1(n_299),
.B2(n_300),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_545),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_547),
.B(n_525),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_577),
.B(n_405),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_545),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_609),
.B(n_405),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_590),
.A2(n_494),
.B(n_477),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_559),
.A2(n_509),
.B(n_504),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_554),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_527),
.B(n_360),
.C(n_424),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_534),
.B(n_509),
.Y(n_674)
);

O2A1O1Ixp5_ASAP7_75t_L g675 ( 
.A1(n_597),
.A2(n_519),
.B(n_509),
.C(n_479),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_532),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_554),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_526),
.B(n_408),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_535),
.A2(n_506),
.B1(n_412),
.B2(n_433),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_537),
.B(n_519),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_595),
.A2(n_499),
.B(n_494),
.Y(n_681)
);

O2A1O1Ixp33_ASAP7_75t_L g682 ( 
.A1(n_615),
.A2(n_403),
.B(n_415),
.C(n_407),
.Y(n_682)
);

AOI21x1_ASAP7_75t_L g683 ( 
.A1(n_560),
.A2(n_394),
.B(n_393),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_587),
.B(n_424),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_595),
.A2(n_499),
.B(n_494),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_549),
.B(n_561),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_528),
.B(n_297),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_556),
.Y(n_688)
);

NOR2xp67_ASAP7_75t_L g689 ( 
.A(n_593),
.B(n_610),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_562),
.Y(n_690)
);

OAI321xp33_ASAP7_75t_L g691 ( 
.A1(n_548),
.A2(n_428),
.A3(n_407),
.B1(n_415),
.B2(n_409),
.C(n_392),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_556),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_566),
.Y(n_693)
);

AO21x2_ASAP7_75t_L g694 ( 
.A1(n_530),
.A2(n_506),
.B(n_393),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_583),
.B(n_298),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_601),
.B(n_433),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_574),
.B(n_519),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_557),
.Y(n_698)
);

AOI33xp33_ASAP7_75t_L g699 ( 
.A1(n_589),
.A2(n_428),
.A3(n_409),
.B1(n_400),
.B2(n_421),
.B3(n_425),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_567),
.A2(n_499),
.B(n_494),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_597),
.A2(n_499),
.B(n_507),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_603),
.A2(n_499),
.B(n_507),
.Y(n_702)
);

OAI21xp33_ASAP7_75t_L g703 ( 
.A1(n_565),
.A2(n_376),
.B(n_365),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_587),
.B(n_424),
.Y(n_704)
);

CKINVDCx10_ASAP7_75t_R g705 ( 
.A(n_540),
.Y(n_705)
);

INVxp67_ASAP7_75t_R g706 ( 
.A(n_566),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_588),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_562),
.B(n_298),
.Y(n_708)
);

AOI21xp33_ASAP7_75t_L g709 ( 
.A1(n_620),
.A2(n_302),
.B(n_376),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_609),
.B(n_302),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_620),
.A2(n_609),
.B1(n_615),
.B2(n_599),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_568),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_617),
.B(n_191),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_532),
.A2(n_222),
.B1(n_269),
.B2(n_394),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_568),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_603),
.A2(n_606),
.B(n_608),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_606),
.A2(n_596),
.B(n_563),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_542),
.B(n_420),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_572),
.B(n_215),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_630),
.B(n_532),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_665),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_663),
.A2(n_579),
.B(n_572),
.C(n_575),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_631),
.B(n_620),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_654),
.B(n_602),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_625),
.B(n_678),
.Y(n_725)
);

BUFx12f_ASAP7_75t_L g726 ( 
.A(n_646),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_628),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_640),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_637),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_668),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_642),
.A2(n_635),
.B(n_626),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_623),
.A2(n_602),
.B(n_542),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_622),
.B(n_643),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_SL g734 ( 
.A(n_663),
.B(n_658),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_695),
.A2(n_602),
.B1(n_575),
.B2(n_579),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_687),
.A2(n_602),
.B(n_619),
.C(n_618),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_710),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_628),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_678),
.B(n_531),
.Y(n_739)
);

NAND2x1p5_ASAP7_75t_L g740 ( 
.A(n_676),
.B(n_542),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_632),
.B(n_377),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_637),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_667),
.Y(n_743)
);

AOI21x1_ASAP7_75t_L g744 ( 
.A1(n_713),
.A2(n_558),
.B(n_553),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_672),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_633),
.A2(n_542),
.B(n_553),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_709),
.A2(n_619),
.B(n_618),
.C(n_594),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_655),
.A2(n_269),
.B1(n_594),
.B2(n_531),
.Y(n_748)
);

A2O1A1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_687),
.A2(n_586),
.B(n_538),
.C(n_591),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_SL g750 ( 
.A(n_664),
.B(n_377),
.C(n_703),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_638),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_666),
.A2(n_591),
.B1(n_621),
.B2(n_558),
.Y(n_752)
);

AOI33xp33_ASAP7_75t_L g753 ( 
.A1(n_696),
.A2(n_667),
.A3(n_707),
.B1(n_645),
.B2(n_669),
.B3(n_698),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_655),
.A2(n_591),
.B1(n_621),
.B2(n_614),
.Y(n_754)
);

AO31x2_ASAP7_75t_L g755 ( 
.A1(n_641),
.A2(n_586),
.A3(n_538),
.B(n_414),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_622),
.B(n_233),
.Y(n_756)
);

OR2x6_ASAP7_75t_SL g757 ( 
.A(n_714),
.B(n_286),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_686),
.B(n_420),
.Y(n_758)
);

OAI21xp5_ASAP7_75t_L g759 ( 
.A1(n_717),
.A2(n_394),
.B(n_396),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_643),
.B(n_233),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_679),
.B(n_287),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_661),
.B(n_420),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_658),
.B(n_640),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_684),
.A2(n_172),
.B1(n_621),
.B2(n_263),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_661),
.B(n_421),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_638),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_676),
.B(n_507),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_R g768 ( 
.A(n_658),
.B(n_287),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_652),
.A2(n_507),
.B(n_419),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_669),
.Y(n_770)
);

NAND2x1p5_ASAP7_75t_L g771 ( 
.A(n_658),
.B(n_507),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_641),
.A2(n_421),
.B(n_425),
.C(n_395),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_708),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_639),
.B(n_425),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_705),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_SL g776 ( 
.A1(n_684),
.A2(n_395),
.B(n_398),
.C(n_392),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_718),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_695),
.B(n_706),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_690),
.B(n_288),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_689),
.B(n_400),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_677),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_SL g782 ( 
.A(n_704),
.B(n_195),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_671),
.A2(n_396),
.B(n_398),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_660),
.A2(n_507),
.B(n_389),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_656),
.A2(n_389),
.B(n_205),
.Y(n_785)
);

AO31x2_ASAP7_75t_L g786 ( 
.A1(n_731),
.A2(n_716),
.A3(n_693),
.B(n_712),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_778),
.B(n_711),
.Y(n_787)
);

BUFx12f_ASAP7_75t_L g788 ( 
.A(n_726),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_746),
.A2(n_627),
.B(n_648),
.Y(n_789)
);

AO31x2_ASAP7_75t_L g790 ( 
.A1(n_736),
.A2(n_749),
.A3(n_723),
.B(n_754),
.Y(n_790)
);

AO31x2_ASAP7_75t_L g791 ( 
.A1(n_762),
.A2(n_677),
.A3(n_693),
.B(n_715),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_732),
.A2(n_649),
.B(n_650),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_722),
.A2(n_634),
.B(n_713),
.Y(n_793)
);

NOR2xp67_ASAP7_75t_L g794 ( 
.A(n_773),
.B(n_673),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_727),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_739),
.B(n_690),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_759),
.A2(n_659),
.B(n_657),
.Y(n_797)
);

OAI21x1_ASAP7_75t_L g798 ( 
.A1(n_784),
.A2(n_653),
.B(n_636),
.Y(n_798)
);

O2A1O1Ixp5_ASAP7_75t_L g799 ( 
.A1(n_734),
.A2(n_719),
.B(n_675),
.C(n_624),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_721),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_737),
.B(n_691),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_733),
.B(n_624),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_774),
.A2(n_700),
.B(n_651),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_742),
.B(n_743),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_765),
.A2(n_783),
.B(n_747),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_725),
.B(n_741),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_772),
.A2(n_682),
.B(n_680),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_SL g808 ( 
.A1(n_720),
.A2(n_697),
.B(n_674),
.C(n_719),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_730),
.Y(n_809)
);

AOI21xp33_ASAP7_75t_L g810 ( 
.A1(n_748),
.A2(n_694),
.B(n_647),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_758),
.A2(n_718),
.B(n_670),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_785),
.A2(n_769),
.B(n_752),
.Y(n_812)
);

AOI21x1_ASAP7_75t_L g813 ( 
.A1(n_744),
.A2(n_683),
.B(n_681),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_725),
.B(n_692),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_728),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_770),
.B(n_644),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_740),
.A2(n_685),
.B(n_662),
.Y(n_817)
);

NOR2x1_ASAP7_75t_SL g818 ( 
.A(n_763),
.B(n_692),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_763),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_763),
.B(n_688),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_748),
.A2(n_715),
.B(n_712),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_729),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_735),
.A2(n_694),
.B(n_701),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_738),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_780),
.Y(n_825)
);

AO32x2_ASAP7_75t_L g826 ( 
.A1(n_755),
.A2(n_699),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_764),
.A2(n_702),
.B(n_699),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_751),
.B(n_399),
.Y(n_828)
);

AO31x2_ASAP7_75t_L g829 ( 
.A1(n_766),
.A2(n_399),
.A3(n_172),
.B(n_246),
.Y(n_829)
);

CKINVDCx8_ASAP7_75t_R g830 ( 
.A(n_780),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_768),
.Y(n_831)
);

AND2x6_ASAP7_75t_L g832 ( 
.A(n_781),
.B(n_629),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_SL g833 ( 
.A1(n_761),
.A2(n_396),
.B(n_172),
.C(n_200),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_741),
.B(n_770),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_776),
.A2(n_764),
.B(n_782),
.Y(n_835)
);

AO31x2_ASAP7_75t_L g836 ( 
.A1(n_745),
.A2(n_779),
.A3(n_755),
.B(n_757),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_729),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_755),
.Y(n_838)
);

AOI21x1_ASAP7_75t_L g839 ( 
.A1(n_724),
.A2(n_397),
.B(n_396),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_740),
.A2(n_396),
.B(n_172),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_806),
.A2(n_756),
.B1(n_760),
.B2(n_779),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_800),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_809),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_795),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_814),
.B(n_777),
.Y(n_845)
);

BUFx12f_ASAP7_75t_L g846 ( 
.A(n_788),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_824),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_837),
.Y(n_848)
);

INVx6_ASAP7_75t_L g849 ( 
.A(n_819),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_787),
.A2(n_288),
.B1(n_246),
.B2(n_263),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_801),
.A2(n_750),
.B1(n_753),
.B2(n_771),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_816),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_819),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_828),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_797),
.A2(n_750),
.B(n_771),
.Y(n_855)
);

INVx6_ASAP7_75t_L g856 ( 
.A(n_819),
.Y(n_856)
);

NAND2x1p5_ASAP7_75t_L g857 ( 
.A(n_820),
.B(n_429),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_802),
.A2(n_246),
.B1(n_253),
.B2(n_263),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_815),
.Y(n_859)
);

OAI22xp33_ASAP7_75t_L g860 ( 
.A1(n_802),
.A2(n_775),
.B1(n_429),
.B2(n_768),
.Y(n_860)
);

BUFx2_ASAP7_75t_SL g861 ( 
.A(n_830),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_825),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_786),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_834),
.A2(n_253),
.B1(n_172),
.B2(n_429),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_828),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_814),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_SL g867 ( 
.A1(n_831),
.A2(n_253),
.B(n_767),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_822),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_804),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_825),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_796),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_796),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_829),
.Y(n_873)
);

INVx8_ASAP7_75t_L g874 ( 
.A(n_820),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_794),
.A2(n_767),
.B1(n_248),
.B2(n_245),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_SL g876 ( 
.A1(n_805),
.A2(n_825),
.B1(n_818),
.B2(n_792),
.Y(n_876)
);

INVx6_ASAP7_75t_L g877 ( 
.A(n_832),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_SL g878 ( 
.A1(n_805),
.A2(n_172),
.B1(n_204),
.B2(n_208),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_832),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_810),
.A2(n_429),
.B1(n_210),
.B2(n_212),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_SL g881 ( 
.A1(n_832),
.A2(n_209),
.B1(n_221),
.B2(n_226),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_832),
.Y(n_882)
);

INVx6_ASAP7_75t_L g883 ( 
.A(n_836),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_836),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_810),
.A2(n_429),
.B1(n_236),
.B2(n_241),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_821),
.B(n_429),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_821),
.A2(n_429),
.B1(n_244),
.B2(n_250),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_835),
.Y(n_888)
);

INVx6_ASAP7_75t_L g889 ( 
.A(n_836),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_829),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_835),
.A2(n_259),
.B1(n_255),
.B2(n_256),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_829),
.B(n_429),
.Y(n_892)
);

INVx3_ASAP7_75t_SL g893 ( 
.A(n_838),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_823),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_840),
.Y(n_895)
);

INVx6_ASAP7_75t_L g896 ( 
.A(n_799),
.Y(n_896)
);

BUFx12f_ASAP7_75t_L g897 ( 
.A(n_833),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_807),
.A2(n_267),
.B1(n_266),
.B2(n_258),
.Y(n_898)
);

BUFx12f_ASAP7_75t_L g899 ( 
.A(n_826),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_893),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_873),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_884),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_894),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_890),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_863),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_871),
.B(n_791),
.Y(n_906)
);

OAI21x1_ASAP7_75t_SL g907 ( 
.A1(n_855),
.A2(n_823),
.B(n_797),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_895),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_893),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_883),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_888),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_899),
.B(n_826),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_883),
.B(n_826),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_896),
.B(n_812),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_883),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_889),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_889),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_841),
.A2(n_807),
.B1(n_827),
.B2(n_234),
.Y(n_918)
);

OA21x2_ASAP7_75t_L g919 ( 
.A1(n_886),
.A2(n_793),
.B(n_798),
.Y(n_919)
);

AOI21x1_ASAP7_75t_L g920 ( 
.A1(n_892),
.A2(n_793),
.B(n_813),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_889),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_872),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_896),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_896),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_842),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_874),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_843),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_874),
.Y(n_928)
);

OR2x6_ASAP7_75t_L g929 ( 
.A(n_874),
.B(n_811),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_866),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_882),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_854),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_845),
.B(n_791),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_848),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_865),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_844),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_897),
.B(n_811),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_841),
.B(n_808),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_931),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_913),
.B(n_876),
.Y(n_940)
);

AND2x4_ASAP7_75t_SL g941 ( 
.A(n_923),
.B(n_853),
.Y(n_941)
);

NAND2xp33_ASAP7_75t_L g942 ( 
.A(n_918),
.B(n_850),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_918),
.A2(n_938),
.B(n_878),
.C(n_911),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_925),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_911),
.B(n_868),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_935),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_908),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_930),
.B(n_869),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_911),
.B(n_852),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_911),
.A2(n_850),
.B1(n_858),
.B2(n_881),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_930),
.B(n_847),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_931),
.B(n_876),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_931),
.B(n_879),
.Y(n_953)
);

NAND2x1_ASAP7_75t_L g954 ( 
.A(n_924),
.B(n_877),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_913),
.B(n_790),
.Y(n_955)
);

BUFx10_ASAP7_75t_L g956 ( 
.A(n_900),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_925),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_938),
.A2(n_860),
.B(n_851),
.C(n_867),
.Y(n_958)
);

AO32x2_ASAP7_75t_L g959 ( 
.A1(n_900),
.A2(n_875),
.A3(n_878),
.B1(n_790),
.B2(n_860),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_916),
.B(n_853),
.Y(n_960)
);

AO32x2_ASAP7_75t_L g961 ( 
.A1(n_900),
.A2(n_790),
.A3(n_791),
.B1(n_885),
.B2(n_880),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_931),
.Y(n_962)
);

OR2x6_ASAP7_75t_L g963 ( 
.A(n_929),
.B(n_877),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_903),
.B(n_922),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_909),
.Y(n_965)
);

NAND4xp25_ASAP7_75t_L g966 ( 
.A(n_934),
.B(n_858),
.C(n_881),
.D(n_898),
.Y(n_966)
);

AO21x2_ASAP7_75t_L g967 ( 
.A1(n_907),
.A2(n_891),
.B(n_827),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_SL g968 ( 
.A1(n_909),
.A2(n_870),
.B(n_877),
.C(n_864),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_909),
.Y(n_969)
);

NOR2xp67_ASAP7_75t_SL g970 ( 
.A(n_923),
.B(n_861),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_924),
.B(n_859),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_916),
.B(n_853),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_908),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_924),
.B(n_849),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_925),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_926),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_927),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_924),
.B(n_849),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_916),
.B(n_862),
.Y(n_979)
);

INVxp67_ASAP7_75t_SL g980 ( 
.A(n_964),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_977),
.B(n_903),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_946),
.B(n_933),
.Y(n_982)
);

INVx5_ASAP7_75t_L g983 ( 
.A(n_963),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_955),
.B(n_913),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_946),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_944),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_963),
.B(n_910),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_942),
.A2(n_912),
.B1(n_937),
.B2(n_907),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_958),
.B(n_928),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_942),
.A2(n_912),
.B1(n_880),
.B2(n_885),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_955),
.B(n_919),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_957),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_975),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_951),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_947),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_940),
.B(n_902),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_947),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_947),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_940),
.B(n_919),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_963),
.B(n_919),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_963),
.B(n_919),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_939),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_954),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_973),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_973),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_SL g1006 ( 
.A1(n_990),
.A2(n_950),
.B(n_943),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_999),
.B(n_973),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_999),
.B(n_984),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_985),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_999),
.B(n_952),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_984),
.B(n_991),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_991),
.B(n_1000),
.Y(n_1012)
);

OAI221xp5_ASAP7_75t_SL g1013 ( 
.A1(n_990),
.A2(n_943),
.B1(n_966),
.B2(n_912),
.C(n_864),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_986),
.Y(n_1014)
);

AOI221xp5_ASAP7_75t_SL g1015 ( 
.A1(n_988),
.A2(n_934),
.B1(n_949),
.B2(n_948),
.C(n_971),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_986),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_992),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_992),
.Y(n_1018)
);

AOI31xp33_ASAP7_75t_L g1019 ( 
.A1(n_989),
.A2(n_945),
.A3(n_965),
.B(n_969),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_984),
.B(n_939),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_985),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_985),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_993),
.Y(n_1023)
);

AOI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_980),
.A2(n_907),
.B(n_967),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_993),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_994),
.B(n_965),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_996),
.A2(n_962),
.B1(n_887),
.B2(n_976),
.Y(n_1027)
);

NOR2x1_ASAP7_75t_L g1028 ( 
.A(n_1019),
.B(n_1006),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1014),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1008),
.B(n_983),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1014),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1022),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1016),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1008),
.B(n_983),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1011),
.B(n_983),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1011),
.B(n_983),
.Y(n_1036)
);

NAND2x1_ASAP7_75t_SL g1037 ( 
.A(n_1009),
.B(n_1021),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1012),
.B(n_983),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1016),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1029),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_1037),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_1037),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1038),
.B(n_1010),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_1029),
.B(n_996),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_1038),
.B(n_1012),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1032),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1040),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1043),
.B(n_1030),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1045),
.B(n_1028),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_1041),
.Y(n_1050)
);

OAI32xp33_ASAP7_75t_L g1051 ( 
.A1(n_1049),
.A2(n_1042),
.A3(n_1041),
.B1(n_1006),
.B2(n_1027),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1050),
.A2(n_1027),
.B1(n_1015),
.B2(n_1042),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1047),
.B(n_1048),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1048),
.Y(n_1054)
);

AOI322xp5_ASAP7_75t_L g1055 ( 
.A1(n_1049),
.A2(n_1015),
.A3(n_1045),
.B1(n_1012),
.B2(n_1030),
.C1(n_1036),
.C2(n_1035),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_1048),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1048),
.B(n_1045),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1047),
.B(n_1031),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1048),
.B(n_1034),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1048),
.B(n_1034),
.Y(n_1060)
);

OAI211xp5_ASAP7_75t_L g1061 ( 
.A1(n_1049),
.A2(n_1013),
.B(n_1024),
.C(n_968),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1056),
.B(n_1044),
.Y(n_1062)
);

AOI32xp33_ASAP7_75t_L g1063 ( 
.A1(n_1056),
.A2(n_1036),
.A3(n_1035),
.B1(n_1026),
.B2(n_1013),
.Y(n_1063)
);

O2A1O1Ixp5_ASAP7_75t_L g1064 ( 
.A1(n_1051),
.A2(n_1046),
.B(n_1024),
.C(n_980),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1053),
.Y(n_1065)
);

OAI32xp33_ASAP7_75t_L g1066 ( 
.A1(n_1053),
.A2(n_1046),
.A3(n_996),
.B1(n_1032),
.B2(n_1003),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1057),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1061),
.A2(n_1019),
.B(n_968),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1058),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1058),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1054),
.B(n_1010),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_1052),
.A2(n_1003),
.B(n_1033),
.C(n_1031),
.Y(n_1072)
);

OAI322xp33_ASAP7_75t_L g1073 ( 
.A1(n_1055),
.A2(n_1039),
.A3(n_1033),
.B1(n_981),
.B2(n_1023),
.C1(n_1018),
.C2(n_1017),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_1059),
.B(n_1039),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1060),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_L g1076 ( 
.A(n_1055),
.B(n_970),
.C(n_969),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1056),
.B(n_1007),
.Y(n_1077)
);

CKINVDCx14_ASAP7_75t_R g1078 ( 
.A(n_1067),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1075),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1071),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_1065),
.B(n_846),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1069),
.B(n_1017),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1062),
.B(n_1018),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_1070),
.B(n_1020),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1063),
.B(n_1023),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1072),
.B(n_1007),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1074),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1077),
.Y(n_1088)
);

OAI221xp5_ASAP7_75t_SL g1089 ( 
.A1(n_1076),
.A2(n_937),
.B1(n_1003),
.B2(n_914),
.C(n_887),
.Y(n_1089)
);

XNOR2x1_ASAP7_75t_L g1090 ( 
.A(n_1068),
.B(n_8),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1064),
.A2(n_978),
.B(n_981),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1066),
.B(n_1025),
.Y(n_1092)
);

OAI22xp33_ASAP7_75t_SL g1093 ( 
.A1(n_1073),
.A2(n_983),
.B1(n_1025),
.B2(n_1022),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1073),
.Y(n_1094)
);

AOI221xp5_ASAP7_75t_L g1095 ( 
.A1(n_1073),
.A2(n_994),
.B1(n_997),
.B2(n_998),
.C(n_1005),
.Y(n_1095)
);

OAI21xp33_ASAP7_75t_SL g1096 ( 
.A1(n_1063),
.A2(n_1020),
.B(n_1009),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1087),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1079),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1078),
.B(n_1022),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1090),
.B(n_1022),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1094),
.B(n_1021),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1082),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1080),
.B(n_997),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1081),
.A2(n_976),
.B1(n_962),
.B2(n_1002),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1088),
.Y(n_1105)
);

BUFx4f_ASAP7_75t_SL g1106 ( 
.A(n_1084),
.Y(n_1106)
);

NAND4xp25_ASAP7_75t_L g1107 ( 
.A(n_1089),
.B(n_953),
.C(n_974),
.D(n_928),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1084),
.B(n_998),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1096),
.B(n_1085),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_1083),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_SL g1111 ( 
.A(n_1095),
.B(n_257),
.C(n_9),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1086),
.A2(n_983),
.B1(n_967),
.B2(n_937),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1096),
.B(n_1092),
.Y(n_1113)
);

AOI221xp5_ASAP7_75t_L g1114 ( 
.A1(n_1113),
.A2(n_1093),
.B1(n_1091),
.B2(n_1002),
.C(n_1004),
.Y(n_1114)
);

AOI221x1_ASAP7_75t_L g1115 ( 
.A1(n_1098),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C(n_17),
.Y(n_1115)
);

AOI211xp5_ASAP7_75t_L g1116 ( 
.A1(n_1109),
.A2(n_862),
.B(n_19),
.C(n_20),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1097),
.B(n_1004),
.Y(n_1117)
);

NAND4xp75_ASAP7_75t_L g1118 ( 
.A(n_1105),
.B(n_17),
.C(n_21),
.D(n_22),
.Y(n_1118)
);

AOI221xp5_ASAP7_75t_L g1119 ( 
.A1(n_1111),
.A2(n_1005),
.B1(n_927),
.B2(n_1000),
.C(n_1001),
.Y(n_1119)
);

AOI21xp33_ASAP7_75t_L g1120 ( 
.A1(n_1110),
.A2(n_21),
.B(n_22),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_SL g1121 ( 
.A1(n_1099),
.A2(n_926),
.B(n_26),
.C(n_28),
.Y(n_1121)
);

OAI211xp5_ASAP7_75t_L g1122 ( 
.A1(n_1101),
.A2(n_1111),
.B(n_1100),
.C(n_1107),
.Y(n_1122)
);

OAI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1106),
.A2(n_937),
.B1(n_914),
.B2(n_929),
.Y(n_1123)
);

OAI222xp33_ASAP7_75t_L g1124 ( 
.A1(n_1104),
.A2(n_937),
.B1(n_914),
.B2(n_929),
.C1(n_960),
.C2(n_972),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_1102),
.A2(n_1103),
.B(n_1108),
.C(n_1112),
.Y(n_1125)
);

NOR2x1_ASAP7_75t_L g1126 ( 
.A(n_1097),
.B(n_24),
.Y(n_1126)
);

O2A1O1Ixp5_ASAP7_75t_L g1127 ( 
.A1(n_1113),
.A2(n_995),
.B(n_936),
.C(n_960),
.Y(n_1127)
);

NAND4xp25_ASAP7_75t_L g1128 ( 
.A(n_1109),
.B(n_928),
.C(n_1001),
.D(n_1000),
.Y(n_1128)
);

AOI221xp5_ASAP7_75t_L g1129 ( 
.A1(n_1113),
.A2(n_1001),
.B1(n_995),
.B2(n_982),
.C(n_922),
.Y(n_1129)
);

NOR4xp25_ASAP7_75t_L g1130 ( 
.A(n_1097),
.B(n_24),
.C(n_26),
.D(n_28),
.Y(n_1130)
);

AOI21xp33_ASAP7_75t_L g1131 ( 
.A1(n_1109),
.A2(n_30),
.B(n_31),
.Y(n_1131)
);

OAI221xp5_ASAP7_75t_SL g1132 ( 
.A1(n_1109),
.A2(n_937),
.B1(n_914),
.B2(n_929),
.C(n_926),
.Y(n_1132)
);

AOI221xp5_ASAP7_75t_L g1133 ( 
.A1(n_1113),
.A2(n_995),
.B1(n_982),
.B2(n_972),
.C(n_960),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1098),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1097),
.Y(n_1135)
);

NAND4xp75_ASAP7_75t_L g1136 ( 
.A(n_1097),
.B(n_33),
.C(n_34),
.D(n_36),
.Y(n_1136)
);

OAI211xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1109),
.A2(n_34),
.B(n_37),
.C(n_38),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1130),
.B(n_37),
.Y(n_1138)
);

AOI221xp5_ASAP7_75t_L g1139 ( 
.A1(n_1131),
.A2(n_862),
.B1(n_972),
.B2(n_41),
.C(n_42),
.Y(n_1139)
);

NOR3xp33_ASAP7_75t_L g1140 ( 
.A(n_1137),
.B(n_928),
.C(n_40),
.Y(n_1140)
);

AOI221xp5_ASAP7_75t_L g1141 ( 
.A1(n_1125),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.C(n_44),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1122),
.A2(n_849),
.B1(n_856),
.B2(n_979),
.Y(n_1142)
);

AOI211xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1116),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1126),
.B(n_45),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1135),
.B(n_987),
.Y(n_1145)
);

AOI222xp33_ASAP7_75t_L g1146 ( 
.A1(n_1119),
.A2(n_956),
.B1(n_47),
.B2(n_48),
.C1(n_49),
.C2(n_50),
.Y(n_1146)
);

NAND4xp25_ASAP7_75t_L g1147 ( 
.A(n_1133),
.B(n_928),
.C(n_979),
.D(n_987),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1136),
.Y(n_1148)
);

AOI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_1114),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.C(n_51),
.Y(n_1149)
);

NAND3xp33_ASAP7_75t_L g1150 ( 
.A(n_1115),
.B(n_51),
.C(n_937),
.Y(n_1150)
);

OAI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_1128),
.A2(n_941),
.B(n_979),
.Y(n_1151)
);

AOI211xp5_ASAP7_75t_L g1152 ( 
.A1(n_1121),
.A2(n_933),
.B(n_991),
.C(n_987),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1118),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1134),
.A2(n_932),
.B1(n_921),
.B2(n_936),
.C(n_917),
.Y(n_1154)
);

AOI222xp33_ASAP7_75t_L g1155 ( 
.A1(n_1129),
.A2(n_1117),
.B1(n_1124),
.B2(n_1123),
.C1(n_1127),
.C2(n_1134),
.Y(n_1155)
);

NAND4xp25_ASAP7_75t_SL g1156 ( 
.A(n_1120),
.B(n_921),
.C(n_917),
.D(n_932),
.Y(n_1156)
);

AOI221xp5_ASAP7_75t_L g1157 ( 
.A1(n_1132),
.A2(n_941),
.B1(n_936),
.B2(n_987),
.C(n_985),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1137),
.A2(n_856),
.B1(n_956),
.B2(n_914),
.Y(n_1158)
);

OAI211xp5_ASAP7_75t_SL g1159 ( 
.A1(n_1122),
.A2(n_936),
.B(n_908),
.C(n_803),
.Y(n_1159)
);

AOI211xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1131),
.A2(n_908),
.B(n_917),
.C(n_987),
.Y(n_1160)
);

OAI221xp5_ASAP7_75t_L g1161 ( 
.A1(n_1137),
.A2(n_856),
.B1(n_914),
.B2(n_929),
.C(n_908),
.Y(n_1161)
);

XNOR2x1_ASAP7_75t_L g1162 ( 
.A(n_1153),
.B(n_56),
.Y(n_1162)
);

XNOR2x1_ASAP7_75t_L g1163 ( 
.A(n_1148),
.B(n_61),
.Y(n_1163)
);

NOR2x1_ASAP7_75t_L g1164 ( 
.A(n_1144),
.B(n_65),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1138),
.Y(n_1165)
);

AOI221xp5_ASAP7_75t_SL g1166 ( 
.A1(n_1141),
.A2(n_904),
.B1(n_901),
.B2(n_902),
.C(n_906),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1150),
.B(n_935),
.Y(n_1167)
);

NOR2x1_ASAP7_75t_L g1168 ( 
.A(n_1156),
.B(n_66),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1145),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1142),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1140),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1139),
.Y(n_1172)
);

NOR2x1_ASAP7_75t_L g1173 ( 
.A(n_1159),
.B(n_67),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1143),
.B(n_956),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1149),
.A2(n_857),
.B(n_914),
.C(n_929),
.Y(n_1175)
);

NAND2xp33_ASAP7_75t_L g1176 ( 
.A(n_1158),
.B(n_857),
.Y(n_1176)
);

NOR2xp67_ASAP7_75t_L g1177 ( 
.A(n_1161),
.B(n_68),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1155),
.Y(n_1178)
);

NOR2x1_ASAP7_75t_L g1179 ( 
.A(n_1147),
.B(n_70),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1154),
.B(n_935),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1152),
.Y(n_1181)
);

XOR2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1146),
.B(n_959),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1151),
.B(n_72),
.Y(n_1183)
);

OAI322xp33_ASAP7_75t_L g1184 ( 
.A1(n_1178),
.A2(n_1160),
.A3(n_1157),
.B1(n_901),
.B2(n_904),
.C1(n_906),
.C2(n_959),
.Y(n_1184)
);

NAND4xp75_ASAP7_75t_L g1185 ( 
.A(n_1164),
.B(n_73),
.C(n_83),
.D(n_85),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1169),
.B(n_1170),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1163),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1174),
.B(n_935),
.Y(n_1188)
);

OAI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1171),
.A2(n_1181),
.B1(n_1172),
.B2(n_1165),
.C(n_1183),
.Y(n_1189)
);

AOI211xp5_ASAP7_75t_L g1190 ( 
.A1(n_1177),
.A2(n_915),
.B(n_910),
.C(n_817),
.Y(n_1190)
);

OAI211xp5_ASAP7_75t_L g1191 ( 
.A1(n_1173),
.A2(n_839),
.B(n_916),
.C(n_902),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1162),
.B(n_1168),
.Y(n_1192)
);

NOR3xp33_ASAP7_75t_L g1193 ( 
.A(n_1179),
.B(n_916),
.C(n_920),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1167),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1173),
.B(n_1166),
.Y(n_1195)
);

NOR3xp33_ASAP7_75t_L g1196 ( 
.A(n_1175),
.B(n_920),
.C(n_915),
.Y(n_1196)
);

OAI221xp5_ASAP7_75t_L g1197 ( 
.A1(n_1176),
.A2(n_929),
.B1(n_915),
.B2(n_910),
.C(n_959),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_SL g1198 ( 
.A1(n_1180),
.A2(n_90),
.B(n_91),
.C(n_94),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1186),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1186),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1192),
.A2(n_1182),
.B1(n_910),
.B2(n_915),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_L g1202 ( 
.A(n_1189),
.B(n_397),
.C(n_96),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1194),
.Y(n_1203)
);

AOI222xp33_ASAP7_75t_L g1204 ( 
.A1(n_1195),
.A2(n_1187),
.B1(n_1188),
.B2(n_1191),
.C1(n_1198),
.C2(n_1197),
.Y(n_1204)
);

OAI211xp5_ASAP7_75t_L g1205 ( 
.A1(n_1190),
.A2(n_95),
.B(n_97),
.C(n_99),
.Y(n_1205)
);

NAND2x1_ASAP7_75t_L g1206 ( 
.A(n_1193),
.B(n_397),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1185),
.Y(n_1207)
);

NAND2x1_ASAP7_75t_L g1208 ( 
.A(n_1196),
.B(n_397),
.Y(n_1208)
);

NAND4xp25_ASAP7_75t_L g1209 ( 
.A(n_1184),
.B(n_100),
.C(n_103),
.D(n_104),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1186),
.B(n_106),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_SL g1211 ( 
.A1(n_1192),
.A2(n_959),
.B(n_920),
.Y(n_1211)
);

NAND2x1p5_ASAP7_75t_SL g1212 ( 
.A(n_1187),
.B(n_108),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1192),
.A2(n_397),
.B(n_789),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1199),
.Y(n_1214)
);

BUFx8_ASAP7_75t_L g1215 ( 
.A(n_1200),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1201),
.A2(n_919),
.B1(n_905),
.B2(n_397),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_SL g1217 ( 
.A1(n_1207),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1210),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1203),
.A2(n_919),
.B1(n_905),
.B2(n_397),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1209),
.A2(n_1204),
.B1(n_1202),
.B2(n_1205),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1206),
.A2(n_905),
.B1(n_961),
.B2(n_119),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1212),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1208),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_SL g1224 ( 
.A(n_1214),
.B(n_1213),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1215),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1222),
.Y(n_1226)
);

OAI22x1_ASAP7_75t_L g1227 ( 
.A1(n_1220),
.A2(n_1211),
.B1(n_116),
.B2(n_120),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_SL g1228 ( 
.A1(n_1218),
.A2(n_1217),
.B1(n_1223),
.B2(n_1221),
.Y(n_1228)
);

XOR2xp5_ASAP7_75t_L g1229 ( 
.A(n_1216),
.B(n_115),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1225),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1227),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1226),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1228),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1230),
.A2(n_1224),
.B(n_1229),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1234),
.Y(n_1235)
);

AOI21xp33_ASAP7_75t_L g1236 ( 
.A1(n_1235),
.A2(n_1233),
.B(n_1232),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1236),
.Y(n_1237)
);

OAI221xp5_ASAP7_75t_R g1238 ( 
.A1(n_1237),
.A2(n_1231),
.B1(n_1219),
.B2(n_126),
.C(n_127),
.Y(n_1238)
);

AOI211xp5_ASAP7_75t_L g1239 ( 
.A1(n_1238),
.A2(n_123),
.B(n_124),
.C(n_128),
.Y(n_1239)
);


endmodule