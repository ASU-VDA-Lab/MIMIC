module fake_jpeg_23755_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_9),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx9p33_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_52),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_28),
.B1(n_19),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_55),
.B1(n_25),
.B2(n_22),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_25),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_54),
.B(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_19),
.B1(n_22),
.B2(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_25),
.B1(n_18),
.B2(n_30),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_30),
.B1(n_23),
.B2(n_18),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_70),
.B1(n_46),
.B2(n_27),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_68),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_84),
.B1(n_59),
.B2(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_30),
.B1(n_23),
.B2(n_18),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_27),
.B(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_22),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_44),
.A2(n_22),
.B1(n_31),
.B2(n_29),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_101)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_81),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_43),
.B1(n_45),
.B2(n_44),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_52),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_43),
.B1(n_45),
.B2(n_52),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_100),
.B1(n_104),
.B2(n_109),
.Y(n_114)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_49),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_95),
.B(n_103),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_101),
.B1(n_107),
.B2(n_83),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_49),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_49),
.B1(n_46),
.B2(n_53),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_27),
.B(n_16),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_67),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_110),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_61),
.A2(n_53),
.B1(n_16),
.B2(n_32),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_0),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_62),
.B1(n_60),
.B2(n_75),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_113),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_117),
.A2(n_110),
.B1(n_114),
.B2(n_88),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_69),
.B1(n_68),
.B2(n_71),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_99),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_71),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_125),
.B1(n_127),
.B2(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_131),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_74),
.B1(n_79),
.B2(n_57),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_74),
.B1(n_79),
.B2(n_57),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_39),
.B1(n_38),
.B2(n_20),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_21),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_28),
.B1(n_32),
.B2(n_21),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_57),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_57),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_20),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_95),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_157),
.C(n_158),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_149),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_86),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_146),
.A2(n_154),
.B(n_162),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_155),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_98),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_28),
.B1(n_10),
.B2(n_3),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_130),
.B(n_118),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_97),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_57),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_103),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_88),
.C(n_97),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_104),
.C(n_109),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_161),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_110),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_112),
.A2(n_102),
.B(n_101),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_112),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_173),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_124),
.C(n_133),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_156),
.C(n_138),
.Y(n_195)
);

OAI322xp33_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_115),
.A3(n_114),
.B1(n_132),
.B2(n_123),
.C1(n_21),
.C2(n_26),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_177),
.B(n_139),
.Y(n_191)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_115),
.B1(n_102),
.B2(n_57),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_177),
.B1(n_185),
.B2(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_179),
.Y(n_190)
);

OAI22x1_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_26),
.B1(n_0),
.B2(n_2),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

AOI322xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_182),
.A3(n_138),
.B1(n_151),
.B2(n_6),
.C1(n_8),
.C2(n_10),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_8),
.A3(n_14),
.B1(n_3),
.B2(n_4),
.C1(n_6),
.C2(n_7),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_145),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_140),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_154),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_187),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_181),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_189),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_168),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_141),
.C(n_149),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_199),
.C(n_172),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_167),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_196),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_201),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

AOI321xp33_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_161),
.A3(n_158),
.B1(n_163),
.B2(n_146),
.C(n_159),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_164),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_160),
.C(n_145),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_202),
.A2(n_204),
.B1(n_166),
.B2(n_185),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_183),
.B(n_11),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_176),
.C(n_184),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_208),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_210),
.C(n_216),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_199),
.C(n_187),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_172),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_215),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_175),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_173),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_217),
.A2(n_204),
.B1(n_202),
.B2(n_200),
.Y(n_219)
);

O2A1O1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_219),
.A2(n_222),
.B(n_225),
.C(n_224),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_213),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_12),
.C(n_13),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_218),
.A2(n_200),
.B1(n_193),
.B2(n_194),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_216),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_227),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_217),
.A2(n_196),
.B1(n_189),
.B2(n_190),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_12),
.Y(n_237)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_179),
.B(n_2),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_15),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_209),
.A2(n_11),
.B(n_4),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_225),
.B(n_6),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_228),
.B(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_233),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_231),
.B(n_12),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_210),
.B(n_206),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_221),
.C(n_219),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_10),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_235),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_11),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_229),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_234),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_235),
.A2(n_220),
.B(n_226),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_244),
.B(n_14),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_14),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_238),
.Y(n_246)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_246),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_249),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_2),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_SL g251 ( 
.A(n_250),
.B(n_15),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_251),
.Y(n_254)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_252),
.Y(n_255)
);

AOI321xp33_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_239),
.A3(n_247),
.B1(n_249),
.B2(n_253),
.C(n_254),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_253),
.Y(n_257)
);


endmodule