module real_jpeg_2272_n_16 (n_5, n_4, n_8, n_0, n_12, n_325, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_325;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_1),
.A2(n_29),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_1),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_1),
.A2(n_39),
.B1(n_63),
.B2(n_65),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_1),
.A2(n_39),
.B1(n_58),
.B2(n_59),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_2),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_2),
.A2(n_35),
.B1(n_63),
.B2(n_65),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_2),
.A2(n_35),
.B1(n_58),
.B2(n_59),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_67),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_3),
.A2(n_29),
.B1(n_36),
.B2(n_67),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_3),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_5),
.A2(n_63),
.B1(n_65),
.B2(n_69),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_5),
.A2(n_29),
.B1(n_36),
.B2(n_69),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_69),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_109),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_6),
.A2(n_29),
.B1(n_36),
.B2(n_109),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_6),
.A2(n_63),
.B1(n_65),
.B2(n_109),
.Y(n_191)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_11),
.A2(n_63),
.B1(n_65),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_11),
.A2(n_29),
.B1(n_36),
.B2(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_72),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_72),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_12),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_12),
.B(n_29),
.C(n_43),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_12),
.B(n_32),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_12),
.B(n_119),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_12),
.B(n_65),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_65),
.B(n_182),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_12),
.B(n_126),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_12),
.A2(n_58),
.B(n_220),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_14),
.A2(n_29),
.B1(n_36),
.B2(n_48),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_14),
.A2(n_48),
.B1(n_63),
.B2(n_65),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_14),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_316),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_306),
.B(n_315),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_272),
.B(n_303),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_249),
.B(n_271),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_135),
.B(n_248),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_110),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_22),
.B(n_110),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_82),
.C(n_93),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_23),
.B(n_82),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_53),
.B2(n_54),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_24),
.B(n_55),
.C(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_26),
.B(n_40),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_37),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_27),
.A2(n_31),
.B(n_86),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_27),
.A2(n_31),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_27),
.A2(n_37),
.B(n_86),
.Y(n_184)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_28),
.B(n_38),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_28),
.A2(n_32),
.B1(n_34),
.B2(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_28),
.A2(n_85),
.B(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_28),
.A2(n_32),
.B1(n_98),
.B2(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_28),
.A2(n_32),
.B1(n_162),
.B2(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_29),
.B(n_160),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_31),
.B(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_31),
.A2(n_88),
.B(n_102),
.Y(n_210)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_38),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B(n_49),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_41),
.A2(n_44),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_41),
.A2(n_91),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_41),
.B(n_199),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_52)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OA22x2_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_46),
.B1(n_75),
.B2(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_45),
.B(n_77),
.Y(n_183)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_46),
.B(n_152),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_46),
.A2(n_65),
.A3(n_75),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_49),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_50),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_51),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_51),
.A2(n_119),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_51),
.A2(n_119),
.B1(n_147),
.B2(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_51),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_51),
.A2(n_119),
.B(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_70),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_62),
.B1(n_66),
.B2(n_68),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_56),
.A2(n_62),
.B1(n_66),
.B2(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_56),
.A2(n_68),
.B(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_56),
.A2(n_62),
.B1(n_108),
.B2(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_56),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_56),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_56),
.A2(n_62),
.B1(n_277),
.B2(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_56),
.A2(n_260),
.B(n_287),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_98),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_61),
.C(n_65),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_60),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_63),
.B(n_97),
.C(n_99),
.Y(n_96)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_62),
.A2(n_277),
.B(n_278),
.Y(n_276)
);

CKINVDCx6p67_ASAP7_75t_R g65 ( 
.A(n_63),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_65),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B(n_79),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_71),
.A2(n_73),
.B(n_78),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_73),
.A2(n_78),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_73),
.A2(n_78),
.B1(n_104),
.B2(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_78),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_78),
.B(n_98),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_79),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_81),
.A2(n_131),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_81),
.A2(n_131),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_90),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_92),
.B(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_91),
.A2(n_118),
.B(n_199),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_93),
.B(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.C(n_107),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_94),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_95),
.A2(n_96),
.B1(n_100),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_97),
.Y(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_100),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_103),
.B(n_107),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_105),
.B(n_130),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_134),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_114),
.B(n_121),
.C(n_134),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_115),
.A2(n_116),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_116),
.B(n_117),
.Y(n_262)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_116),
.A2(n_257),
.B(n_262),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_132),
.B2(n_133),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_124),
.B(n_128),
.C(n_133),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_125),
.B(n_278),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_126),
.B(n_261),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_127),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_129),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_131),
.A2(n_268),
.B(n_281),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_132),
.Y(n_133)
);

AOI321xp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_230),
.A3(n_240),
.B1(n_246),
.B2(n_247),
.C(n_325),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_213),
.B(n_229),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_193),
.B(n_212),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_175),
.B(n_192),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_156),
.B(n_174),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_149),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_149),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_146),
.C(n_177),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_143),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_168),
.B(n_173),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_163),
.B(n_167),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_166),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_172),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_178),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_186),
.C(n_189),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_211),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_211),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_200),
.C(n_201),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_198),
.B(n_265),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_199),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_208),
.C(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_215),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_224),
.B2(n_225),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_226),
.C(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_222),
.C(n_223),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_233),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_239),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_235),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_270),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_270),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_255),
.C(n_263),
.Y(n_301)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_263),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_261),
.B(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_266),
.B(n_269),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_266),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_295),
.C(n_299),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_269),
.B(n_295),
.CI(n_299),
.CON(n_302),
.SN(n_302)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_300),
.Y(n_272)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_273),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_294),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_294),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_284),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_276),
.C(n_293),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_280),
.C(n_282),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_285),
.B1(n_292),
.B2(n_293),
.Y(n_284)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_276),
.A2(n_292),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_282),
.B1(n_291),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_282),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_286),
.C(n_290),
.Y(n_314)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_302),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_302),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_308),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_314),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_312),
.C(n_314),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_321),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_320),
.Y(n_322)
);


endmodule