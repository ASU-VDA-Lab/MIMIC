module fake_ibex_489_n_957 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_957);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_957;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_375;
wire n_280;
wire n_317;
wire n_340;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_497;
wire n_243;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_562;
wire n_506;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_520;
wire n_411;
wire n_927;
wire n_684;
wire n_775;
wire n_934;
wire n_784;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_288;
wire n_379;
wire n_247;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_164;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_8),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_5),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_34),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_1),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_70),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_53),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_33),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_35),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_3),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_46),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_65),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_34),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_56),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_76),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_31),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_125),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_2),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_35),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_71),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_87),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_121),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_119),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_59),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_95),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_143),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_88),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_50),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_81),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_84),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_141),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_7),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_54),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_49),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_7),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_14),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_66),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_100),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_10),
.B(n_110),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_28),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_130),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_41),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_27),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_61),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_30),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_13),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_148),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_99),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_5),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_101),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_107),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_147),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_85),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_21),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_78),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_45),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_123),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_97),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_106),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_55),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_62),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_115),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_137),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_11),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_118),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_159),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_68),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_144),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_112),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_21),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_94),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_51),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_91),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_127),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_8),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_38),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_77),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_129),
.B(n_4),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_153),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_116),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_15),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_48),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_82),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_73),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_24),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_L g262 ( 
.A(n_86),
.B(n_1),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_29),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_80),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_105),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_52),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_142),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_64),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_3),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_30),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_19),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_89),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_138),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_63),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_39),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_149),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_13),
.B(n_44),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_160),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_31),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_104),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_74),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_58),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_14),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_98),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_27),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_120),
.Y(n_286)
);

AND2x6_ASAP7_75t_L g287 ( 
.A(n_176),
.B(n_40),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_233),
.B(n_0),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_213),
.B(n_0),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_213),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_163),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_168),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_168),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_239),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_176),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_227),
.B(n_2),
.Y(n_297)
);

OAI22x1_ASAP7_75t_L g298 ( 
.A1(n_163),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_298)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_195),
.B(n_42),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_185),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_169),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_231),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_170),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_179),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_195),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_188),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_193),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_175),
.Y(n_310)
);

AOI22x1_ASAP7_75t_SL g311 ( 
.A1(n_172),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_311)
);

AOI22x1_ASAP7_75t_SL g312 ( 
.A1(n_173),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_261),
.B(n_12),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_175),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_184),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_185),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_194),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_248),
.B(n_16),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_17),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_185),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_241),
.B(n_232),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_241),
.B(n_17),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g323 ( 
.A1(n_184),
.A2(n_92),
.B(n_157),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_196),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_189),
.Y(n_325)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_182),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_164),
.Y(n_327)
);

AND2x4_ASAP7_75t_L g328 ( 
.A(n_189),
.B(n_18),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_191),
.B(n_18),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_191),
.B(n_19),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_166),
.Y(n_331)
);

BUFx8_ASAP7_75t_L g332 ( 
.A(n_277),
.Y(n_332)
);

OA21x2_ASAP7_75t_L g333 ( 
.A1(n_197),
.A2(n_93),
.B(n_152),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_197),
.Y(n_334)
);

AO22x1_ASAP7_75t_L g335 ( 
.A1(n_171),
.A2(n_283),
.B1(n_277),
.B2(n_246),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_177),
.B(n_20),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_200),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_201),
.B(n_20),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_167),
.Y(n_339)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_226),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_203),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_206),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_165),
.B(n_174),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_187),
.B(n_22),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_177),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_226),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_234),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_204),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_204),
.B(n_23),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_234),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_249),
.B(n_25),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_249),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_207),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_205),
.B(n_25),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_210),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_205),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_212),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_214),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_217),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_180),
.B(n_26),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_218),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_219),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_183),
.B(n_26),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_220),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_221),
.B(n_28),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_223),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_230),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_242),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_222),
.B(n_228),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_285),
.B(n_29),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_244),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_222),
.B(n_32),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_199),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_245),
.Y(n_374)
);

BUFx8_ASAP7_75t_L g375 ( 
.A(n_250),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_253),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_329),
.B(n_266),
.Y(n_377)
);

BUFx4f_ASAP7_75t_L g378 ( 
.A(n_300),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_302),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_306),
.B(n_224),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_289),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_289),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_289),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_287),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_289),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_323),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_334),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_305),
.B(n_257),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_329),
.B(n_272),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_306),
.B(n_257),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_329),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_326),
.A2(n_263),
.B1(n_269),
.B2(n_275),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_316),
.B(n_263),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_330),
.Y(n_394)
);

INVxp33_ASAP7_75t_SL g395 ( 
.A(n_343),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_332),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_330),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_334),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_330),
.B(n_273),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_330),
.B(n_274),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g402 ( 
.A(n_351),
.B(n_276),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_351),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_351),
.A2(n_252),
.B1(n_209),
.B2(n_279),
.Y(n_404)
);

BUFx4f_ASAP7_75t_L g405 ( 
.A(n_300),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_328),
.B(n_281),
.Y(n_407)
);

OR2x6_ASAP7_75t_L g408 ( 
.A(n_335),
.B(n_215),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_334),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_369),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_323),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_307),
.Y(n_412)
);

NOR3xp33_ASAP7_75t_L g413 ( 
.A(n_348),
.B(n_269),
.C(n_216),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_307),
.Y(n_414)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_316),
.Y(n_415)
);

INVxp67_ASAP7_75t_R g416 ( 
.A(n_344),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_307),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_287),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_316),
.B(n_300),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_320),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_L g421 ( 
.A1(n_305),
.A2(n_270),
.B1(n_271),
.B2(n_251),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_320),
.B(n_165),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_328),
.A2(n_284),
.B1(n_208),
.B2(n_202),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_328),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

OR2x6_ASAP7_75t_L g427 ( 
.A(n_335),
.B(n_254),
.Y(n_427)
);

NAND2x1_ASAP7_75t_L g428 ( 
.A(n_344),
.B(n_262),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_301),
.B(n_174),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_321),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_320),
.B(n_178),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_307),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_301),
.B(n_186),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_375),
.B(n_181),
.Y(n_436)
);

BUFx4f_ASAP7_75t_L g437 ( 
.A(n_326),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_321),
.B(n_186),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_302),
.B(n_192),
.Y(n_440)
);

BUFx8_ASAP7_75t_SL g441 ( 
.A(n_313),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_321),
.B(n_190),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_355),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_333),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_355),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_292),
.B(n_190),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_355),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_303),
.A2(n_240),
.B1(n_282),
.B2(n_280),
.Y(n_448)
);

AND3x2_ASAP7_75t_L g449 ( 
.A(n_313),
.B(n_238),
.C(n_258),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_333),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_L g451 ( 
.A(n_287),
.B(n_211),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_303),
.B(n_286),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_355),
.Y(n_454)
);

INVxp33_ASAP7_75t_SL g455 ( 
.A(n_345),
.Y(n_455)
);

BUFx4f_ASAP7_75t_L g456 ( 
.A(n_326),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_304),
.B(n_308),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_327),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_358),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_327),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_333),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_287),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_339),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_304),
.B(n_225),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_308),
.B(n_225),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_339),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_296),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_309),
.B(n_286),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_356),
.B(n_229),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_358),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_287),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_332),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_358),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_309),
.B(n_282),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_331),
.B(n_280),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_332),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_317),
.B(n_278),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_317),
.B(n_278),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_287),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_373),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_373),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_375),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_346),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_297),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_299),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_324),
.B(n_268),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_368),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_346),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_368),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_368),
.Y(n_490)
);

OAI21xp33_ASAP7_75t_SL g491 ( 
.A1(n_337),
.A2(n_32),
.B(n_33),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_299),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_350),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_350),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_322),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_299),
.Y(n_496)
);

OAI22xp33_ASAP7_75t_L g497 ( 
.A1(n_288),
.A2(n_336),
.B1(n_354),
.B2(n_372),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_368),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_375),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_340),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_410),
.B(n_297),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_441),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_384),
.B(n_319),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_384),
.B(n_319),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_467),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_388),
.B(n_349),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_495),
.B(n_337),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_464),
.B(n_349),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_464),
.B(n_341),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_474),
.B(n_341),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_474),
.B(n_342),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_467),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_430),
.Y(n_513)
);

AND2x6_ASAP7_75t_SL g514 ( 
.A(n_408),
.B(n_370),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_475),
.B(n_359),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_402),
.A2(n_359),
.B1(n_374),
.B2(n_371),
.Y(n_516)
);

A2O1A1Ixp33_ASAP7_75t_L g517 ( 
.A1(n_425),
.A2(n_362),
.B(n_367),
.C(n_366),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_384),
.B(n_318),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_437),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_442),
.B(n_361),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_392),
.B(n_370),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_408),
.B(n_298),
.Y(n_522)
);

BUFx12f_ASAP7_75t_L g523 ( 
.A(n_379),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_442),
.B(n_361),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_460),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_438),
.B(n_362),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_472),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_476),
.B(n_366),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_438),
.B(n_367),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_481),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_393),
.B(n_353),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_497),
.A2(n_338),
.B1(n_365),
.B2(n_259),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_481),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_402),
.A2(n_376),
.B1(n_364),
.B2(n_357),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_491),
.A2(n_312),
.B1(n_311),
.B2(n_290),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_458),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_408),
.A2(n_376),
.B1(n_364),
.B2(n_357),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_382),
.Y(n_538)
);

O2A1O1Ixp33_ASAP7_75t_L g539 ( 
.A1(n_381),
.A2(n_295),
.B(n_290),
.C(n_291),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_463),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_466),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_438),
.B(n_296),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_396),
.B(n_290),
.Y(n_543)
);

CKINVDCx11_ASAP7_75t_R g544 ( 
.A(n_427),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_480),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_419),
.B(n_235),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_402),
.A2(n_299),
.B1(n_347),
.B2(n_293),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_484),
.B(n_291),
.Y(n_549)
);

OAI221xp5_ASAP7_75t_L g550 ( 
.A1(n_404),
.A2(n_295),
.B1(n_291),
.B2(n_294),
.C(n_352),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_455),
.A2(n_440),
.B1(n_427),
.B2(n_395),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_415),
.B(n_264),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_390),
.B(n_380),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_427),
.A2(n_298),
.B1(n_311),
.B2(n_312),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_415),
.B(n_260),
.Y(n_555)
);

AO22x1_ASAP7_75t_L g556 ( 
.A1(n_395),
.A2(n_299),
.B1(n_236),
.B2(n_243),
.Y(n_556)
);

A2O1A1Ixp33_ASAP7_75t_L g557 ( 
.A1(n_426),
.A2(n_294),
.B(n_325),
.C(n_315),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_413),
.A2(n_299),
.B1(n_236),
.B2(n_243),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_446),
.A2(n_299),
.B1(n_247),
.B2(n_256),
.Y(n_559)
);

O2A1O1Ixp33_ASAP7_75t_L g560 ( 
.A1(n_383),
.A2(n_314),
.B(n_310),
.C(n_315),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_500),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_420),
.B(n_325),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_451),
.A2(n_333),
.B(n_314),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_469),
.A2(n_256),
.B1(n_255),
.B2(n_247),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_493),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_422),
.B(n_198),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_431),
.B(n_340),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_429),
.B(n_340),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_494),
.B(n_340),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_434),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_416),
.B(n_340),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_428),
.B(n_113),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_434),
.B(n_36),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_452),
.B(n_36),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_378),
.B(n_114),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_418),
.B(n_111),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_452),
.B(n_37),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_465),
.B(n_37),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_433),
.A2(n_38),
.B1(n_43),
.B2(n_47),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_441),
.Y(n_580)
);

BUFx8_ASAP7_75t_L g581 ( 
.A(n_436),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_418),
.B(n_57),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_439),
.A2(n_60),
.B1(n_67),
.B2(n_69),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_468),
.B(n_72),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_451),
.A2(n_75),
.B(n_79),
.Y(n_585)
);

A2O1A1Ixp33_ASAP7_75t_L g586 ( 
.A1(n_435),
.A2(n_90),
.B(n_102),
.C(n_103),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_456),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_468),
.B(n_124),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_404),
.A2(n_126),
.B1(n_128),
.B2(n_132),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_L g590 ( 
.A1(n_424),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_462),
.B(n_136),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_477),
.B(n_478),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_423),
.A2(n_140),
.B1(n_145),
.B2(n_146),
.Y(n_593)
);

BUFx8_ASAP7_75t_L g594 ( 
.A(n_523),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_563),
.A2(n_444),
.B(n_450),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_538),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_563),
.A2(n_444),
.B(n_450),
.Y(n_597)
);

OA21x2_ASAP7_75t_L g598 ( 
.A1(n_585),
.A2(n_394),
.B(n_406),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_501),
.B(n_448),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_538),
.Y(n_600)
);

O2A1O1Ixp33_ASAP7_75t_L g601 ( 
.A1(n_517),
.A2(n_407),
.B(n_391),
.C(n_403),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_513),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_513),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_507),
.B(n_448),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_528),
.B(n_499),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_565),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_508),
.B(n_486),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_562),
.Y(n_608)
);

O2A1O1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_550),
.A2(n_407),
.B(n_397),
.C(n_377),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_506),
.B(n_477),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_553),
.B(n_515),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_545),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_509),
.A2(n_461),
.B(n_444),
.Y(n_613)
);

O2A1O1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_550),
.A2(n_389),
.B(n_400),
.C(n_399),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_545),
.B(n_482),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_526),
.B(n_439),
.Y(n_616)
);

NOR3xp33_ASAP7_75t_L g617 ( 
.A(n_554),
.B(n_421),
.C(n_457),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_529),
.B(n_385),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_570),
.B(n_457),
.Y(n_619)
);

O2A1O1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_520),
.A2(n_389),
.B(n_399),
.C(n_488),
.Y(n_620)
);

NAND2x1p5_ASAP7_75t_L g621 ( 
.A(n_528),
.B(n_462),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_510),
.A2(n_450),
.B(n_461),
.Y(n_622)
);

NOR2xp67_ASAP7_75t_L g623 ( 
.A(n_502),
.B(n_483),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_527),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_570),
.B(n_405),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_516),
.A2(n_479),
.B1(n_496),
.B2(n_471),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_511),
.B(n_405),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_564),
.B(n_449),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_524),
.A2(n_450),
.B(n_461),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_535),
.A2(n_411),
.B1(n_386),
.B2(n_444),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_505),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_581),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_592),
.A2(n_461),
.B(n_492),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_562),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_543),
.Y(n_635)
);

A2O1A1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_531),
.A2(n_386),
.B(n_411),
.C(n_490),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_522),
.A2(n_485),
.B1(n_479),
.B2(n_386),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_534),
.B(n_411),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_549),
.Y(n_639)
);

BUFx12f_ASAP7_75t_L g640 ( 
.A(n_544),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_536),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_512),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_537),
.B(n_489),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_540),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_519),
.B(n_587),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_581),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_518),
.A2(n_498),
.B(n_487),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_569),
.Y(n_648)
);

BUFx12f_ASAP7_75t_L g649 ( 
.A(n_514),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_569),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_548),
.B(n_473),
.C(n_470),
.Y(n_651)
);

NOR2x1_ASAP7_75t_L g652 ( 
.A(n_522),
.B(n_573),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_559),
.B(n_470),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_503),
.A2(n_459),
.B(n_454),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_558),
.B(n_454),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_541),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_504),
.A2(n_453),
.B(n_447),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_521),
.Y(n_658)
);

CKINVDCx14_ASAP7_75t_R g659 ( 
.A(n_522),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_532),
.B(n_453),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_542),
.B(n_447),
.Y(n_661)
);

AO22x1_ASAP7_75t_L g662 ( 
.A1(n_580),
.A2(n_445),
.B1(n_443),
.B2(n_412),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_551),
.B(n_432),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_557),
.A2(n_567),
.B(n_568),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_560),
.A2(n_539),
.B(n_590),
.C(n_578),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_547),
.A2(n_417),
.B1(n_414),
.B2(n_412),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_556),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_535),
.A2(n_387),
.B1(n_398),
.B2(n_401),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_539),
.B(n_398),
.Y(n_669)
);

INVxp33_ASAP7_75t_SL g670 ( 
.A(n_566),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_561),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_571),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_546),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_624),
.B(n_574),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_612),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_648),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_629),
.A2(n_560),
.B(n_577),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_621),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_658),
.B(n_533),
.Y(n_679)
);

NOR2x1_ASAP7_75t_L g680 ( 
.A(n_652),
.B(n_590),
.Y(n_680)
);

AOI221x1_ASAP7_75t_L g681 ( 
.A1(n_630),
.A2(n_586),
.B1(n_589),
.B2(n_584),
.C(n_588),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_606),
.Y(n_682)
);

O2A1O1Ixp33_ASAP7_75t_SL g683 ( 
.A1(n_636),
.A2(n_591),
.B(n_582),
.C(n_576),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_L g684 ( 
.A(n_621),
.B(n_611),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_599),
.B(n_525),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_615),
.B(n_552),
.Y(n_686)
);

AO31x2_ASAP7_75t_L g687 ( 
.A1(n_595),
.A2(n_575),
.A3(n_572),
.B(n_409),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_604),
.B(n_530),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_670),
.B(n_610),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_668),
.A2(n_593),
.B1(n_579),
.B2(n_583),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_594),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_617),
.B(n_555),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_622),
.A2(n_158),
.B(n_629),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_594),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_639),
.B(n_635),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_660),
.A2(n_628),
.B1(n_607),
.B2(n_627),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_641),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_SL g698 ( 
.A1(n_626),
.A2(n_598),
.B(n_665),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_648),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_672),
.B(n_608),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_640),
.Y(n_701)
);

AO31x2_ASAP7_75t_L g702 ( 
.A1(n_664),
.A2(n_633),
.A3(n_669),
.B(n_666),
.Y(n_702)
);

O2A1O1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_665),
.A2(n_620),
.B(n_601),
.C(n_609),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_623),
.B(n_634),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_644),
.B(n_656),
.Y(n_705)
);

NAND2x1p5_ASAP7_75t_L g706 ( 
.A(n_632),
.B(n_650),
.Y(n_706)
);

O2A1O1Ixp5_ASAP7_75t_L g707 ( 
.A1(n_662),
.A2(n_655),
.B(n_653),
.C(n_667),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_673),
.B(n_645),
.Y(n_708)
);

O2A1O1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_620),
.A2(n_601),
.B(n_609),
.C(n_614),
.Y(n_709)
);

OAI221xp5_ASAP7_75t_L g710 ( 
.A1(n_618),
.A2(n_616),
.B1(n_625),
.B2(n_663),
.C(n_614),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_619),
.B(n_645),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_646),
.Y(n_712)
);

CKINVDCx12_ASAP7_75t_R g713 ( 
.A(n_663),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_637),
.A2(n_598),
.B1(n_659),
.B2(n_643),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_596),
.B(n_600),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_647),
.A2(n_657),
.B(n_654),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_L g717 ( 
.A1(n_654),
.A2(n_657),
.B(n_651),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_631),
.A2(n_642),
.B1(n_661),
.B2(n_603),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_631),
.A2(n_642),
.B1(n_602),
.B2(n_671),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_649),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_606),
.Y(n_721)
);

AO31x2_ASAP7_75t_L g722 ( 
.A1(n_636),
.A2(n_595),
.A3(n_597),
.B(n_613),
.Y(n_722)
);

NAND3xp33_ASAP7_75t_SL g723 ( 
.A(n_605),
.B(n_379),
.C(n_436),
.Y(n_723)
);

AO31x2_ASAP7_75t_L g724 ( 
.A1(n_636),
.A2(n_595),
.A3(n_597),
.B(n_613),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_624),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_595),
.A2(n_597),
.B(n_638),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_648),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_624),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_606),
.Y(n_729)
);

OAI22x1_ASAP7_75t_L g730 ( 
.A1(n_624),
.A2(n_545),
.B1(n_370),
.B2(n_440),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_611),
.B(n_599),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_611),
.B(n_599),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_611),
.B(n_599),
.Y(n_733)
);

OAI21xp33_ASAP7_75t_L g734 ( 
.A1(n_611),
.A2(n_604),
.B(n_599),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_611),
.B(n_599),
.Y(n_735)
);

NAND3xp33_ASAP7_75t_L g736 ( 
.A(n_636),
.B(n_665),
.C(n_668),
.Y(n_736)
);

CKINVDCx11_ASAP7_75t_R g737 ( 
.A(n_640),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_611),
.B(n_599),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_606),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_606),
.Y(n_740)
);

AND2x2_ASAP7_75t_SL g741 ( 
.A(n_624),
.B(n_436),
.Y(n_741)
);

INVx5_ASAP7_75t_L g742 ( 
.A(n_648),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_606),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_595),
.A2(n_597),
.B(n_613),
.Y(n_744)
);

AO31x2_ASAP7_75t_L g745 ( 
.A1(n_636),
.A2(n_595),
.A3(n_597),
.B(n_613),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_611),
.B(n_599),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_658),
.B(n_545),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_612),
.B(n_545),
.Y(n_748)
);

AO31x2_ASAP7_75t_L g749 ( 
.A1(n_636),
.A2(n_595),
.A3(n_597),
.B(n_613),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_595),
.A2(n_597),
.B(n_613),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_606),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_594),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_595),
.A2(n_597),
.B(n_638),
.Y(n_753)
);

CKINVDCx6p67_ASAP7_75t_R g754 ( 
.A(n_640),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_595),
.A2(n_597),
.B(n_613),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_611),
.A2(n_553),
.B(n_665),
.C(n_620),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_611),
.B(n_599),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_611),
.B(n_599),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_606),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_611),
.A2(n_553),
.B(n_665),
.C(n_620),
.Y(n_760)
);

AOI221xp5_ASAP7_75t_SL g761 ( 
.A1(n_665),
.A2(n_630),
.B1(n_609),
.B2(n_604),
.C(n_550),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_682),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_737),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_731),
.B(n_732),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_678),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_752),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_689),
.B(n_725),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_759),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_697),
.Y(n_769)
);

NOR2xp67_ASAP7_75t_L g770 ( 
.A(n_694),
.B(n_730),
.Y(n_770)
);

AO21x2_ASAP7_75t_L g771 ( 
.A1(n_698),
.A2(n_753),
.B(n_726),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_676),
.Y(n_772)
);

OAI21x1_ASAP7_75t_SL g773 ( 
.A1(n_680),
.A2(n_719),
.B(n_758),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_721),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_728),
.B(n_748),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_676),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_756),
.A2(n_760),
.B(n_693),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_691),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_717),
.A2(n_734),
.B(n_683),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_744),
.A2(n_755),
.B(n_750),
.Y(n_780)
);

AOI21xp33_ASAP7_75t_SL g781 ( 
.A1(n_741),
.A2(n_720),
.B(n_712),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_733),
.B(n_735),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_717),
.A2(n_734),
.B(n_684),
.Y(n_783)
);

OR2x6_ASAP7_75t_L g784 ( 
.A(n_701),
.B(n_706),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_729),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_675),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_699),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_708),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_739),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_747),
.B(n_708),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_740),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_743),
.Y(n_792)
);

AO21x2_ASAP7_75t_L g793 ( 
.A1(n_736),
.A2(n_714),
.B(n_677),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_738),
.B(n_746),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_757),
.B(n_696),
.Y(n_795)
);

CKINVDCx6p67_ASAP7_75t_R g796 ( 
.A(n_754),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_696),
.B(n_692),
.Y(n_797)
);

OA21x2_ASAP7_75t_L g798 ( 
.A1(n_761),
.A2(n_681),
.B(n_716),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_710),
.A2(n_703),
.B(n_709),
.C(n_690),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_751),
.B(n_705),
.Y(n_800)
);

OA21x2_ASAP7_75t_L g801 ( 
.A1(n_761),
.A2(n_677),
.B(n_707),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_680),
.B(n_690),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_711),
.B(n_686),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_676),
.Y(n_804)
);

AO31x2_ASAP7_75t_L g805 ( 
.A1(n_719),
.A2(n_685),
.A3(n_688),
.B(n_715),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_713),
.Y(n_806)
);

AOI21xp33_ASAP7_75t_L g807 ( 
.A1(n_679),
.A2(n_674),
.B(n_700),
.Y(n_807)
);

AO31x2_ASAP7_75t_L g808 ( 
.A1(n_702),
.A2(n_687),
.A3(n_749),
.B(n_745),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_742),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_695),
.Y(n_810)
);

INVx6_ASAP7_75t_L g811 ( 
.A(n_742),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_718),
.A2(n_742),
.B1(n_704),
.B2(n_699),
.Y(n_812)
);

AO21x2_ASAP7_75t_L g813 ( 
.A1(n_722),
.A2(n_749),
.B(n_745),
.Y(n_813)
);

OAI21x1_ASAP7_75t_L g814 ( 
.A1(n_722),
.A2(n_724),
.B(n_727),
.Y(n_814)
);

AO31x2_ASAP7_75t_L g815 ( 
.A1(n_702),
.A2(n_687),
.A3(n_722),
.B(n_724),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_727),
.B(n_723),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_699),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_756),
.A2(n_760),
.B(n_611),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_748),
.B(n_545),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_731),
.B(n_732),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_731),
.B(n_732),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_748),
.B(n_545),
.Y(n_822)
);

BUFx8_ASAP7_75t_L g823 ( 
.A(n_691),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_748),
.B(n_545),
.Y(n_824)
);

OAI21xp33_ASAP7_75t_L g825 ( 
.A1(n_747),
.A2(n_455),
.B(n_545),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_725),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_809),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_L g828 ( 
.A(n_818),
.B(n_825),
.C(n_795),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_773),
.B(n_799),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_797),
.B(n_799),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_802),
.B(n_805),
.Y(n_831)
);

INVxp33_ASAP7_75t_L g832 ( 
.A(n_819),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_777),
.A2(n_783),
.B(n_802),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_765),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_805),
.B(n_813),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_814),
.B(n_771),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_769),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_785),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_791),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_808),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_808),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_777),
.A2(n_783),
.B(n_779),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_779),
.A2(n_821),
.B(n_820),
.Y(n_843)
);

NOR2xp67_ASAP7_75t_L g844 ( 
.A(n_816),
.B(n_817),
.Y(n_844)
);

OR2x6_ASAP7_75t_L g845 ( 
.A(n_812),
.B(n_780),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_770),
.A2(n_807),
.B1(n_790),
.B2(n_803),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_764),
.B(n_782),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_794),
.B(n_800),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_808),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_817),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_815),
.B(n_798),
.Y(n_851)
);

CKINVDCx6p67_ASAP7_75t_R g852 ( 
.A(n_796),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_809),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_815),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_787),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_850),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_840),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_830),
.B(n_793),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_847),
.B(n_778),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_840),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_841),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_835),
.B(n_801),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_855),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_843),
.B(n_789),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_836),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_850),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_849),
.B(n_775),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_843),
.B(n_792),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_835),
.B(n_774),
.Y(n_869)
);

NAND2x1_ASAP7_75t_L g870 ( 
.A(n_845),
.B(n_811),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_851),
.B(n_762),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_827),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_851),
.B(n_768),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_867),
.B(n_854),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_863),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_857),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_856),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_869),
.B(n_831),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_867),
.B(n_869),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_869),
.B(n_831),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_871),
.B(n_847),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_857),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_860),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_860),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_865),
.B(n_836),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_861),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_861),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_871),
.B(n_831),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_876),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_888),
.B(n_862),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_879),
.B(n_856),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_888),
.B(n_862),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_876),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_881),
.B(n_871),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_882),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_875),
.B(n_844),
.Y(n_896)
);

NAND4xp25_ASAP7_75t_L g897 ( 
.A(n_874),
.B(n_846),
.C(n_859),
.D(n_828),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_879),
.B(n_873),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_878),
.B(n_873),
.Y(n_899)
);

NAND2xp33_ASAP7_75t_SL g900 ( 
.A(n_875),
.B(n_870),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_882),
.Y(n_901)
);

NOR2x1_ASAP7_75t_L g902 ( 
.A(n_874),
.B(n_872),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_890),
.B(n_878),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_889),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_891),
.B(n_890),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_892),
.B(n_880),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_893),
.Y(n_907)
);

OR2x2_ASAP7_75t_L g908 ( 
.A(n_899),
.B(n_880),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_895),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_901),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_892),
.B(n_877),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_898),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_897),
.B(n_846),
.C(n_858),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_894),
.B(n_862),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_905),
.Y(n_915)
);

OAI221xp5_ASAP7_75t_L g916 ( 
.A1(n_913),
.A2(n_900),
.B1(n_902),
.B2(n_896),
.C(n_781),
.Y(n_916)
);

AOI221xp5_ASAP7_75t_L g917 ( 
.A1(n_912),
.A2(n_786),
.B1(n_826),
.B2(n_900),
.C(n_828),
.Y(n_917)
);

NOR2x2_ASAP7_75t_L g918 ( 
.A(n_904),
.B(n_829),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_905),
.A2(n_896),
.B1(n_872),
.B2(n_852),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_914),
.B(n_866),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_911),
.A2(n_844),
.B(n_848),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_904),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_907),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_908),
.B(n_903),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_907),
.Y(n_925)
);

AOI322xp5_ASAP7_75t_L g926 ( 
.A1(n_903),
.A2(n_806),
.A3(n_872),
.B1(n_827),
.B2(n_853),
.C1(n_838),
.C2(n_839),
.Y(n_926)
);

AOI322xp5_ASAP7_75t_L g927 ( 
.A1(n_924),
.A2(n_906),
.A3(n_914),
.B1(n_909),
.B2(n_806),
.C1(n_910),
.C2(n_827),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_920),
.Y(n_928)
);

O2A1O1Ixp5_ASAP7_75t_L g929 ( 
.A1(n_919),
.A2(n_924),
.B(n_921),
.C(n_915),
.Y(n_929)
);

AOI221x1_ASAP7_75t_L g930 ( 
.A1(n_922),
.A2(n_837),
.B1(n_838),
.B2(n_839),
.C(n_910),
.Y(n_930)
);

AOI221xp5_ASAP7_75t_L g931 ( 
.A1(n_916),
.A2(n_906),
.B1(n_832),
.B2(n_886),
.C(n_884),
.Y(n_931)
);

AOI222xp33_ASAP7_75t_L g932 ( 
.A1(n_917),
.A2(n_853),
.B1(n_832),
.B2(n_823),
.C1(n_837),
.C2(n_848),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_923),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_930),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_931),
.A2(n_918),
.B1(n_852),
.B2(n_925),
.Y(n_935)
);

NOR2x1_ASAP7_75t_L g936 ( 
.A(n_929),
.B(n_766),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_928),
.B(n_926),
.Y(n_937)
);

NOR4xp75_ASAP7_75t_L g938 ( 
.A(n_929),
.B(n_852),
.C(n_870),
.D(n_823),
.Y(n_938)
);

NAND4xp75_ASAP7_75t_L g939 ( 
.A(n_933),
.B(n_918),
.C(n_868),
.D(n_864),
.Y(n_939)
);

NAND5xp2_ASAP7_75t_L g940 ( 
.A(n_937),
.B(n_932),
.C(n_927),
.D(n_763),
.E(n_833),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_936),
.A2(n_853),
.B1(n_829),
.B2(n_885),
.Y(n_941)
);

NAND5xp2_ASAP7_75t_L g942 ( 
.A(n_934),
.B(n_833),
.C(n_842),
.D(n_822),
.E(n_824),
.Y(n_942)
);

AOI221xp5_ASAP7_75t_L g943 ( 
.A1(n_935),
.A2(n_887),
.B1(n_886),
.B2(n_883),
.C(n_884),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_941),
.A2(n_943),
.B(n_939),
.Y(n_944)
);

NOR3xp33_ASAP7_75t_L g945 ( 
.A(n_940),
.B(n_938),
.C(n_804),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_L g946 ( 
.A(n_942),
.B(n_776),
.C(n_772),
.Y(n_946)
);

NAND4xp25_ASAP7_75t_L g947 ( 
.A(n_940),
.B(n_834),
.C(n_767),
.D(n_766),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_944),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_SL g949 ( 
.A(n_947),
.B(n_945),
.C(n_946),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_948),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_949),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_SL g952 ( 
.A1(n_951),
.A2(n_784),
.B1(n_811),
.B2(n_834),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_952),
.A2(n_951),
.B1(n_950),
.B2(n_784),
.Y(n_953)
);

AOI21xp33_ASAP7_75t_L g954 ( 
.A1(n_953),
.A2(n_784),
.B(n_776),
.Y(n_954)
);

XNOR2xp5_ASAP7_75t_L g955 ( 
.A(n_954),
.B(n_788),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_955),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_SL g957 ( 
.A1(n_956),
.A2(n_810),
.B1(n_772),
.B2(n_765),
.Y(n_957)
);


endmodule