module fake_jpeg_1358_n_385 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_385);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_385;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_2),
.B(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_16),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_45),
.B(n_61),
.Y(n_125)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_66),
.Y(n_89)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_29),
.B(n_12),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_11),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_62),
.Y(n_99)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_34),
.Y(n_62)
);

CKINVDCx9p33_ASAP7_75t_R g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_26),
.B(n_11),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_82),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_39),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_32),
.B(n_11),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_17),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_83),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_40),
.B1(n_39),
.B2(n_41),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_84),
.A2(n_92),
.B1(n_96),
.B2(n_107),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_90),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_27),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_91),
.B(n_103),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_47),
.A2(n_39),
.B1(n_34),
.B2(n_41),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_63),
.A2(n_39),
.B1(n_38),
.B2(n_22),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_93),
.A2(n_104),
.B1(n_120),
.B2(n_55),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_36),
.B1(n_32),
.B2(n_28),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_94),
.A2(n_65),
.B1(n_44),
.B2(n_3),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_48),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_52),
.B(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_27),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_61),
.A2(n_38),
.B1(n_20),
.B2(n_18),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_58),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_57),
.A2(n_28),
.B1(n_42),
.B2(n_35),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_109),
.A2(n_118),
.B1(n_44),
.B2(n_5),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_30),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_132),
.B(n_78),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_17),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_103),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_30),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_33),
.B1(n_42),
.B2(n_35),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_51),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_33),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_56),
.B(n_10),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_78),
.A2(n_23),
.B(n_17),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_59),
.B(n_10),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_0),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_134),
.B(n_137),
.Y(n_184)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_85),
.B(n_73),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_138),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_89),
.B(n_10),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_139),
.B(n_141),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_140),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_97),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_142),
.B(n_162),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_60),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_169),
.Y(n_179)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_154),
.Y(n_186)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_81),
.B1(n_77),
.B2(n_46),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_148),
.A2(n_164),
.B1(n_126),
.B2(n_121),
.Y(n_204)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_96),
.A2(n_23),
.B1(n_80),
.B2(n_44),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_153),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_102),
.Y(n_154)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_165),
.Y(n_188)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_122),
.Y(n_189)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

CKINVDCx12_ASAP7_75t_R g201 ( 
.A(n_161),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_108),
.B1(n_113),
.B2(n_84),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_44),
.B1(n_1),
.B2(n_3),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_100),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_99),
.B(n_0),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_171),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_0),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_100),
.B(n_3),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_174),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_118),
.B(n_4),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_173),
.Y(n_180)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_119),
.B(n_4),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_92),
.A2(n_128),
.B1(n_86),
.B2(n_131),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_98),
.B1(n_116),
.B2(n_105),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_86),
.B(n_4),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_4),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_95),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_159),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_189),
.B(n_203),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_131),
.C(n_122),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_194),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_128),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_134),
.B(n_130),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_205),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_141),
.B(n_130),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_6),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_106),
.Y(n_211)
);

A2O1A1O1Ixp25_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_169),
.B(n_145),
.C(n_146),
.D(n_174),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_177),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_212),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_154),
.B(n_106),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_217),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_142),
.B(n_98),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_170),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_152),
.B(n_88),
.C(n_121),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_136),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_88),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_183),
.A2(n_163),
.B1(n_140),
.B2(n_167),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_218),
.A2(n_244),
.B1(n_180),
.B2(n_203),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_163),
.B1(n_135),
.B2(n_155),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_221),
.A2(n_224),
.B1(n_240),
.B2(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_230),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_135),
.B1(n_155),
.B2(n_172),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_194),
.B(n_183),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_249),
.Y(n_258)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_193),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_145),
.B1(n_171),
.B2(n_143),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_248),
.B(n_189),
.Y(n_251)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_235),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_139),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_232),
.B(n_241),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_188),
.A2(n_160),
.B(n_158),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_233),
.A2(n_246),
.B(n_184),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_209),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_209),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_238),
.Y(n_276)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_186),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_247),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_185),
.A2(n_148),
.B1(n_137),
.B2(n_164),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_168),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_185),
.A2(n_178),
.B1(n_173),
.B2(n_157),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_206),
.A2(n_116),
.B1(n_105),
.B2(n_166),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_144),
.B(n_138),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_215),
.A2(n_147),
.B1(n_156),
.B2(n_87),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_184),
.B(n_166),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_182),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_253),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_219),
.Y(n_252)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_196),
.B1(n_214),
.B2(n_211),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_259),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_SL g257 ( 
.A1(n_233),
.A2(n_196),
.B(n_189),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_257),
.B(n_272),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_207),
.B1(n_216),
.B2(n_180),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_267),
.B1(n_277),
.B2(n_242),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_225),
.A2(n_201),
.B(n_190),
.Y(n_262)
);

AOI21x1_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_263),
.B(n_264),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_221),
.A2(n_179),
.B(n_180),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_220),
.A2(n_179),
.B(n_181),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_218),
.A2(n_181),
.B1(n_199),
.B2(n_187),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_266),
.A2(n_278),
.B1(n_242),
.B2(n_243),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_228),
.A2(n_182),
.B1(n_187),
.B2(n_126),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_191),
.C(n_201),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_275),
.C(n_222),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_245),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_231),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_226),
.C(n_249),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_240),
.A2(n_182),
.B1(n_126),
.B2(n_197),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_191),
.B1(n_200),
.B2(n_208),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_298),
.C(n_269),
.Y(n_304)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_280),
.Y(n_310)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_276),
.Y(n_281)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_238),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_282),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_241),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_283),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_287),
.Y(n_315)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_289),
.A2(n_290),
.B1(n_293),
.B2(n_297),
.Y(n_306)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_261),
.A2(n_224),
.B1(n_223),
.B2(n_230),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_291),
.A2(n_292),
.B1(n_299),
.B2(n_300),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_266),
.A2(n_245),
.B1(n_248),
.B2(n_246),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_227),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_258),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_262),
.A2(n_229),
.B(n_200),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_SL g321 ( 
.A(n_296),
.B(n_271),
.C(n_136),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_244),
.B1(n_236),
.B2(n_235),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_237),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_254),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_304),
.C(n_317),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_265),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_307),
.C(n_309),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_253),
.B(n_273),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_284),
.B(n_295),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_298),
.B(n_265),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_289),
.A2(n_263),
.B1(n_251),
.B2(n_274),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_308),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_264),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_297),
.A2(n_272),
.B1(n_278),
.B2(n_268),
.Y(n_312)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_312),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_287),
.B1(n_281),
.B2(n_293),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_316),
.A2(n_299),
.B1(n_285),
.B2(n_301),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_277),
.C(n_267),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_286),
.B(n_268),
.C(n_260),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_284),
.C(n_300),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_288),
.A2(n_260),
.B1(n_255),
.B2(n_271),
.Y(n_320)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_290),
.Y(n_322)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_316),
.B1(n_306),
.B2(n_311),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_323),
.A2(n_336),
.B1(n_302),
.B2(n_208),
.Y(n_350)
);

NAND3xp33_ASAP7_75t_SL g347 ( 
.A(n_324),
.B(n_337),
.C(n_303),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_288),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_326),
.B(n_332),
.Y(n_344)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_331),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_307),
.B(n_292),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_338),
.Y(n_348)
);

INVx13_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_335),
.Y(n_346)
);

XNOR2x2_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_301),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_320),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_333),
.A2(n_325),
.B1(n_327),
.B2(n_315),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_339),
.B(n_343),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_315),
.Y(n_342)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_325),
.A2(n_308),
.B1(n_312),
.B2(n_319),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_317),
.Y(n_345)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_345),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_347),
.A2(n_328),
.B(n_210),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_329),
.B(n_304),
.C(n_309),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_329),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_350),
.A2(n_330),
.B1(n_327),
.B2(n_324),
.Y(n_352)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_337),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_351),
.B(n_87),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_360),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_353),
.B(n_349),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_350),
.A2(n_330),
.B1(n_323),
.B2(n_334),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_361),
.Y(n_362)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_341),
.Y(n_357)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_357),
.Y(n_370)
);

NAND4xp25_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_335),
.C(n_332),
.D(n_328),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_346),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_364),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_344),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_367),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_343),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_348),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_368),
.B(n_369),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_352),
.B(n_339),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_370),
.B(n_356),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_371),
.B(n_374),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_355),
.C(n_346),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_340),
.C(n_360),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_372),
.Y(n_377)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_377),
.Y(n_381)
);

AOI322xp5_ASAP7_75t_L g378 ( 
.A1(n_373),
.A2(n_375),
.A3(n_340),
.B1(n_362),
.B2(n_342),
.C1(n_358),
.C2(n_351),
.Y(n_378)
);

AOI322xp5_ASAP7_75t_L g382 ( 
.A1(n_378),
.A2(n_379),
.A3(n_7),
.B1(n_8),
.B2(n_150),
.C1(n_161),
.C2(n_380),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_372),
.A2(n_362),
.B1(n_361),
.B2(n_210),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_382),
.A2(n_161),
.B(n_7),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_381),
.C(n_8),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_384),
.B(n_8),
.Y(n_385)
);


endmodule