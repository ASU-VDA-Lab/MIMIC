module fake_jpeg_19830_n_70 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_70);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_70;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_10),
.B(n_4),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_5),
.C(n_6),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_18),
.C(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_8),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_20),
.B(n_14),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_16),
.B(n_12),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_36),
.B(n_25),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_33)
);

OA21x2_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_38),
.B(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_9),
.Y(n_36)
);

AND2x6_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_9),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_47),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_49),
.B1(n_33),
.B2(n_35),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_56),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_49),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_39),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_46),
.C(n_42),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_45),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_61),
.C(n_55),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_40),
.B(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_57),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_53),
.Y(n_66)
);

HAxp5_ASAP7_75t_SL g68 ( 
.A(n_65),
.B(n_48),
.CON(n_68),
.SN(n_68)
);

OAI211xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_62),
.B(n_41),
.C(n_46),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_66),
.Y(n_70)
);


endmodule