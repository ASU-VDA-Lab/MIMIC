module real_aes_975_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_231;
wire n_547;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_0), .A2(n_181), .B1(n_257), .B2(n_399), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_1), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_2), .A2(n_184), .B1(n_286), .B2(n_287), .Y(n_479) );
AO22x2_ASAP7_75t_L g247 ( .A1(n_3), .A2(n_140), .B1(n_248), .B2(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g606 ( .A(n_3), .Y(n_606) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_4), .A2(n_223), .B(n_233), .C(n_608), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_5), .A2(n_178), .B1(n_372), .B2(n_375), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_6), .A2(n_52), .B1(n_577), .B2(n_578), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_7), .A2(n_208), .B1(n_282), .B2(n_293), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_8), .A2(n_127), .B1(n_365), .B2(n_407), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_9), .A2(n_56), .B1(n_286), .B2(n_294), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_10), .A2(n_83), .B1(n_358), .B2(n_575), .Y(n_574) );
OA22x2_ASAP7_75t_L g238 ( .A1(n_11), .A2(n_239), .B1(n_240), .B2(n_241), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_11), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_12), .A2(n_22), .B1(n_293), .B2(n_294), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_13), .A2(n_71), .B1(n_319), .B2(n_322), .Y(n_318) );
AO22x2_ASAP7_75t_L g261 ( .A1(n_14), .A2(n_53), .B1(n_248), .B2(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_14), .B(n_605), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_15), .A2(n_42), .B1(n_287), .B2(n_293), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_16), .A2(n_50), .B1(n_461), .B2(n_646), .Y(n_645) );
AOI22xp5_ASAP7_75t_SL g641 ( .A1(n_17), .A2(n_194), .B1(n_642), .B2(n_643), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_18), .A2(n_129), .B1(n_361), .B2(n_364), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g349 ( .A1(n_19), .A2(n_39), .B1(n_350), .B2(n_351), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_20), .A2(n_104), .B1(n_310), .B2(n_404), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_21), .A2(n_155), .B1(n_289), .B2(n_291), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_23), .A2(n_69), .B1(n_407), .B2(n_408), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_24), .A2(n_133), .B1(n_383), .B2(n_559), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_25), .A2(n_47), .B1(n_282), .B2(n_283), .Y(n_281) );
AOI222xp33_ASAP7_75t_L g243 ( .A1(n_26), .A2(n_182), .B1(n_215), .B2(n_244), .C1(n_257), .C2(n_263), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_27), .A2(n_161), .B1(n_289), .B2(n_291), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_28), .A2(n_221), .B1(n_286), .B2(n_287), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_29), .A2(n_94), .B1(n_286), .B2(n_287), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_30), .A2(n_190), .B1(n_372), .B2(n_375), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_31), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_32), .A2(n_144), .B1(n_286), .B2(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_33), .B(n_431), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_34), .A2(n_204), .B1(n_286), .B2(n_287), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_35), .A2(n_134), .B1(n_271), .B2(n_397), .Y(n_488) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_36), .A2(n_44), .B1(n_545), .B2(n_546), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_37), .A2(n_207), .B1(n_378), .B2(n_382), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_38), .A2(n_154), .B1(n_461), .B2(n_462), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_40), .A2(n_214), .B1(n_437), .B2(n_438), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_41), .A2(n_153), .B1(n_440), .B2(n_466), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g275 ( .A1(n_43), .A2(n_218), .B1(n_276), .B2(n_279), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_45), .A2(n_72), .B1(n_346), .B2(n_348), .Y(n_345) );
AO222x2_ASAP7_75t_L g613 ( .A1(n_46), .A2(n_62), .B1(n_146), .B2(n_263), .C1(n_279), .C2(n_394), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_48), .A2(n_158), .B1(n_287), .B2(n_301), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_49), .A2(n_98), .B1(n_283), .B2(n_367), .Y(n_482) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_51), .A2(n_147), .B1(n_283), .B2(n_303), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_54), .A2(n_90), .B1(n_399), .B2(n_487), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_55), .A2(n_111), .B1(n_426), .B2(n_456), .Y(n_455) );
XNOR2x2_ASAP7_75t_L g416 ( .A(n_57), .B(n_417), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_58), .A2(n_217), .B1(n_289), .B2(n_291), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_59), .A2(n_151), .B1(n_354), .B2(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_60), .B(n_431), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_61), .A2(n_200), .B1(n_279), .B2(n_394), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_63), .A2(n_65), .B1(n_244), .B2(n_487), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_64), .A2(n_126), .B1(n_283), .B2(n_303), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_66), .A2(n_121), .B1(n_441), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_67), .A2(n_175), .B1(n_404), .B2(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g248 ( .A(n_68), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_70), .A2(n_201), .B1(n_368), .B2(n_379), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_73), .A2(n_131), .B1(n_282), .B2(n_283), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_74), .B(n_426), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_75), .A2(n_137), .B1(n_293), .B2(n_294), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_76), .A2(n_114), .B1(n_364), .B2(n_638), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_77), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_78), .B(n_580), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_79), .A2(n_92), .B1(n_441), .B2(n_634), .Y(n_633) );
AO22x1_ASAP7_75t_L g419 ( .A1(n_80), .A2(n_112), .B1(n_420), .B2(n_421), .Y(n_419) );
INVx1_ASAP7_75t_SL g253 ( .A(n_81), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_81), .B(n_97), .Y(n_607) );
INVx2_ASAP7_75t_L g232 ( .A(n_82), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_84), .A2(n_174), .B1(n_325), .B2(n_327), .Y(n_324) );
XOR2x2_ASAP7_75t_L g552 ( .A(n_85), .B(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_86), .A2(n_160), .B1(n_361), .B2(n_443), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_87), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_88), .A2(n_99), .B1(n_526), .B2(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_89), .A2(n_102), .B1(n_589), .B2(n_591), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_91), .A2(n_193), .B1(n_271), .B2(n_397), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_93), .B(n_343), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_95), .A2(n_177), .B1(n_282), .B2(n_283), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_96), .B(n_263), .Y(n_502) );
AO22x2_ASAP7_75t_L g255 ( .A1(n_97), .A2(n_149), .B1(n_248), .B2(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_100), .B(n_315), .Y(n_314) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_101), .A2(n_119), .B1(n_429), .B2(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_103), .A2(n_170), .B1(n_279), .B2(n_394), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_105), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_106), .A2(n_187), .B1(n_367), .B2(n_368), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_107), .A2(n_113), .B1(n_289), .B2(n_620), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_108), .Y(n_392) );
INVx1_ASAP7_75t_L g254 ( .A(n_109), .Y(n_254) );
AOI22xp33_ASAP7_75t_SL g402 ( .A1(n_110), .A2(n_157), .B1(n_289), .B2(n_305), .Y(n_402) );
XNOR2xp5_ASAP7_75t_L g515 ( .A(n_115), .B(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_116), .A2(n_186), .B1(n_319), .B2(n_397), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_117), .A2(n_213), .B1(n_305), .B2(n_307), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_118), .B(n_431), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_120), .A2(n_124), .B1(n_271), .B2(n_397), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_122), .A2(n_172), .B1(n_301), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g396 ( .A1(n_123), .A2(n_210), .B1(n_271), .B2(n_397), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_125), .A2(n_138), .B1(n_289), .B2(n_291), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_128), .A2(n_171), .B1(n_583), .B2(n_586), .Y(n_582) );
XNOR2x1_ASAP7_75t_L g499 ( .A(n_130), .B(n_500), .Y(n_499) );
AO22x1_ASAP7_75t_L g423 ( .A1(n_132), .A2(n_205), .B1(n_424), .B2(n_426), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_135), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_136), .A2(n_203), .B1(n_267), .B2(n_271), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_139), .A2(n_165), .B1(n_468), .B2(n_469), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_141), .A2(n_183), .B1(n_354), .B2(n_356), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_142), .A2(n_202), .B1(n_440), .B2(n_441), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_143), .A2(n_180), .B1(n_434), .B2(n_435), .Y(n_433) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_145), .A2(n_197), .B1(n_352), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_148), .A2(n_185), .B1(n_548), .B2(n_549), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_150), .A2(n_162), .B1(n_594), .B2(n_595), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_152), .A2(n_196), .B1(n_276), .B2(n_279), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_156), .A2(n_189), .B1(n_538), .B2(n_539), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_159), .B(n_431), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_163), .A2(n_610), .B1(n_611), .B2(n_625), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_163), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_164), .Y(n_648) );
AO22x2_ASAP7_75t_L g476 ( .A1(n_166), .A2(n_477), .B1(n_489), .B2(n_490), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_166), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_167), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g602 ( .A(n_167), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_168), .A2(n_198), .B1(n_244), .B2(n_257), .Y(n_565) );
XOR2x2_ASAP7_75t_L g569 ( .A(n_169), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g228 ( .A(n_173), .Y(n_228) );
AND2x2_ASAP7_75t_R g627 ( .A(n_173), .B(n_602), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_176), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_179), .A2(n_339), .B1(n_340), .B2(n_384), .Y(n_338) );
INVx1_ASAP7_75t_L g384 ( .A(n_179), .Y(n_384) );
INVxp67_ASAP7_75t_L g230 ( .A(n_188), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_191), .A2(n_206), .B1(n_325), .B2(n_352), .Y(n_644) );
INVx1_ASAP7_75t_L g410 ( .A(n_192), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_195), .A2(n_220), .B1(n_244), .B2(n_257), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_199), .A2(n_209), .B1(n_286), .B2(n_287), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_211), .A2(n_216), .B1(n_244), .B2(n_487), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_212), .Y(n_524) );
OA22x2_ASAP7_75t_L g295 ( .A1(n_219), .A2(n_296), .B1(n_297), .B2(n_331), .Y(n_295) );
INVx1_ASAP7_75t_L g331 ( .A(n_219), .Y(n_331) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_225), .Y(n_224) );
AND2x4_ASAP7_75t_SL g225 ( .A(n_226), .B(n_229), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g652 ( .A(n_227), .B(n_229), .Y(n_652) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_228), .B(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_494), .B1(n_597), .B2(n_598), .C(n_599), .Y(n_233) );
INVx1_ASAP7_75t_L g597 ( .A(n_234), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_413), .B1(n_414), .B2(n_493), .Y(n_234) );
INVx1_ASAP7_75t_L g493 ( .A(n_235), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_334), .B1(n_335), .B2(n_412), .Y(n_235) );
INVx1_ASAP7_75t_L g412 ( .A(n_236), .Y(n_412) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OAI22xp33_ASAP7_75t_SL g237 ( .A1(n_238), .A2(n_295), .B1(n_332), .B2(n_333), .Y(n_237) );
INVx1_ASAP7_75t_L g332 ( .A(n_238), .Y(n_332) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2x1_ASAP7_75t_L g241 ( .A(n_242), .B(n_280), .Y(n_241) );
NAND3xp33_ASAP7_75t_L g242 ( .A(n_243), .B(n_266), .C(n_275), .Y(n_242) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_250), .Y(n_244) );
AND2x4_ASAP7_75t_L g358 ( .A(n_245), .B(n_250), .Y(n_358) );
AND2x2_ASAP7_75t_L g399 ( .A(n_245), .B(n_250), .Y(n_399) );
INVxp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x4_ASAP7_75t_L g260 ( .A(n_246), .B(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g264 ( .A(n_246), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g272 ( .A(n_247), .B(n_270), .Y(n_272) );
AND2x2_ASAP7_75t_L g278 ( .A(n_247), .B(n_261), .Y(n_278) );
INVx1_ASAP7_75t_L g249 ( .A(n_248), .Y(n_249) );
OAI22x1_ASAP7_75t_L g251 ( .A1(n_248), .A2(n_252), .B1(n_253), .B2(n_254), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_248), .Y(n_252) );
INVx1_ASAP7_75t_L g256 ( .A(n_248), .Y(n_256) );
INVx2_ASAP7_75t_L g262 ( .A(n_248), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_250), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g267 ( .A(n_250), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g317 ( .A(n_250), .B(n_264), .Y(n_317) );
AND2x4_ASAP7_75t_L g323 ( .A(n_250), .B(n_268), .Y(n_323) );
AND2x2_ASAP7_75t_L g397 ( .A(n_250), .B(n_268), .Y(n_397) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_255), .Y(n_250) );
INVx2_ASAP7_75t_L g259 ( .A(n_251), .Y(n_259) );
AND2x2_ASAP7_75t_L g273 ( .A(n_251), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_251), .Y(n_277) );
AND2x2_ASAP7_75t_L g258 ( .A(n_255), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g274 ( .A(n_255), .Y(n_274) );
BUFx2_ASAP7_75t_L g290 ( .A(n_255), .Y(n_290) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
AND2x6_ASAP7_75t_L g287 ( .A(n_258), .B(n_264), .Y(n_287) );
AND2x2_ASAP7_75t_L g291 ( .A(n_258), .B(n_272), .Y(n_291) );
AND2x2_ASAP7_75t_L g306 ( .A(n_258), .B(n_272), .Y(n_306) );
AND2x4_ASAP7_75t_L g355 ( .A(n_258), .B(n_260), .Y(n_355) );
AND2x2_ASAP7_75t_L g381 ( .A(n_258), .B(n_264), .Y(n_381) );
AND2x2_ASAP7_75t_L g487 ( .A(n_258), .B(n_260), .Y(n_487) );
AND2x2_ASAP7_75t_SL g620 ( .A(n_258), .B(n_272), .Y(n_620) );
AND2x4_ASAP7_75t_L g284 ( .A(n_259), .B(n_274), .Y(n_284) );
AND2x4_ASAP7_75t_L g279 ( .A(n_260), .B(n_273), .Y(n_279) );
AND2x2_ASAP7_75t_L g293 ( .A(n_260), .B(n_284), .Y(n_293) );
AND2x4_ASAP7_75t_L g301 ( .A(n_260), .B(n_284), .Y(n_301) );
AND2x2_ASAP7_75t_L g326 ( .A(n_260), .B(n_273), .Y(n_326) );
INVx1_ASAP7_75t_L g265 ( .A(n_261), .Y(n_265) );
INVx1_ASAP7_75t_L g270 ( .A(n_261), .Y(n_270) );
INVx2_ASAP7_75t_SL g391 ( .A(n_263), .Y(n_391) );
AND2x2_ASAP7_75t_L g282 ( .A(n_264), .B(n_273), .Y(n_282) );
AND2x2_ASAP7_75t_L g294 ( .A(n_264), .B(n_284), .Y(n_294) );
AND2x2_ASAP7_75t_L g303 ( .A(n_264), .B(n_273), .Y(n_303) );
AND2x4_ASAP7_75t_L g312 ( .A(n_264), .B(n_284), .Y(n_312) );
AND2x4_ASAP7_75t_L g363 ( .A(n_264), .B(n_273), .Y(n_363) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AND2x6_ASAP7_75t_L g286 ( .A(n_272), .B(n_284), .Y(n_286) );
AND2x2_ASAP7_75t_L g321 ( .A(n_272), .B(n_273), .Y(n_321) );
AND2x4_ASAP7_75t_L g370 ( .A(n_272), .B(n_284), .Y(n_370) );
AND2x2_ASAP7_75t_SL g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g329 ( .A(n_277), .B(n_278), .Y(n_329) );
AND2x2_ASAP7_75t_SL g394 ( .A(n_277), .B(n_278), .Y(n_394) );
AND2x4_ASAP7_75t_L g283 ( .A(n_278), .B(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g289 ( .A(n_278), .B(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g308 ( .A(n_278), .B(n_290), .Y(n_308) );
AND2x4_ASAP7_75t_L g365 ( .A(n_278), .B(n_284), .Y(n_365) );
NAND4xp25_ASAP7_75t_L g280 ( .A(n_281), .B(n_285), .C(n_288), .D(n_292), .Y(n_280) );
INVx2_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NOR2xp67_ASAP7_75t_L g297 ( .A(n_298), .B(n_313), .Y(n_297) );
NAND3xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_304), .C(n_309), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_301), .Y(n_383) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_301), .Y(n_404) );
BUFx3_ASAP7_75t_L g438 ( .A(n_301), .Y(n_438) );
BUFx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g374 ( .A(n_306), .Y(n_374) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_306), .Y(n_634) );
BUFx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx5_ASAP7_75t_SL g376 ( .A(n_308), .Y(n_376) );
INVx3_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx4_ASAP7_75t_L g367 ( .A(n_311), .Y(n_367) );
INVx2_ASAP7_75t_SL g437 ( .A(n_311), .Y(n_437) );
INVx2_ASAP7_75t_L g473 ( .A(n_311), .Y(n_473) );
INVx2_ASAP7_75t_SL g545 ( .A(n_311), .Y(n_545) );
INVx3_ASAP7_75t_L g559 ( .A(n_311), .Y(n_559) );
INVx8_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND4xp25_ASAP7_75t_L g313 ( .A(n_314), .B(n_318), .C(n_324), .D(n_330), .Y(n_313) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g344 ( .A(n_316), .Y(n_344) );
INVx4_ASAP7_75t_SL g431 ( .A(n_316), .Y(n_431) );
INVx3_ASAP7_75t_SL g453 ( .A(n_316), .Y(n_453) );
INVx6_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx4_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g420 ( .A(n_320), .Y(n_420) );
INVx1_ASAP7_75t_L g527 ( .A(n_320), .Y(n_527) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_321), .Y(n_347) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_321), .Y(n_461) );
BUFx2_ASAP7_75t_SL g348 ( .A(n_322), .Y(n_348) );
BUFx6f_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g422 ( .A(n_323), .Y(n_422) );
BUFx3_ASAP7_75t_L g462 ( .A(n_323), .Y(n_462) );
INVx1_ASAP7_75t_L g647 ( .A(n_323), .Y(n_647) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_325), .Y(n_350) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g425 ( .A(n_326), .Y(n_425) );
BUFx3_ASAP7_75t_L g456 ( .A(n_326), .Y(n_456) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_327), .Y(n_578) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g352 ( .A(n_328), .Y(n_352) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx12f_ASAP7_75t_L g426 ( .A(n_329), .Y(n_426) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
OAI22x1_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_385), .B2(n_411), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_359), .Y(n_340) );
NAND4xp25_ASAP7_75t_SL g341 ( .A(n_342), .B(n_345), .C(n_349), .D(n_353), .Y(n_341) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx4f_ASAP7_75t_SL g533 ( .A(n_354), .Y(n_533) );
BUFx2_ASAP7_75t_L g575 ( .A(n_354), .Y(n_575) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g459 ( .A(n_355), .Y(n_459) );
BUFx2_ASAP7_75t_L g642 ( .A(n_355), .Y(n_642) );
INVx2_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g429 ( .A(n_357), .Y(n_429) );
OAI22xp33_ASAP7_75t_L g530 ( .A1(n_357), .A2(n_531), .B1(n_532), .B2(n_534), .Y(n_530) );
INVx1_ASAP7_75t_L g643 ( .A(n_357), .Y(n_643) );
INVx6_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND4xp25_ASAP7_75t_L g359 ( .A(n_360), .B(n_366), .C(n_371), .D(n_377), .Y(n_359) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g538 ( .A(n_362), .Y(n_538) );
INVx1_ASAP7_75t_SL g594 ( .A(n_362), .Y(n_594) );
INVx3_ASAP7_75t_L g638 ( .A(n_362), .Y(n_638) );
INVx6_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx3_ASAP7_75t_L g407 ( .A(n_363), .Y(n_407) );
BUFx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx3_ASAP7_75t_L g408 ( .A(n_365), .Y(n_408) );
INVx2_ASAP7_75t_L g444 ( .A(n_365), .Y(n_444) );
BUFx2_ASAP7_75t_SL g539 ( .A(n_365), .Y(n_539) );
BUFx2_ASAP7_75t_SL g595 ( .A(n_365), .Y(n_595) );
INVx2_ASAP7_75t_L g590 ( .A(n_367), .Y(n_590) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g435 ( .A(n_369), .Y(n_435) );
INVx2_ASAP7_75t_L g469 ( .A(n_369), .Y(n_469) );
INVx1_ASAP7_75t_SL g546 ( .A(n_369), .Y(n_546) );
INVx2_ASAP7_75t_L g586 ( .A(n_369), .Y(n_586) );
INVx8_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g440 ( .A(n_374), .Y(n_440) );
INVx2_ASAP7_75t_L g542 ( .A(n_374), .Y(n_542) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx3_ASAP7_75t_L g441 ( .A(n_376), .Y(n_441) );
INVx2_ASAP7_75t_L g466 ( .A(n_376), .Y(n_466) );
BUFx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g434 ( .A(n_380), .Y(n_434) );
INVx2_ASAP7_75t_SL g548 ( .A(n_380), .Y(n_548) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g468 ( .A(n_381), .Y(n_468) );
BUFx2_ASAP7_75t_L g585 ( .A(n_381), .Y(n_585) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g550 ( .A(n_383), .Y(n_550) );
INVx1_ASAP7_75t_SL g411 ( .A(n_385), .Y(n_411) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
XOR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_410), .Y(n_387) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_400), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_395), .Y(n_389) );
OAI21xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_392), .B(n_393), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_401), .B(n_405), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx2_ASAP7_75t_L g592 ( .A(n_404), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_409), .Y(n_405) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_445), .B1(n_446), .B2(n_492), .Y(n_414) );
INVx1_ASAP7_75t_L g492 ( .A(n_415), .Y(n_492) );
BUFx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_432), .Y(n_417) );
NOR3xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_423), .C(n_427), .Y(n_418) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx2_ASAP7_75t_L g529 ( .A(n_422), .Y(n_529) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g562 ( .A(n_425), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_428), .B(n_430), .Y(n_427) );
AND4x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_436), .C(n_439), .D(n_442), .Y(n_432) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22x1_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_475), .B1(n_476), .B2(n_491), .Y(n_447) );
INVx2_ASAP7_75t_L g491 ( .A(n_448), .Y(n_491) );
XNOR2x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_474), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_463), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_457), .Y(n_450) );
OAI21xp33_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_454), .B(n_455), .Y(n_451) );
OAI221xp5_ASAP7_75t_L g518 ( .A1(n_452), .A2(n_519), .B1(n_520), .B2(n_521), .C(n_522), .Y(n_518) );
INVx2_ASAP7_75t_L g580 ( .A(n_452), .Y(n_580) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g521 ( .A(n_456), .Y(n_521) );
BUFx6f_ASAP7_75t_SL g577 ( .A(n_456), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
BUFx6f_ASAP7_75t_SL g573 ( .A(n_462), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_470), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g490 ( .A(n_477), .Y(n_490) );
NOR2xp67_ASAP7_75t_L g477 ( .A(n_478), .B(n_483), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .C(n_481), .D(n_482), .Y(n_478) );
NAND4xp25_ASAP7_75t_SL g483 ( .A(n_484), .B(n_485), .C(n_486), .D(n_488), .Y(n_483) );
INVx1_ASAP7_75t_L g598 ( .A(n_494), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_511), .B2(n_596), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_506), .Y(n_500) );
NAND4xp25_ASAP7_75t_SL g501 ( .A(n_502), .B(n_503), .C(n_504), .D(n_505), .Y(n_501) );
NAND4xp25_ASAP7_75t_SL g506 ( .A(n_507), .B(n_508), .C(n_509), .D(n_510), .Y(n_506) );
INVxp67_ASAP7_75t_L g596 ( .A(n_511), .Y(n_596) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OA22x2_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B1(n_568), .B2(n_569), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_551), .B1(n_552), .B2(n_567), .Y(n_514) );
INVx1_ASAP7_75t_L g567 ( .A(n_515), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_535), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_523), .C(n_530), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_528), .B2(n_529), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_543), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_547), .Y(n_543) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NOR3xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_560), .C(n_564), .Y(n_553) );
NAND4xp25_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .C(n_557), .D(n_558), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx4_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_581), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .C(n_576), .D(n_579), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g581 ( .A(n_582), .B(n_587), .C(n_588), .D(n_593), .Y(n_581) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_601), .B(n_604), .Y(n_651) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
OAI222xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_626), .B1(n_628), .B2(n_648), .C1(n_649), .C2(n_652), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2x1_ASAP7_75t_L g611 ( .A(n_612), .B(n_617), .Y(n_611) );
NOR2x1_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_622), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
XNOR2x1_ASAP7_75t_L g630 ( .A(n_631), .B(n_648), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_639), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .C(n_636), .D(n_637), .Y(n_632) );
NAND4xp25_ASAP7_75t_SL g639 ( .A(n_640), .B(n_641), .C(n_644), .D(n_645), .Y(n_639) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
CKINVDCx6p67_ASAP7_75t_R g650 ( .A(n_651), .Y(n_650) );
endmodule