module fake_jpeg_6408_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_241;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_38),
.CON(n_51),
.SN(n_51)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_30),
.Y(n_53)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_16),
.A2(n_17),
.B1(n_30),
.B2(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_29),
.B1(n_28),
.B2(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_56),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_16),
.B1(n_29),
.B2(n_28),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_24),
.B(n_22),
.Y(n_71)
);

AO22x1_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_16),
.B1(n_21),
.B2(n_23),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_41),
.B1(n_39),
.B2(n_23),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_21),
.B1(n_23),
.B2(n_27),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_55),
.B1(n_24),
.B2(n_22),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_19),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_22),
.B1(n_29),
.B2(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_66),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_15),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_63),
.C(n_1),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_19),
.Y(n_72)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_47),
.B1(n_51),
.B2(n_57),
.Y(n_89)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_81),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_48),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_53),
.B(n_25),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_46),
.B1(n_61),
.B2(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_34),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_46),
.Y(n_95)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_47),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_87),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_98),
.B1(n_99),
.B2(n_75),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_104),
.B(n_71),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_103),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_61),
.B1(n_46),
.B2(n_60),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_102),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_61),
.B1(n_50),
.B2(n_52),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_90),
.B1(n_65),
.B2(n_87),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_34),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_54),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_125),
.B1(n_86),
.B2(n_101),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_106),
.A2(n_79),
.B1(n_69),
.B2(n_85),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_113),
.B1(n_79),
.B2(n_65),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_79),
.B1(n_69),
.B2(n_85),
.Y(n_113)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_84),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_88),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_121),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_73),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_78),
.B1(n_83),
.B2(n_76),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_99),
.B1(n_98),
.B2(n_87),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_104),
.B(n_92),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_70),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_130),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_105),
.B(n_54),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_88),
.A2(n_70),
.B(n_78),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_34),
.B(n_31),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_140),
.B1(n_115),
.B2(n_116),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_154),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_77),
.Y(n_184)
);

NAND2xp33_ASAP7_75t_SL g179 ( 
.A(n_137),
.B(n_54),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_155),
.B(n_121),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_86),
.B1(n_97),
.B2(n_100),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_117),
.B1(n_109),
.B2(n_124),
.Y(n_176)
);

AO22x1_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_97),
.B1(n_66),
.B2(n_101),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_146),
.B(n_156),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_66),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_114),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_148),
.B(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_125),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_157),
.C(n_131),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_110),
.A2(n_97),
.B1(n_107),
.B2(n_80),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_107),
.B(n_77),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_128),
.C(n_132),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_42),
.B1(n_23),
.B2(n_62),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_162),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_120),
.C(n_130),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_184),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_169),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_120),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_166),
.B(n_168),
.Y(n_195)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_156),
.C(n_158),
.Y(n_196)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_133),
.B1(n_117),
.B2(n_62),
.Y(n_172)
);

AO22x1_ASAP7_75t_SL g202 ( 
.A1(n_172),
.A2(n_137),
.B1(n_142),
.B2(n_145),
.Y(n_202)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_182),
.Y(n_192)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_175),
.A2(n_176),
.B(n_179),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_178),
.A2(n_183),
.B1(n_154),
.B2(n_150),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_34),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_196),
.C(n_199),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_135),
.B1(n_170),
.B2(n_172),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_187),
.A2(n_190),
.B1(n_202),
.B2(n_204),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_155),
.B1(n_138),
.B2(n_134),
.Y(n_190)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_207),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_148),
.C(n_141),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_166),
.A2(n_145),
.B1(n_142),
.B2(n_137),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_152),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_169),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_31),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_208),
.Y(n_214)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_31),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_223),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_112),
.Y(n_213)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_216),
.A2(n_227),
.B(n_228),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_192),
.A2(n_167),
.B1(n_162),
.B2(n_173),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_217),
.A2(n_209),
.B1(n_222),
.B2(n_219),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_167),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_164),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_183),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_206),
.C(n_196),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_112),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_194),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_194),
.B(n_112),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_232),
.C(n_221),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_197),
.B1(n_201),
.B2(n_188),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_233),
.B1(n_210),
.B2(n_215),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_192),
.C(n_185),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_190),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_235),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_217),
.B(n_208),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_189),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_245),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_189),
.B(n_204),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_241),
.A2(n_240),
.B(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_159),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_183),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_250),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_209),
.B1(n_201),
.B2(n_211),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_249),
.A2(n_67),
.B1(n_21),
.B2(n_2),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_174),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_252),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_67),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_232),
.B(n_214),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_260),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_256),
.A2(n_236),
.B(n_239),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_237),
.A2(n_221),
.B(n_159),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_258),
.B(n_259),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_195),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_230),
.B(n_42),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_234),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_239),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_241),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_263),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_270),
.B(n_272),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_259),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_20),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_245),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_67),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_255),
.B(n_9),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_255),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_281),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_20),
.B(n_1),
.Y(n_291)
);

AOI221xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_283),
.B1(n_10),
.B2(n_14),
.C(n_12),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_49),
.B(n_20),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_12),
.A3(n_11),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_21),
.B(n_1),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_285),
.Y(n_295)
);

AOI221xp5_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_267),
.B1(n_265),
.B2(n_263),
.C(n_271),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_289),
.A3(n_290),
.B1(n_291),
.B2(n_2),
.C1(n_4),
.C2(n_5),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_20),
.A3(n_11),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_278),
.C(n_277),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.C(n_296),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_0),
.B(n_1),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_5),
.B(n_6),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_279),
.C2(n_267),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_295),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_297),
.C(n_7),
.Y(n_300)
);


endmodule