module fake_aes_6758_n_783 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_39, n_783);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_39;
output n_783;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_223;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g95 ( .A(n_36), .Y(n_95) );
BUFx6f_ASAP7_75t_L g96 ( .A(n_76), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_36), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_48), .Y(n_98) );
BUFx2_ASAP7_75t_L g99 ( .A(n_49), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_15), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_60), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_74), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_59), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_65), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_10), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_47), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_58), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_66), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_33), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_79), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_83), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_69), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_53), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_11), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_29), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_6), .Y(n_116) );
CKINVDCx14_ASAP7_75t_R g117 ( .A(n_20), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_85), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_82), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_55), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_31), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_87), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_75), .Y(n_124) );
INVx2_ASAP7_75t_SL g125 ( .A(n_57), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_51), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_88), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_84), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_80), .Y(n_129) );
INVx2_ASAP7_75t_SL g130 ( .A(n_35), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_17), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_94), .Y(n_132) );
CKINVDCx12_ASAP7_75t_R g133 ( .A(n_56), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_7), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_27), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_2), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_4), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_68), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_33), .Y(n_139) );
BUFx12f_ASAP7_75t_L g140 ( .A(n_125), .Y(n_140) );
NOR2xp33_ASAP7_75t_SL g141 ( .A(n_103), .B(n_39), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_99), .B(n_0), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_98), .Y(n_143) );
BUFx12f_ASAP7_75t_L g144 ( .A(n_125), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_99), .B(n_1), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_125), .B(n_1), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_96), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_130), .B(n_2), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_130), .B(n_3), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_105), .Y(n_151) );
BUFx8_ASAP7_75t_SL g152 ( .A(n_100), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_96), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_105), .B(n_3), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_108), .Y(n_155) );
BUFx12f_ASAP7_75t_L g156 ( .A(n_96), .Y(n_156) );
INVxp67_ASAP7_75t_L g157 ( .A(n_130), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_96), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_117), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_96), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_95), .B(n_4), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_115), .B(n_5), .Y(n_162) );
AO22x2_ASAP7_75t_L g163 ( .A1(n_142), .A2(n_95), .B1(n_97), .B2(n_116), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_151), .B(n_115), .Y(n_164) );
BUFx10_ASAP7_75t_L g165 ( .A(n_159), .Y(n_165) );
OAI22xp33_ASAP7_75t_L g166 ( .A1(n_151), .A2(n_109), .B1(n_97), .B2(n_116), .Y(n_166) );
AO22x2_ASAP7_75t_L g167 ( .A1(n_142), .A2(n_136), .B1(n_102), .B2(n_104), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_148), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_142), .A2(n_139), .B1(n_114), .B2(n_137), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_142), .A2(n_121), .B1(n_135), .B2(n_134), .Y(n_171) );
BUFx10_ASAP7_75t_L g172 ( .A(n_159), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_142), .A2(n_122), .B1(n_131), .B2(n_136), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_140), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_151), .B(n_101), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_154), .B(n_106), .Y(n_177) );
OAI22xp33_ASAP7_75t_SL g178 ( .A1(n_141), .A2(n_119), .B1(n_102), .B2(n_104), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_155), .Y(n_179) );
BUFx6f_ASAP7_75t_SL g180 ( .A(n_142), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_142), .A2(n_138), .B1(n_128), .B2(n_133), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_142), .A2(n_133), .B1(n_119), .B2(n_118), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_154), .A2(n_118), .B1(n_110), .B2(n_127), .Y(n_184) );
INVxp67_ASAP7_75t_SL g185 ( .A(n_145), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_154), .A2(n_98), .B1(n_110), .B2(n_127), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g188 ( .A1(n_145), .A2(n_111), .B1(n_124), .B2(n_123), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
OAI22xp33_ASAP7_75t_SL g190 ( .A1(n_141), .A2(n_111), .B1(n_112), .B2(n_124), .Y(n_190) );
AO22x2_ASAP7_75t_L g191 ( .A1(n_148), .A2(n_112), .B1(n_123), .B2(n_108), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_157), .B(n_107), .Y(n_192) );
OAI22xp33_ASAP7_75t_SL g193 ( .A1(n_141), .A2(n_132), .B1(n_129), .B2(n_126), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_157), .B(n_108), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_155), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_154), .A2(n_120), .B1(n_113), .B2(n_7), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_157), .B(n_5), .Y(n_197) );
CKINVDCx6p67_ASAP7_75t_R g198 ( .A(n_162), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_148), .A2(n_6), .B1(n_8), .B2(n_9), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_140), .B(n_40), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_162), .B(n_8), .Y(n_201) );
NOR2xp33_ASAP7_75t_SL g202 ( .A(n_162), .B(n_41), .Y(n_202) );
AO22x2_ASAP7_75t_L g203 ( .A1(n_148), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_148), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_162), .B(n_12), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_145), .B(n_12), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_156), .Y(n_207) );
OAI22xp33_ASAP7_75t_L g208 ( .A1(n_161), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_185), .B(n_143), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_168), .B(n_143), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_168), .B(n_143), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_168), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_175), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_169), .A2(n_146), .B(n_149), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_164), .B(n_163), .Y(n_215) );
INVx4_ASAP7_75t_SL g216 ( .A(n_180), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_163), .B(n_161), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_175), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_179), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_174), .B(n_140), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_163), .B(n_161), .Y(n_221) );
NOR2xp67_ASAP7_75t_L g222 ( .A(n_187), .B(n_140), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_182), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_182), .Y(n_224) );
XOR2xp5_ASAP7_75t_L g225 ( .A(n_181), .B(n_152), .Y(n_225) );
INVx1_ASAP7_75t_SL g226 ( .A(n_198), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_195), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_174), .Y(n_228) );
BUFx3_ASAP7_75t_L g229 ( .A(n_191), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_195), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_189), .Y(n_231) );
HAxp5_ASAP7_75t_SL g232 ( .A(n_196), .B(n_152), .CON(n_232), .SN(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_198), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_165), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_204), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_191), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_165), .B(n_144), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_177), .B(n_149), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_191), .Y(n_239) );
INVxp67_ASAP7_75t_L g240 ( .A(n_180), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_188), .B(n_146), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_167), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_207), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_167), .Y(n_244) );
INVxp33_ASAP7_75t_L g245 ( .A(n_176), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_206), .B(n_149), .Y(n_246) );
INVx2_ASAP7_75t_SL g247 ( .A(n_207), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_165), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_167), .B(n_146), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_172), .B(n_144), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_203), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_203), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_203), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_172), .B(n_155), .Y(n_254) );
NOR2xp67_ASAP7_75t_L g255 ( .A(n_183), .B(n_144), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_207), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_172), .B(n_155), .Y(n_257) );
XOR2xp5_ASAP7_75t_L g258 ( .A(n_170), .B(n_13), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_171), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_194), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_194), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_194), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_199), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_205), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_197), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_205), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_201), .B(n_155), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_192), .B(n_144), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_208), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_178), .A2(n_160), .B(n_153), .Y(n_270) );
BUFx5_ASAP7_75t_L g271 ( .A(n_190), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_246), .B(n_173), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_246), .B(n_184), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_209), .B(n_188), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_227), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_209), .B(n_238), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_209), .B(n_186), .Y(n_277) );
INVx4_ASAP7_75t_L g278 ( .A(n_229), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_229), .B(n_200), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_229), .B(n_200), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_212), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_243), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_212), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_254), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_238), .B(n_193), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_217), .B(n_166), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_231), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_245), .B(n_166), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_231), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_247), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_217), .B(n_202), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_221), .B(n_156), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_269), .A2(n_208), .B1(n_156), .B2(n_160), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_215), .B(n_156), .Y(n_294) );
INVx4_ASAP7_75t_L g295 ( .A(n_216), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_231), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_235), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_271), .B(n_147), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_247), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_254), .B(n_153), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_215), .B(n_14), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_227), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_216), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_257), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_248), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_263), .B(n_16), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_270), .A2(n_160), .B(n_153), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_257), .B(n_153), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_263), .B(n_16), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_227), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_213), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_226), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_249), .B(n_17), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_247), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_264), .B(n_153), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_226), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_264), .B(n_266), .Y(n_317) );
BUFx4_ASAP7_75t_SL g318 ( .A(n_234), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_266), .B(n_160), .Y(n_319) );
AND2x2_ASAP7_75t_SL g320 ( .A(n_251), .B(n_160), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_249), .B(n_18), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_241), .B(n_18), .Y(n_322) );
AND2x2_ASAP7_75t_SL g323 ( .A(n_251), .B(n_147), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_213), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_235), .Y(n_325) );
AND2x2_ASAP7_75t_SL g326 ( .A(n_278), .B(n_252), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_284), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_318), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_278), .B(n_216), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_276), .B(n_214), .Y(n_330) );
AND2x6_ASAP7_75t_L g331 ( .A(n_291), .B(n_242), .Y(n_331) );
INVx2_ASAP7_75t_SL g332 ( .A(n_278), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_275), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_311), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_295), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_276), .B(n_214), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_286), .B(n_241), .Y(n_337) );
AND2x6_ASAP7_75t_L g338 ( .A(n_291), .B(n_244), .Y(n_338) );
OR2x6_ASAP7_75t_L g339 ( .A(n_278), .B(n_244), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_273), .B(n_267), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_284), .Y(n_341) );
NOR2xp33_ASAP7_75t_SL g342 ( .A(n_278), .B(n_295), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_286), .B(n_269), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_274), .B(n_271), .Y(n_344) );
BUFx4f_ASAP7_75t_L g345 ( .A(n_303), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_278), .Y(n_346) );
OR2x6_ASAP7_75t_L g347 ( .A(n_295), .B(n_252), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_311), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_273), .B(n_259), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_295), .Y(n_350) );
NOR2xp67_ASAP7_75t_L g351 ( .A(n_295), .B(n_253), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_305), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_273), .B(n_233), .Y(n_353) );
BUFx4f_ASAP7_75t_L g354 ( .A(n_303), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_275), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_311), .Y(n_356) );
NOR2x1_ASAP7_75t_L g357 ( .A(n_295), .B(n_236), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_272), .B(n_267), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_304), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_304), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_335), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_341), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_341), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_339), .Y(n_364) );
BUFx4f_ASAP7_75t_L g365 ( .A(n_329), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_330), .B(n_274), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_334), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_329), .Y(n_368) );
INVx4_ASAP7_75t_L g369 ( .A(n_329), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_334), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_329), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_333), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_330), .B(n_277), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_348), .B(n_303), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_339), .Y(n_375) );
INVx4_ASAP7_75t_L g376 ( .A(n_329), .Y(n_376) );
INVx5_ASAP7_75t_L g377 ( .A(n_339), .Y(n_377) );
AND2x6_ASAP7_75t_L g378 ( .A(n_348), .B(n_291), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_335), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_346), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
INVx6_ASAP7_75t_L g382 ( .A(n_335), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_349), .B(n_272), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_349), .A2(n_285), .B1(n_321), .B2(n_313), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_339), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_335), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_356), .B(n_311), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_339), .Y(n_388) );
INVx2_ASAP7_75t_SL g389 ( .A(n_345), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_335), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_356), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_361), .Y(n_392) );
BUFx2_ASAP7_75t_L g393 ( .A(n_364), .Y(n_393) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_361), .Y(n_394) );
CKINVDCx11_ASAP7_75t_R g395 ( .A(n_362), .Y(n_395) );
BUFx12f_ASAP7_75t_L g396 ( .A(n_369), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_383), .A2(n_353), .B1(n_358), .B2(n_340), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_384), .A2(n_293), .B1(n_305), .B2(n_360), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_372), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_384), .A2(n_293), .B1(n_360), .B2(n_312), .Y(n_400) );
OAI21xp5_ASAP7_75t_SL g401 ( .A1(n_364), .A2(n_225), .B(n_258), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_372), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_361), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_383), .A2(n_353), .B1(n_358), .B2(n_340), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_367), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_362), .Y(n_406) );
INVx3_ASAP7_75t_SL g407 ( .A(n_377), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_361), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_372), .Y(n_409) );
BUFx8_ASAP7_75t_L g410 ( .A(n_364), .Y(n_410) );
BUFx6f_ASAP7_75t_SL g411 ( .A(n_387), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_367), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_378), .A2(n_358), .B1(n_340), .B2(n_338), .Y(n_413) );
BUFx2_ASAP7_75t_SL g414 ( .A(n_377), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_377), .A2(n_313), .B1(n_321), .B2(n_327), .Y(n_415) );
BUFx12f_ASAP7_75t_L g416 ( .A(n_369), .Y(n_416) );
BUFx12f_ASAP7_75t_L g417 ( .A(n_369), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_363), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_387), .Y(n_419) );
NAND2x1p5_ASAP7_75t_L g420 ( .A(n_377), .B(n_346), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_367), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_375), .Y(n_422) );
CKINVDCx14_ASAP7_75t_R g423 ( .A(n_365), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_377), .A2(n_313), .B1(n_321), .B2(n_327), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_378), .A2(n_338), .B1(n_331), .B2(n_306), .Y(n_425) );
INVx4_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_370), .Y(n_427) );
CKINVDCx8_ASAP7_75t_R g428 ( .A(n_377), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_370), .Y(n_429) );
INVx3_ASAP7_75t_L g430 ( .A(n_387), .Y(n_430) );
INVx4_ASAP7_75t_L g431 ( .A(n_365), .Y(n_431) );
BUFx12f_ASAP7_75t_L g432 ( .A(n_369), .Y(n_432) );
INVx6_ASAP7_75t_L g433 ( .A(n_369), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_365), .A2(n_375), .B1(n_385), .B2(n_381), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_399), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g436 ( .A1(n_423), .A2(n_375), .B1(n_385), .B2(n_381), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_395), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_410), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_398), .A2(n_378), .B1(n_338), .B2(n_331), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_405), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_401), .A2(n_285), .B1(n_258), .B2(n_288), .Y(n_441) );
OAI21xp5_ASAP7_75t_SL g442 ( .A1(n_401), .A2(n_225), .B(n_306), .Y(n_442) );
AOI211xp5_ASAP7_75t_L g443 ( .A1(n_400), .A2(n_309), .B(n_232), .C(n_272), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_410), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_396), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_430), .B(n_387), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_405), .Y(n_447) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_397), .B(n_232), .C(n_270), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_406), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_404), .B(n_370), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_425), .A2(n_365), .B1(n_388), .B2(n_385), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_413), .A2(n_388), .B1(n_373), .B2(n_369), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_411), .A2(n_376), .B1(n_326), .B2(n_391), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_393), .B(n_391), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_430), .B(n_387), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_411), .A2(n_376), .B1(n_326), .B2(n_391), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_428), .A2(n_376), .B1(n_366), .B2(n_387), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_431), .A2(n_378), .B1(n_338), .B2(n_331), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_412), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_414), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_396), .Y(n_462) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_431), .A2(n_376), .B1(n_342), .B2(n_389), .Y(n_463) );
BUFx4f_ASAP7_75t_L g464 ( .A(n_416), .Y(n_464) );
BUFx12f_ASAP7_75t_L g465 ( .A(n_416), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_431), .A2(n_378), .B1(n_338), .B2(n_331), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_414), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g468 ( .A1(n_417), .A2(n_432), .B1(n_431), .B2(n_410), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_419), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_428), .A2(n_376), .B1(n_366), .B2(n_389), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_410), .A2(n_378), .B1(n_331), .B2(n_338), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_415), .A2(n_389), .B1(n_339), .B2(n_332), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_424), .A2(n_332), .B1(n_371), .B2(n_359), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_421), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_421), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_399), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_417), .A2(n_378), .B1(n_338), .B2(n_331), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_432), .B(n_316), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_427), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_426), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_429), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_402), .Y(n_482) );
BUFx4f_ASAP7_75t_SL g483 ( .A(n_407), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_429), .B(n_343), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_393), .A2(n_378), .B1(n_338), .B2(n_331), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_422), .A2(n_378), .B1(n_331), .B2(n_338), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_422), .A2(n_378), .B1(n_331), .B2(n_338), .Y(n_487) );
CKINVDCx8_ASAP7_75t_R g488 ( .A(n_392), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_434), .A2(n_378), .B1(n_331), .B2(n_330), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_419), .Y(n_490) );
NAND2x1_ASAP7_75t_L g491 ( .A(n_426), .B(n_433), .Y(n_491) );
BUFx4f_ASAP7_75t_SL g492 ( .A(n_426), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_433), .A2(n_336), .B1(n_371), .B2(n_368), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_409), .B(n_368), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_433), .A2(n_336), .B1(n_368), .B2(n_280), .Y(n_495) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_433), .A2(n_368), .B1(n_380), .B2(n_382), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_426), .A2(n_336), .B1(n_280), .B2(n_279), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_440), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g499 ( .A1(n_442), .A2(n_301), .B1(n_317), .B2(n_277), .C(n_322), .Y(n_499) );
AOI221xp5_ASAP7_75t_L g500 ( .A1(n_443), .A2(n_301), .B1(n_317), .B2(n_322), .C(n_232), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_464), .A2(n_420), .B1(n_380), .B2(n_382), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_440), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_464), .A2(n_420), .B1(n_380), .B2(n_382), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_448), .A2(n_301), .B1(n_294), .B2(n_337), .C(n_315), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_492), .A2(n_420), .B1(n_352), .B2(n_382), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_438), .A2(n_382), .B1(n_380), .B2(n_328), .Y(n_506) );
NAND3xp33_ASAP7_75t_SL g507 ( .A(n_437), .B(n_318), .C(n_237), .Y(n_507) );
OA222x2_ASAP7_75t_L g508 ( .A1(n_454), .A2(n_409), .B1(n_347), .B2(n_390), .C1(n_379), .C2(n_346), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_438), .A2(n_382), .B1(n_361), .B2(n_386), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_439), .A2(n_347), .B1(n_280), .B2(n_279), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g511 ( .A1(n_444), .A2(n_374), .B1(n_347), .B2(n_382), .Y(n_511) );
OAI222xp33_ASAP7_75t_L g512 ( .A1(n_444), .A2(n_347), .B1(n_374), .B2(n_379), .C1(n_390), .C2(n_357), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_451), .A2(n_347), .B1(n_279), .B2(n_346), .Y(n_513) );
OAI221xp5_ASAP7_75t_SL g514 ( .A1(n_441), .A2(n_337), .B1(n_344), .B2(n_315), .C(n_319), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_447), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_450), .B(n_337), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_452), .A2(n_279), .B1(n_346), .B2(n_320), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_457), .A2(n_456), .B1(n_453), .B2(n_489), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_447), .B(n_392), .Y(n_519) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_483), .A2(n_361), .B1(n_386), .B2(n_394), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_472), .A2(n_320), .B1(n_271), .B2(n_357), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_464), .A2(n_374), .B1(n_390), .B2(n_379), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_473), .A2(n_320), .B1(n_271), .B2(n_351), .Y(n_523) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_480), .A2(n_386), .B1(n_361), .B2(n_394), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_436), .A2(n_320), .B1(n_271), .B2(n_351), .Y(n_525) );
NAND3xp33_ASAP7_75t_SL g526 ( .A(n_437), .B(n_374), .C(n_292), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_497), .A2(n_271), .B1(n_379), .B2(n_390), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_468), .A2(n_374), .B1(n_379), .B2(n_390), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_470), .A2(n_271), .B1(n_361), .B2(n_386), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_480), .A2(n_386), .B1(n_403), .B2(n_394), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_495), .A2(n_271), .B1(n_386), .B2(n_350), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_445), .B(n_19), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_493), .A2(n_271), .B1(n_386), .B2(n_350), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_471), .A2(n_271), .B1(n_386), .B2(n_350), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_485), .A2(n_255), .B1(n_403), .B2(n_394), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_435), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_465), .A2(n_408), .B1(n_403), .B2(n_394), .Y(n_537) );
AO22x1_ASAP7_75t_L g538 ( .A1(n_445), .A2(n_408), .B1(n_403), .B2(n_392), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_486), .A2(n_408), .B1(n_403), .B2(n_392), .Y(n_539) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_465), .A2(n_408), .B1(n_392), .B2(n_335), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_477), .A2(n_355), .B1(n_333), .B2(n_408), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_487), .A2(n_355), .B1(n_354), .B2(n_345), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_458), .A2(n_355), .B1(n_354), .B2(n_345), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g544 ( .A1(n_478), .A2(n_261), .B1(n_260), .B2(n_300), .C(n_308), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_466), .A2(n_335), .B1(n_297), .B2(n_296), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_446), .A2(n_289), .B1(n_287), .B2(n_325), .Y(n_546) );
OAI222xp33_ASAP7_75t_L g547 ( .A1(n_461), .A2(n_239), .B1(n_236), .B2(n_296), .C1(n_297), .C2(n_287), .Y(n_547) );
OAI21xp33_ASAP7_75t_L g548 ( .A1(n_462), .A2(n_150), .B(n_147), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_462), .A2(n_345), .B1(n_354), .B2(n_324), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_446), .A2(n_325), .B1(n_289), .B2(n_287), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_455), .A2(n_289), .B1(n_325), .B2(n_323), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_459), .B(n_307), .Y(n_552) );
OAI22xp33_ASAP7_75t_L g553 ( .A1(n_467), .A2(n_345), .B1(n_354), .B2(n_324), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_469), .A2(n_323), .B1(n_298), .B2(n_324), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_490), .A2(n_323), .B1(n_324), .B2(n_265), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_474), .B(n_307), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_474), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_490), .A2(n_265), .B1(n_354), .B2(n_281), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_449), .B(n_19), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_475), .B(n_479), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_496), .A2(n_310), .B1(n_302), .B2(n_275), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_463), .A2(n_281), .B1(n_283), .B2(n_262), .Y(n_562) );
OAI211xp5_ASAP7_75t_SL g563 ( .A1(n_460), .A2(n_262), .B(n_250), .C(n_283), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_454), .A2(n_275), .B1(n_310), .B2(n_302), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_491), .A2(n_310), .B1(n_302), .B2(n_303), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_479), .A2(n_282), .B1(n_307), .B2(n_235), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_481), .A2(n_282), .B1(n_307), .B2(n_299), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_481), .A2(n_282), .B1(n_299), .B2(n_290), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_484), .A2(n_282), .B1(n_299), .B2(n_290), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_494), .A2(n_314), .B1(n_299), .B2(n_290), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_476), .B(n_147), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_476), .A2(n_211), .B1(n_210), .B2(n_222), .Y(n_572) );
BUFx8_ASAP7_75t_SL g573 ( .A(n_482), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_488), .B(n_20), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_488), .A2(n_314), .B1(n_299), .B2(n_290), .Y(n_575) );
NAND3xp33_ASAP7_75t_L g576 ( .A(n_442), .B(n_147), .C(n_150), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_442), .B(n_21), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_577), .A2(n_576), .B1(n_559), .B2(n_499), .C(n_500), .Y(n_578) );
AOI21xp5_ASAP7_75t_SL g579 ( .A1(n_526), .A2(n_240), .B(n_22), .Y(n_579) );
NAND3xp33_ASAP7_75t_SL g580 ( .A(n_532), .B(n_21), .C(n_22), .Y(n_580) );
OAI221xp5_ASAP7_75t_SL g581 ( .A1(n_518), .A2(n_23), .B1(n_24), .B2(n_25), .C(n_26), .Y(n_581) );
NOR3xp33_ASAP7_75t_L g582 ( .A(n_574), .B(n_218), .C(n_219), .Y(n_582) );
NAND4xp25_ASAP7_75t_L g583 ( .A(n_514), .B(n_268), .C(n_25), .D(n_26), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_511), .A2(n_158), .B1(n_150), .B2(n_314), .Y(n_584) );
OA211x2_ASAP7_75t_L g585 ( .A1(n_548), .A2(n_24), .B(n_27), .C(n_28), .Y(n_585) );
AND2x2_ASAP7_75t_SL g586 ( .A(n_508), .B(n_314), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_508), .B(n_150), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_519), .B(n_158), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_504), .A2(n_158), .B1(n_314), .B2(n_230), .Y(n_589) );
NOR3xp33_ASAP7_75t_SL g590 ( .A(n_507), .B(n_30), .C(n_31), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_515), .B(n_30), .Y(n_591) );
AOI21xp5_ASAP7_75t_SL g592 ( .A1(n_528), .A2(n_32), .B(n_34), .Y(n_592) );
NAND2xp33_ASAP7_75t_SL g593 ( .A(n_511), .B(n_34), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_560), .B(n_37), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_557), .B(n_38), .Y(n_595) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_506), .A2(n_158), .B(n_38), .Y(n_596) );
NOR3xp33_ASAP7_75t_L g597 ( .A(n_544), .B(n_223), .C(n_230), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_552), .B(n_42), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_516), .B(n_224), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_556), .B(n_43), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_556), .B(n_44), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_573), .B(n_45), .Y(n_602) );
AND2x2_ASAP7_75t_SL g603 ( .A(n_573), .B(n_216), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_529), .B(n_220), .C(n_243), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_513), .A2(n_243), .B1(n_256), .B2(n_228), .C(n_46), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_563), .B(n_256), .C(n_228), .Y(n_606) );
OAI21xp5_ASAP7_75t_SL g607 ( .A1(n_512), .A2(n_216), .B(n_50), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_536), .B(n_52), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_564), .B(n_54), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_571), .B(n_61), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_509), .B(n_228), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_540), .A2(n_62), .B(n_63), .Y(n_612) );
OAI21xp5_ASAP7_75t_SL g613 ( .A1(n_520), .A2(n_64), .B(n_67), .Y(n_613) );
OA21x2_ASAP7_75t_L g614 ( .A1(n_539), .A2(n_70), .B(n_71), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_524), .B(n_72), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_530), .B(n_73), .Y(n_616) );
AOI21xp5_ASAP7_75t_SL g617 ( .A1(n_501), .A2(n_77), .B(n_78), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_537), .B(n_81), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_522), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_503), .A2(n_86), .B1(n_89), .B2(n_90), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_553), .B(n_91), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_517), .B(n_93), .Y(n_622) );
NOR2xp33_ASAP7_75t_SL g623 ( .A(n_547), .B(n_92), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_562), .B(n_527), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_546), .B(n_550), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_565), .B(n_543), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_566), .B(n_567), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_533), .B(n_534), .C(n_535), .Y(n_628) );
OAI21xp5_ASAP7_75t_SL g629 ( .A1(n_549), .A2(n_542), .B(n_525), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_541), .B(n_561), .Y(n_630) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_531), .A2(n_558), .B(n_545), .Y(n_631) );
NAND3xp33_ASAP7_75t_L g632 ( .A(n_521), .B(n_523), .C(n_572), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_538), .B(n_510), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_551), .A2(n_569), .B1(n_555), .B2(n_554), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_538), .B(n_570), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_575), .B(n_568), .Y(n_636) );
OAI221xp5_ASAP7_75t_L g637 ( .A1(n_577), .A2(n_442), .B1(n_401), .B2(n_576), .C(n_443), .Y(n_637) );
NAND2xp33_ASAP7_75t_SL g638 ( .A(n_511), .B(n_438), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g639 ( .A(n_576), .B(n_442), .C(n_577), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_576), .B(n_442), .C(n_577), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_500), .A2(n_576), .B1(n_448), .B2(n_499), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_577), .B(n_576), .C(n_442), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_508), .B(n_449), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_498), .B(n_502), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_508), .B(n_449), .Y(n_645) );
OAI221xp5_ASAP7_75t_SL g646 ( .A1(n_499), .A2(n_442), .B1(n_576), .B2(n_443), .C(n_500), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_500), .A2(n_576), .B1(n_448), .B2(n_499), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_505), .A2(n_576), .B1(n_464), .B2(n_468), .Y(n_648) );
NAND4xp75_ASAP7_75t_L g649 ( .A(n_603), .B(n_587), .C(n_586), .D(n_621), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_596), .A2(n_607), .B(n_592), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_643), .B(n_645), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_639), .B(n_640), .C(n_642), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_619), .B(n_586), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_637), .B(n_646), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_638), .B(n_593), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_644), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_638), .A2(n_593), .B1(n_578), .B2(n_648), .Y(n_657) );
NAND4xp75_ASAP7_75t_L g658 ( .A(n_603), .B(n_633), .C(n_626), .D(n_590), .Y(n_658) );
NAND3xp33_ASAP7_75t_L g659 ( .A(n_629), .B(n_647), .C(n_641), .Y(n_659) );
NOR3xp33_ASAP7_75t_L g660 ( .A(n_580), .B(n_583), .C(n_581), .Y(n_660) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_641), .A2(n_647), .B(n_579), .C(n_613), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_635), .B(n_588), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_598), .B(n_627), .Y(n_663) );
AOI211xp5_ASAP7_75t_L g664 ( .A1(n_617), .A2(n_626), .B(n_623), .C(n_621), .Y(n_664) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_591), .A2(n_595), .B1(n_632), .B2(n_614), .Y(n_665) );
NAND4xp75_ASAP7_75t_L g666 ( .A(n_585), .B(n_602), .C(n_611), .D(n_614), .Y(n_666) );
INVx1_ASAP7_75t_SL g667 ( .A(n_594), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_608), .B(n_630), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_624), .B(n_600), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_584), .B(n_628), .C(n_582), .Y(n_670) );
BUFx3_ASAP7_75t_L g671 ( .A(n_618), .Y(n_671) );
NAND4xp75_ASAP7_75t_L g672 ( .A(n_636), .B(n_616), .C(n_615), .D(n_631), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_601), .B(n_634), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_599), .B(n_589), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_589), .B(n_597), .Y(n_675) );
NAND4xp75_ASAP7_75t_L g676 ( .A(n_625), .B(n_622), .C(n_609), .D(n_610), .Y(n_676) );
AO21x2_ASAP7_75t_L g677 ( .A1(n_612), .A2(n_604), .B(n_605), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_620), .B(n_606), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_586), .B(n_587), .Y(n_679) );
OR2x2_ASAP7_75t_L g680 ( .A(n_619), .B(n_643), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_643), .B(n_645), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_643), .B(n_645), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_643), .B(n_645), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_587), .A2(n_648), .B(n_638), .C(n_607), .Y(n_684) );
NOR3xp33_ASAP7_75t_SL g685 ( .A(n_637), .B(n_646), .C(n_638), .Y(n_685) );
OAI22xp33_ASAP7_75t_L g686 ( .A1(n_607), .A2(n_648), .B1(n_587), .B2(n_623), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_643), .B(n_645), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_643), .B(n_645), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_587), .B(n_640), .C(n_639), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_643), .B(n_645), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_587), .B(n_640), .C(n_639), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_643), .B(n_645), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_643), .B(n_645), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_619), .B(n_643), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_643), .B(n_645), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_643), .B(n_645), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g697 ( .A(n_580), .B(n_646), .C(n_583), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_637), .B(n_437), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_643), .B(n_645), .Y(n_699) );
NOR2x1_ASAP7_75t_L g700 ( .A(n_648), .B(n_607), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_643), .B(n_645), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_643), .B(n_645), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_619), .B(n_643), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_662), .Y(n_704) );
INVx3_ASAP7_75t_L g705 ( .A(n_653), .Y(n_705) );
XNOR2xp5_ASAP7_75t_L g706 ( .A(n_685), .B(n_657), .Y(n_706) );
NOR4xp25_ASAP7_75t_L g707 ( .A(n_659), .B(n_652), .C(n_687), .D(n_701), .Y(n_707) );
INVx2_ASAP7_75t_SL g708 ( .A(n_679), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_656), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_681), .B(n_683), .Y(n_710) );
NAND4xp75_ASAP7_75t_L g711 ( .A(n_700), .B(n_655), .C(n_650), .D(n_679), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_680), .B(n_703), .Y(n_712) );
NAND4xp75_ASAP7_75t_L g713 ( .A(n_655), .B(n_654), .C(n_678), .D(n_698), .Y(n_713) );
NOR2x1p5_ASAP7_75t_L g714 ( .A(n_649), .B(n_658), .Y(n_714) );
AND4x1_ASAP7_75t_L g715 ( .A(n_684), .B(n_664), .C(n_691), .D(n_689), .Y(n_715) );
NAND4xp75_ASAP7_75t_SL g716 ( .A(n_678), .B(n_661), .C(n_686), .D(n_690), .Y(n_716) );
INVx1_ASAP7_75t_SL g717 ( .A(n_667), .Y(n_717) );
OR2x2_ASAP7_75t_L g718 ( .A(n_703), .B(n_694), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_680), .Y(n_719) );
NOR4xp25_ASAP7_75t_L g720 ( .A(n_651), .B(n_688), .C(n_699), .D(n_696), .Y(n_720) );
NAND4xp25_ASAP7_75t_SL g721 ( .A(n_682), .B(n_693), .C(n_665), .D(n_702), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_692), .B(n_695), .Y(n_722) );
INVx4_ASAP7_75t_L g723 ( .A(n_677), .Y(n_723) );
NAND4xp75_ASAP7_75t_L g724 ( .A(n_673), .B(n_675), .C(n_674), .D(n_663), .Y(n_724) );
INVx1_ASAP7_75t_SL g725 ( .A(n_671), .Y(n_725) );
XNOR2x2_ASAP7_75t_L g726 ( .A(n_649), .B(n_672), .Y(n_726) );
XNOR2xp5_ASAP7_75t_L g727 ( .A(n_706), .B(n_697), .Y(n_727) );
XNOR2xp5_ASAP7_75t_L g728 ( .A(n_706), .B(n_669), .Y(n_728) );
INVxp33_ASAP7_75t_SL g729 ( .A(n_711), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_713), .B(n_670), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_720), .B(n_668), .Y(n_731) );
INVxp67_ASAP7_75t_L g732 ( .A(n_713), .Y(n_732) );
XNOR2x2_ASAP7_75t_L g733 ( .A(n_726), .B(n_666), .Y(n_733) );
XOR2x2_ASAP7_75t_L g734 ( .A(n_716), .B(n_660), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_704), .Y(n_735) );
INVx1_ASAP7_75t_SL g736 ( .A(n_717), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_709), .Y(n_737) );
XNOR2x1_ASAP7_75t_L g738 ( .A(n_726), .B(n_676), .Y(n_738) );
INVx1_ASAP7_75t_SL g739 ( .A(n_725), .Y(n_739) );
XOR2x2_ASAP7_75t_L g740 ( .A(n_715), .B(n_671), .Y(n_740) );
INVx4_ASAP7_75t_L g741 ( .A(n_740), .Y(n_741) );
INVxp67_ASAP7_75t_SL g742 ( .A(n_733), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_729), .A2(n_714), .B1(n_721), .B2(n_724), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_730), .A2(n_724), .B1(n_707), .B2(n_708), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_735), .Y(n_745) );
INVx3_ASAP7_75t_SL g746 ( .A(n_736), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_737), .B(n_719), .Y(n_747) );
OA22x2_ASAP7_75t_L g748 ( .A1(n_732), .A2(n_723), .B1(n_710), .B2(n_722), .Y(n_748) );
OAI22xp33_ASAP7_75t_L g749 ( .A1(n_731), .A2(n_705), .B1(n_712), .B2(n_718), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_745), .Y(n_750) );
OA22x2_ASAP7_75t_L g751 ( .A1(n_741), .A2(n_727), .B1(n_728), .B2(n_733), .Y(n_751) );
INVx2_ASAP7_75t_SL g752 ( .A(n_746), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_742), .Y(n_753) );
INVx1_ASAP7_75t_SL g754 ( .A(n_741), .Y(n_754) );
INVxp67_ASAP7_75t_SL g755 ( .A(n_742), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_744), .Y(n_756) );
INVxp67_ASAP7_75t_SL g757 ( .A(n_748), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_747), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_756), .A2(n_734), .B1(n_751), .B2(n_743), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_752), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_755), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_753), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_756), .A2(n_734), .B1(n_738), .B2(n_740), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_760), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_763), .A2(n_751), .B1(n_754), .B2(n_738), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_759), .B(n_727), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_764), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_766), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_765), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g770 ( .A(n_769), .B(n_752), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_767), .Y(n_771) );
OAI31xp33_ASAP7_75t_L g772 ( .A1(n_770), .A2(n_761), .A3(n_768), .B(n_762), .Y(n_772) );
AND2x4_ASAP7_75t_L g773 ( .A(n_771), .B(n_767), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_773), .Y(n_774) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_773), .Y(n_775) );
INVxp67_ASAP7_75t_SL g776 ( .A(n_775), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_776), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_777), .A2(n_774), .B1(n_775), .B2(n_750), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_778), .Y(n_779) );
OAI22xp33_ASAP7_75t_L g780 ( .A1(n_779), .A2(n_775), .B1(n_757), .B2(n_772), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_780), .Y(n_781) );
AOI221xp5_ASAP7_75t_L g782 ( .A1(n_781), .A2(n_775), .B1(n_749), .B2(n_758), .C(n_728), .Y(n_782) );
AOI211xp5_ASAP7_75t_L g783 ( .A1(n_782), .A2(n_775), .B(n_749), .C(n_739), .Y(n_783) );
endmodule