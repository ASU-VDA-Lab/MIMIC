module fake_jpeg_563_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_54),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_0),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_58),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_0),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_55),
.A2(n_44),
.B1(n_42),
.B2(n_45),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_65),
.B1(n_69),
.B2(n_40),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_44),
.B1(n_52),
.B2(n_47),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_47),
.B1(n_43),
.B2(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_49),
.B1(n_48),
.B2(n_3),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_73),
.Y(n_88)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_46),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_46),
.B1(n_40),
.B2(n_3),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_1),
.B(n_2),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_9),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_61),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_40),
.C(n_15),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_82),
.B1(n_68),
.B2(n_62),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_68),
.B(n_6),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_5),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_75),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_96),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_94),
.B1(n_76),
.B2(n_12),
.Y(n_110)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_94),
.Y(n_100)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_80),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_106),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_11),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_110),
.A2(n_105),
.B(n_108),
.Y(n_112)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_113),
.C(n_121),
.Y(n_124)
);

NOR4xp25_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_27),
.C(n_13),
.D(n_14),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_96),
.B(n_91),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_97),
.C(n_102),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_12),
.A3(n_16),
.B1(n_17),
.B2(n_19),
.C1(n_21),
.C2(n_22),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_99),
.B1(n_110),
.B2(n_32),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_125),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_99),
.C(n_30),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_124),
.B(n_114),
.Y(n_126)
);

NAND4xp25_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_116),
.C(n_118),
.D(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_128),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_127),
.C(n_121),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_34),
.C(n_29),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_133),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_33),
.Y(n_135)
);


endmodule