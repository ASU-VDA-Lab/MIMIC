module fake_jpeg_27719_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_55),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_20),
.B1(n_25),
.B2(n_32),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_60),
.B1(n_25),
.B2(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_21),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_28),
.B1(n_32),
.B2(n_19),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_41),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_25),
.B1(n_27),
.B2(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_34),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_63),
.A2(n_65),
.B(n_73),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_19),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_77),
.Y(n_104)
);

NAND2x1p5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_28),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_36),
.B1(n_43),
.B2(n_42),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_91),
.B1(n_50),
.B2(n_57),
.Y(n_100)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_46),
.B(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_16),
.B1(n_33),
.B2(n_18),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_18),
.B1(n_33),
.B2(n_16),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_57),
.B1(n_53),
.B2(n_18),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_47),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_86),
.Y(n_114)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_34),
.C(n_41),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_31),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_18),
.B1(n_33),
.B2(n_22),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_95),
.A2(n_78),
.B(n_90),
.C(n_39),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_106),
.Y(n_130)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_68),
.B(n_34),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_111),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_34),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_116),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_41),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_117),
.A2(n_87),
.B1(n_92),
.B2(n_71),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_74),
.A2(n_57),
.B1(n_39),
.B2(n_26),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_72),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_110),
.B(n_64),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_122),
.B(n_135),
.Y(n_157)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_68),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_143),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_128),
.A2(n_133),
.B(n_146),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_129),
.B(n_134),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_64),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_98),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_145),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_75),
.Y(n_139)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_86),
.Y(n_140)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_141),
.B(n_142),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_63),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_147),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

AOI22x1_ASAP7_75t_SL g146 ( 
.A1(n_97),
.A2(n_74),
.B1(n_63),
.B2(n_88),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_115),
.B1(n_99),
.B2(n_83),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_97),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

OR2x6_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_97),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_152),
.A2(n_154),
.B(n_158),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_121),
.B(n_102),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_132),
.A2(n_94),
.B1(n_102),
.B2(n_111),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_132),
.A2(n_94),
.B1(n_119),
.B2(n_105),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_9),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_103),
.C(n_39),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_173),
.C(n_180),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_8),
.C(n_15),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_163),
.B(n_11),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_125),
.B(n_134),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_164),
.B(n_17),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_31),
.A3(n_29),
.B1(n_22),
.B2(n_93),
.C1(n_117),
.C2(n_26),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_183),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_113),
.B1(n_103),
.B2(n_99),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_145),
.B1(n_136),
.B2(n_123),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_137),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_168),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_58),
.C(n_85),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_124),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_174),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_98),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_178),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_128),
.B1(n_136),
.B2(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_26),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_115),
.C(n_17),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_31),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_184),
.Y(n_201)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_22),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_205),
.B1(n_158),
.B2(n_156),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_186),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_192),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_154),
.A2(n_149),
.B1(n_123),
.B2(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_149),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_195),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_152),
.A2(n_29),
.A3(n_17),
.B1(n_7),
.B2(n_12),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_203),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_152),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_199)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_6),
.C(n_14),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_206),
.C(n_159),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_152),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_204)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_152),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_6),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_164),
.A2(n_179),
.B1(n_176),
.B2(n_180),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_0),
.Y(n_210)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_160),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_160),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_SL g240 ( 
.A1(n_214),
.A2(n_178),
.B(n_182),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_171),
.B(n_153),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_215),
.Y(n_228)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_230),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_220),
.A2(n_199),
.B1(n_204),
.B2(n_214),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_155),
.B1(n_181),
.B2(n_184),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_155),
.B1(n_197),
.B2(n_185),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_151),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_206),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_190),
.Y(n_230)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_194),
.C(n_191),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_251),
.C(n_256),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_257),
.Y(n_264)
);

XOR2x2_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_193),
.Y(n_245)
);

OAI31xp33_ASAP7_75t_L g277 ( 
.A1(n_245),
.A2(n_237),
.A3(n_238),
.B(n_196),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_225),
.B1(n_221),
.B2(n_227),
.Y(n_272)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_194),
.C(n_193),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_201),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_173),
.C(n_195),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_229),
.B(n_202),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_151),
.C(n_189),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_260),
.C(n_236),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_225),
.B1(n_222),
.B2(n_227),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_183),
.C(n_172),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_231),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_270),
.Y(n_283)
);

FAx1_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_221),
.CI(n_222),
.CON(n_263),
.SN(n_263)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_263),
.B(n_277),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_266),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_244),
.B1(n_242),
.B2(n_250),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_258),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_257),
.C(n_256),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_254),
.C(n_228),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_273),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_238),
.B1(n_237),
.B2(n_214),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_279),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_219),
.B1(n_216),
.B2(n_232),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_243),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_263),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_259),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_289),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_290),
.C(n_271),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

INVx11_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_177),
.C(n_165),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_212),
.B1(n_211),
.B2(n_156),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_261),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_293),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_276),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_263),
.B(n_275),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_294),
.A2(n_6),
.B(n_12),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_299),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_210),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_302),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_264),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_303),
.B(n_9),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_296),
.B1(n_293),
.B2(n_297),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_13),
.B1(n_15),
.B2(n_5),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g306 ( 
.A(n_295),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_309),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_290),
.B1(n_284),
.B2(n_279),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_281),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_311),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_304),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_296),
.B1(n_303),
.B2(n_298),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_316),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_13),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_320),
.B(n_315),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_307),
.B(n_15),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_318),
.C(n_314),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_307),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_313),
.B(n_3),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_4),
.C(n_323),
.Y(n_326)
);


endmodule