module fake_jpeg_24786_n_99 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_99);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_99;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_3),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_22),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_27),
.Y(n_29)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_26),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_9),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_14),
.B(n_18),
.Y(n_33)
);

AND2x6_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_35),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_10),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_13),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_27),
.B1(n_24),
.B2(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_15),
.B1(n_26),
.B2(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_31),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

FAx1_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_30),
.CI(n_25),
.CON(n_52),
.SN(n_52)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_60),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_38),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_49),
.B(n_40),
.C(n_43),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_59),
.B(n_54),
.C(n_38),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_42),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_69),
.C(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_61),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_39),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_58),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_54),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_31),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_64),
.Y(n_80)
);

BUFx24_ASAP7_75t_SL g83 ( 
.A(n_80),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_31),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_71),
.C(n_76),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_17),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_74),
.B(n_76),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_87),
.Y(n_89)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_88),
.Y(n_91)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_17),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_6),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_93),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_89),
.B(n_83),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_93),
.B1(n_1),
.B2(n_2),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_0),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_0),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_95),
.Y(n_99)
);


endmodule