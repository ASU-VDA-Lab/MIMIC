module fake_jpeg_21273_n_39 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_39);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx3_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_6),
.B1(n_12),
.B2(n_9),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_17),
.B1(n_21),
.B2(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_26),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_1),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_34),
.B(n_30),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_33),
.B1(n_32),
.B2(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

OAI222xp33_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_7),
.B1(n_8),
.B2(n_4),
.C1(n_22),
.C2(n_18),
.Y(n_38)
);

AOI322xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_19),
.C1(n_22),
.C2(n_23),
.Y(n_39)
);


endmodule