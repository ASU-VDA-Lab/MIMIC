module fake_jpeg_3414_n_178 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_46),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_56),
.B1(n_47),
.B2(n_52),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_72),
.B1(n_69),
.B2(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_61),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_84),
.Y(n_98)
);

FAx1_ASAP7_75t_SL g84 ( 
.A(n_80),
.B(n_57),
.CI(n_50),
.CON(n_84),
.SN(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_47),
.B1(n_56),
.B2(n_50),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_85),
.A2(n_90),
.B1(n_20),
.B2(n_34),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_54),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_89),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_54),
.B1(n_57),
.B2(n_2),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_92),
.B1(n_4),
.B2(n_5),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_0),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_95),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_1),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_19),
.A3(n_41),
.B1(n_38),
.B2(n_35),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_28),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_17),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_116),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_18),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_3),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_115),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_114),
.B1(n_8),
.B2(n_10),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_4),
.B(n_5),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_6),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_6),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_23),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_114),
.A2(n_85),
.B1(n_96),
.B2(n_9),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_126),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_105),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_133),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_129),
.B(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_11),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_132),
.B1(n_116),
.B2(n_15),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_27),
.B1(n_33),
.B2(n_32),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_13),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_126),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_137),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_112),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_138),
.B(n_44),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_109),
.B(n_112),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_151),
.B(n_29),
.C(n_30),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_99),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_149),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_144),
.B1(n_131),
.B2(n_121),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_15),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_128),
.B(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_147),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_125),
.B1(n_121),
.B2(n_127),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_155),
.B1(n_151),
.B2(n_150),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_16),
.B1(n_24),
.B2(n_25),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_144),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_139),
.C(n_146),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_162),
.B(n_163),
.Y(n_168)
);

OA21x2_ASAP7_75t_SL g162 ( 
.A1(n_153),
.A2(n_140),
.B(n_160),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_166),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_156),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_157),
.C(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_168),
.A2(n_166),
.B1(n_138),
.B2(n_159),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_164),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_170),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_169),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g176 ( 
.A(n_175),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_157),
.C(n_145),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_145),
.Y(n_178)
);


endmodule