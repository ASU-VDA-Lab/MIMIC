module fake_jpeg_11197_n_190 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_190);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_10),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_17),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_88),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_0),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_72),
.B1(n_78),
.B2(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_65),
.B1(n_64),
.B2(n_68),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_60),
.B1(n_77),
.B2(n_78),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_76),
.B1(n_80),
.B2(n_79),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_113),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_111),
.Y(n_135)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_66),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_117),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_81),
.B1(n_60),
.B2(n_77),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_127),
.B1(n_6),
.B2(n_8),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_53),
.B1(n_68),
.B2(n_64),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_129),
.B1(n_2),
.B2(n_4),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_69),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_124),
.B1(n_89),
.B2(n_1),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_126),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_84),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_122),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_54),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_89),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_56),
.B1(n_71),
.B2(n_57),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_55),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_5),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_73),
.B1(n_63),
.B2(n_59),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_147),
.Y(n_155)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_145),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_21),
.B(n_48),
.C(n_46),
.D(n_45),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_140),
.B(n_28),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_0),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_137),
.B(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_151),
.B1(n_9),
.B2(n_10),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_5),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_6),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_152),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_29),
.C(n_39),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_165),
.C(n_167),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_160),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_8),
.B(n_9),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_149),
.B(n_138),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_30),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_11),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_31),
.C(n_37),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_135),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_155),
.C(n_162),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_154),
.A2(n_144),
.B1(n_134),
.B2(n_140),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_172),
.C(n_173),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_166),
.A2(n_141),
.B(n_139),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_153),
.A2(n_16),
.B(n_35),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_177),
.A2(n_180),
.B1(n_159),
.B2(n_168),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_156),
.B(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_182),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_179),
.C(n_174),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_184),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_175),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_153),
.B1(n_161),
.B2(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_51),
.B(n_13),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_15),
.Y(n_190)
);


endmodule