module fake_jpeg_14382_n_580 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_580);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_580;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_55),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_80),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_96),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx2_ASAP7_75t_R g173 ( 
.A(n_63),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_26),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_65),
.B(n_72),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_69),
.Y(n_172)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_70),
.Y(n_161)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_16),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_75),
.Y(n_167)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_79),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_40),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_99),
.Y(n_110)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_53),
.B(n_16),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_101),
.B(n_103),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_104),
.Y(n_166)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_108),
.Y(n_111)
);

BUFx6f_ASAP7_75t_SL g106 ( 
.A(n_42),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_SL g154 ( 
.A(n_106),
.Y(n_154)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_45),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_53),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_50),
.B(n_38),
.C(n_48),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_139),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_62),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_119),
.B(n_120),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_50),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_41),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_126),
.B(n_128),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_41),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_62),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_130),
.B(n_136),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_55),
.Y(n_136)
);

OR2x2_ASAP7_75t_SL g137 ( 
.A(n_63),
.B(n_33),
.Y(n_137)
);

OR2x2_ASAP7_75t_SL g228 ( 
.A(n_137),
.B(n_139),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_85),
.A2(n_51),
.B(n_48),
.C(n_46),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_77),
.A2(n_81),
.B1(n_66),
.B2(n_60),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_157),
.B1(n_170),
.B2(n_87),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_143),
.B(n_45),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_102),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_153),
.B(n_159),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_93),
.A2(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_97),
.B(n_41),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_97),
.B(n_41),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_163),
.B(n_171),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_107),
.A2(n_28),
.B1(n_46),
.B2(n_24),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_170),
.A2(n_23),
.B1(n_28),
.B2(n_45),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_54),
.B(n_41),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_33),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_174),
.B(n_184),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_175),
.A2(n_204),
.B1(n_213),
.B2(n_167),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_176),
.Y(n_283)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g255 ( 
.A(n_177),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_178),
.Y(n_276)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_137),
.A2(n_32),
.B1(n_36),
.B2(n_38),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_180),
.A2(n_209),
.B1(n_222),
.B2(n_227),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_36),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_188),
.Y(n_261)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_189),
.Y(n_271)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_156),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_191),
.B(n_193),
.Y(n_258)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_192),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_145),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_125),
.A2(n_67),
.B1(n_64),
.B2(n_73),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_194),
.A2(n_195),
.B1(n_151),
.B2(n_142),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_125),
.A2(n_75),
.B1(n_91),
.B2(n_90),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_196),
.Y(n_274)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_199),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_115),
.B(n_103),
.C(n_89),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_200),
.B(n_135),
.C(n_132),
.Y(n_253)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_201),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_134),
.B(n_32),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_203),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_121),
.B(n_51),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_118),
.A2(n_28),
.B1(n_22),
.B2(n_23),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_205),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_131),
.Y(n_206)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_206),
.Y(n_275)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_207),
.Y(n_288)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_208),
.B(n_212),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_161),
.A2(n_69),
.B1(n_43),
.B2(n_29),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_217),
.Y(n_238)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_114),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_111),
.B(n_12),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_215),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_133),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_220),
.Y(n_272)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_219),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_113),
.B(n_13),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_221),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_45),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_223),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_122),
.B(n_45),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_224),
.Y(n_290)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_129),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_225),
.Y(n_291)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_129),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_229),
.Y(n_240)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_158),
.A2(n_43),
.B1(n_29),
.B2(n_21),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_236),
.B1(n_114),
.B2(n_162),
.Y(n_250)
);

INVx6_ASAP7_75t_SL g231 ( 
.A(n_160),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_233),
.Y(n_243)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_158),
.A2(n_144),
.B1(n_138),
.B2(n_142),
.Y(n_232)
);

AO22x1_ASAP7_75t_SL g266 ( 
.A1(n_232),
.A2(n_166),
.B1(n_58),
.B2(n_54),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_122),
.B(n_43),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_138),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_235),
.Y(n_264)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_169),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_186),
.A2(n_147),
.B1(n_144),
.B2(n_169),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_237),
.A2(n_248),
.B1(n_251),
.B2(n_286),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_245),
.A2(n_250),
.B1(n_262),
.B2(n_263),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_186),
.A2(n_167),
.B1(n_141),
.B2(n_152),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_218),
.A2(n_141),
.B1(n_152),
.B2(n_149),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_253),
.B(n_265),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_207),
.C(n_208),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_259),
.B(n_260),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_147),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_213),
.A2(n_149),
.B1(n_117),
.B2(n_127),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_211),
.A2(n_162),
.B1(n_117),
.B2(n_127),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_217),
.B(n_146),
.Y(n_265)
);

AO21x2_ASAP7_75t_L g334 ( 
.A1(n_266),
.A2(n_6),
.B(n_8),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_232),
.A2(n_29),
.B1(n_21),
.B2(n_146),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_278),
.A2(n_292),
.B1(n_4),
.B2(n_5),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_200),
.B(n_58),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_282),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_190),
.B(n_1),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_199),
.B(n_1),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_287),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_229),
.B(n_2),
.C(n_3),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_181),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_232),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_181),
.B(n_2),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_232),
.A2(n_225),
.B1(n_227),
.B2(n_197),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_293),
.B(n_297),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_244),
.A2(n_188),
.B1(n_235),
.B2(n_210),
.Y(n_294)
);

OAI22x1_ASAP7_75t_L g375 ( 
.A1(n_294),
.A2(n_307),
.B1(n_312),
.B2(n_325),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_182),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_295),
.Y(n_366)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_296),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_198),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_245),
.A2(n_234),
.B1(n_189),
.B2(n_179),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_298),
.A2(n_311),
.B1(n_326),
.B2(n_333),
.Y(n_365)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_299),
.Y(n_385)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_244),
.Y(n_300)
);

INVx8_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_276),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_302),
.B(n_314),
.Y(n_350)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_261),
.A2(n_188),
.B1(n_231),
.B2(n_192),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_268),
.B(n_201),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_308),
.B(n_320),
.Y(n_369)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_261),
.Y(n_309)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_309),
.Y(n_378)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_310),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_292),
.A2(n_222),
.B1(n_206),
.B2(n_187),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_286),
.A2(n_236),
.B1(n_212),
.B2(n_220),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_264),
.Y(n_313)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_313),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_280),
.Y(n_314)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

INVx4_ASAP7_75t_SL g316 ( 
.A(n_266),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_316),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_240),
.B(n_196),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_317),
.B(n_318),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_240),
.B(n_183),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_288),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_319),
.B(n_324),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_259),
.B(n_176),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_267),
.B(n_215),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_248),
.A2(n_177),
.B1(n_205),
.B2(n_219),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_281),
.B(n_4),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_327),
.B(n_328),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_272),
.B(n_284),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_238),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_336),
.Y(n_352)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_260),
.B(n_11),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_SL g357 ( 
.A(n_330),
.B(n_342),
.C(n_270),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_266),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_332),
.A2(n_247),
.B1(n_277),
.B2(n_275),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_289),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_334),
.A2(n_339),
.B1(n_249),
.B2(n_255),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_272),
.B(n_11),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_335),
.B(n_340),
.Y(n_382)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_241),
.Y(n_336)
);

BUFx24_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_337),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_238),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_341),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_251),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_272),
.B(n_9),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_241),
.Y(n_341)
);

AND2x6_ASAP7_75t_L g342 ( 
.A(n_254),
.B(n_10),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_253),
.A2(n_250),
.B1(n_263),
.B2(n_282),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_343),
.A2(n_265),
.B1(n_238),
.B2(n_258),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_321),
.A2(n_243),
.B1(n_287),
.B2(n_257),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_345),
.B(n_348),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g346 ( 
.A1(n_316),
.A2(n_321),
.B(n_323),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_346),
.A2(n_379),
.B(n_348),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_351),
.A2(n_340),
.B1(n_335),
.B2(n_330),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_239),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_354),
.B(n_361),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_322),
.A2(n_243),
.B(n_274),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_355),
.Y(n_403)
);

OAI21xp33_ASAP7_75t_SL g425 ( 
.A1(n_357),
.A2(n_371),
.B(n_370),
.Y(n_425)
);

OAI22x1_ASAP7_75t_SL g360 ( 
.A1(n_334),
.A2(n_255),
.B1(n_273),
.B2(n_246),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_306),
.B(n_291),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_331),
.B(n_285),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_363),
.B(n_376),
.C(n_355),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_318),
.B(n_274),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_374),
.Y(n_402)
);

OA22x2_ASAP7_75t_L g368 ( 
.A1(n_334),
.A2(n_246),
.B1(n_271),
.B2(n_277),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g417 ( 
.A1(n_368),
.A2(n_353),
.B(n_360),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_306),
.B(n_271),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_373),
.B(n_304),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_299),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_322),
.B(n_283),
.C(n_331),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_303),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_380),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_322),
.A2(n_301),
.B(n_296),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_303),
.B(n_309),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_327),
.B(n_343),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_298),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_323),
.A2(n_313),
.B1(n_334),
.B2(n_339),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_387),
.A2(n_365),
.B1(n_347),
.B2(n_334),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_350),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_388),
.B(n_389),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_352),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_390),
.B(n_411),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_391),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_392),
.B(n_416),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_359),
.B(n_361),
.Y(n_393)
);

CKINVDCx14_ASAP7_75t_R g436 ( 
.A(n_393),
.Y(n_436)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_381),
.Y(n_394)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_394),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_395),
.B(n_372),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_379),
.A2(n_311),
.B1(n_342),
.B2(n_319),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_396),
.A2(n_420),
.B1(n_422),
.B2(n_368),
.Y(n_450)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_381),
.Y(n_397)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_397),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_358),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_398),
.B(n_400),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_359),
.B(n_310),
.Y(n_399)
);

OAI21xp33_ASAP7_75t_L g442 ( 
.A1(n_399),
.A2(n_407),
.B(n_408),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_341),
.Y(n_400)
);

CKINVDCx12_ASAP7_75t_R g401 ( 
.A(n_385),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_401),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_344),
.B(n_337),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_406),
.B(n_421),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_347),
.B(n_315),
.Y(n_407)
);

OAI21xp33_ASAP7_75t_L g408 ( 
.A1(n_356),
.A2(n_300),
.B(n_333),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_367),
.Y(n_409)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_409),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_365),
.A2(n_305),
.B1(n_337),
.B2(n_356),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_412),
.Y(n_445)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_384),
.Y(n_413)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_413),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_383),
.B(n_363),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_415),
.B(n_418),
.C(n_386),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_374),
.B(n_385),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_417),
.A2(n_362),
.B(n_349),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_384),
.A2(n_346),
.B1(n_373),
.B2(n_387),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_425),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_346),
.A2(n_376),
.B1(n_369),
.B2(n_344),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_369),
.B(n_345),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_358),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_424),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_346),
.B(n_382),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_416),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_426),
.A2(n_433),
.B1(n_451),
.B2(n_453),
.Y(n_474)
);

FAx1_ASAP7_75t_SL g427 ( 
.A(n_418),
.B(n_372),
.CI(n_382),
.CON(n_427),
.SN(n_427)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_414),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_410),
.A2(n_357),
.B1(n_368),
.B2(n_375),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_428),
.A2(n_390),
.B1(n_417),
.B2(n_396),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_424),
.A2(n_375),
.B(n_370),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_431),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_402),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_452),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_SL g440 ( 
.A1(n_404),
.A2(n_403),
.B1(n_398),
.B2(n_388),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_440),
.A2(n_450),
.B1(n_422),
.B2(n_410),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_424),
.A2(n_378),
.B(n_368),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_456),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_393),
.B(n_378),
.Y(n_448)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_448),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_402),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_419),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_386),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_405),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_349),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_455),
.B(n_458),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_395),
.B(n_420),
.C(n_405),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_413),
.Y(n_459)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_459),
.Y(n_477)
);

XNOR2x1_ASAP7_75t_L g501 ( 
.A(n_462),
.B(n_457),
.Y(n_501)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_439),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_463),
.B(n_476),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_457),
.A2(n_417),
.B(n_423),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_464),
.B(n_466),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_453),
.A2(n_432),
.B1(n_428),
.B2(n_443),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_467),
.B(n_488),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_399),
.Y(n_469)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_470),
.A2(n_437),
.B1(n_456),
.B2(n_431),
.Y(n_498)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_444),
.Y(n_471)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_471),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_485),
.Y(n_491)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_444),
.Y(n_473)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_473),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_457),
.A2(n_417),
.B(n_407),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_439),
.Y(n_478)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_478),
.Y(n_502)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_479),
.Y(n_506)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_430),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_482),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_446),
.A2(n_389),
.B1(n_392),
.B2(n_411),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_481),
.Y(n_510)
);

NOR2x1_ASAP7_75t_L g482 ( 
.A(n_436),
.B(n_391),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_394),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_483),
.Y(n_507)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_449),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_484),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_452),
.B(n_397),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_432),
.A2(n_409),
.B1(n_412),
.B2(n_362),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_486),
.A2(n_441),
.B1(n_442),
.B2(n_429),
.Y(n_494)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_447),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_446),
.A2(n_349),
.B1(n_401),
.B2(n_433),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_454),
.C(n_458),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_492),
.B(n_493),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_460),
.B(n_435),
.C(n_426),
.Y(n_493)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_494),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_460),
.B(n_437),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_497),
.B(n_505),
.Y(n_526)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_498),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_475),
.B(n_447),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_499),
.B(n_474),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_501),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_471),
.A2(n_429),
.B1(n_434),
.B2(n_459),
.Y(n_503)
);

OAI22x1_ASAP7_75t_L g524 ( 
.A1(n_503),
.A2(n_509),
.B1(n_484),
.B2(n_465),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_472),
.B(n_427),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_473),
.A2(n_434),
.B1(n_438),
.B2(n_445),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_512),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_503),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_513),
.B(n_519),
.Y(n_541)
);

BUFx12_ASAP7_75t_L g517 ( 
.A(n_507),
.Y(n_517)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_517),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_518),
.Y(n_540)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_502),
.Y(n_519)
);

OA21x2_ASAP7_75t_SL g521 ( 
.A1(n_506),
.A2(n_427),
.B(n_483),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_521),
.A2(n_527),
.B1(n_508),
.B2(n_500),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_493),
.B(n_461),
.C(n_468),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_522),
.B(n_525),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_524),
.B(n_494),
.Y(n_532)
);

INVx8_ASAP7_75t_L g525 ( 
.A(n_510),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_509),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_492),
.B(n_461),
.C(n_468),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_528),
.B(n_530),
.C(n_497),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_469),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_529),
.B(n_531),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_491),
.B(n_461),
.C(n_467),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_486),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_532),
.B(n_536),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_533),
.A2(n_534),
.B1(n_537),
.B2(n_517),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_515),
.A2(n_462),
.B1(n_498),
.B2(n_489),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_525),
.A2(n_495),
.B1(n_496),
.B2(n_504),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_491),
.C(n_504),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_538),
.B(n_543),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_526),
.B(n_530),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_542),
.B(n_536),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_505),
.C(n_501),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_SL g545 ( 
.A(n_526),
.B(n_490),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_545),
.B(n_517),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_520),
.B(n_482),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_546),
.A2(n_529),
.B(n_476),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_515),
.A2(n_523),
.B1(n_527),
.B2(n_514),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_547),
.A2(n_535),
.B1(n_523),
.B2(n_531),
.Y(n_548)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_548),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_538),
.B(n_516),
.C(n_524),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_549),
.B(n_554),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_551),
.B(n_553),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_464),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_519),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_555),
.B(n_558),
.Y(n_561)
);

INVx11_ASAP7_75t_L g556 ( 
.A(n_544),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_556),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_557),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_543),
.B(n_438),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_559),
.A2(n_541),
.B(n_534),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_562),
.A2(n_549),
.B(n_559),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_564),
.B(n_551),
.C(n_550),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_567),
.B(n_570),
.Y(n_571)
);

OAI21x1_ASAP7_75t_SL g568 ( 
.A1(n_566),
.A2(n_556),
.B(n_552),
.Y(n_568)
);

AOI21x1_ASAP7_75t_SL g572 ( 
.A1(n_568),
.A2(n_569),
.B(n_561),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_565),
.A2(n_540),
.B1(n_547),
.B2(n_532),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_572),
.B(n_563),
.C(n_553),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_567),
.B(n_560),
.C(n_563),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_573),
.B(n_550),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_574),
.B(n_575),
.C(n_571),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_576),
.B(n_545),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_577),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_445),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_579),
.B(n_477),
.Y(n_580)
);


endmodule