module real_aes_15674_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_0), .Y(n_562) );
AND2x4_ASAP7_75t_L g112 ( .A(n_1), .B(n_113), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_2), .A2(n_4), .B1(n_288), .B2(n_289), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_3), .A2(n_21), .B1(n_215), .B2(n_224), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_5), .A2(n_52), .B1(n_173), .B2(n_174), .Y(n_172) );
BUFx3_ASAP7_75t_L g513 ( .A(n_6), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_7), .A2(n_15), .B1(n_145), .B2(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_9), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_10), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_11), .B(n_198), .Y(n_519) );
BUFx2_ASAP7_75t_L g104 ( .A(n_12), .Y(n_104) );
OR2x2_ASAP7_75t_L g122 ( .A(n_12), .B(n_30), .Y(n_122) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_13), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_14), .Y(n_847) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_16), .B(n_180), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_17), .B(n_189), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_18), .A2(n_84), .B1(n_180), .B2(n_224), .Y(n_577) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_19), .A2(n_47), .B(n_158), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_20), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_22), .B(n_215), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_23), .B(n_150), .Y(n_244) );
INVx4_ASAP7_75t_R g197 ( .A(n_24), .Y(n_197) );
AO32x2_ASAP7_75t_L g574 ( .A1(n_25), .A2(n_226), .A3(n_227), .B1(n_575), .B2(n_578), .Y(n_574) );
AO32x1_ASAP7_75t_L g596 ( .A1(n_25), .A2(n_226), .A3(n_227), .B1(n_575), .B2(n_578), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_26), .B(n_215), .Y(n_250) );
INVx1_ASAP7_75t_L g293 ( .A(n_27), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_SL g221 ( .A1(n_28), .A2(n_145), .B(n_149), .C(n_222), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_29), .A2(n_44), .B1(n_145), .B2(n_152), .Y(n_233) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_30), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_31), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_32), .A2(n_51), .B1(n_199), .B2(n_215), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_33), .A2(n_89), .B1(n_152), .B2(n_224), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_34), .B(n_521), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_35), .B(n_543), .Y(n_587) );
INVx1_ASAP7_75t_L g247 ( .A(n_36), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_37), .B(n_145), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_38), .A2(n_67), .B1(n_152), .B2(n_568), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_39), .Y(n_266) );
INVx2_ASAP7_75t_L g127 ( .A(n_40), .Y(n_127) );
INVx1_ASAP7_75t_L g107 ( .A(n_41), .Y(n_107) );
BUFx3_ASAP7_75t_L g130 ( .A(n_41), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_42), .A2(n_100), .B1(n_114), .B2(n_854), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_43), .B(n_589), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_45), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_46), .A2(n_83), .B1(n_145), .B2(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_48), .B(n_837), .Y(n_836) );
OAI31xp67_ASAP7_75t_SL g842 ( .A1(n_48), .A2(n_838), .A3(n_840), .B(n_843), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_49), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_50), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_53), .A2(n_77), .B1(n_182), .B2(n_543), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_54), .Y(n_163) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_55), .A2(n_81), .B1(n_180), .B2(n_224), .Y(n_509) );
INVx1_ASAP7_75t_L g158 ( .A(n_56), .Y(n_158) );
AND2x4_ASAP7_75t_L g160 ( .A(n_57), .B(n_161), .Y(n_160) );
XNOR2xp5_ASAP7_75t_L g131 ( .A(n_58), .B(n_132), .Y(n_131) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_59), .A2(n_88), .B1(n_152), .B2(n_286), .Y(n_285) );
AO22x1_ASAP7_75t_L g178 ( .A1(n_60), .A2(n_72), .B1(n_179), .B2(n_181), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_61), .B(n_224), .Y(n_518) );
INVx1_ASAP7_75t_L g161 ( .A(n_62), .Y(n_161) );
AND2x2_ASAP7_75t_L g225 ( .A(n_63), .B(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_64), .B(n_226), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_65), .A2(n_170), .B(n_173), .C(n_561), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_66), .B(n_224), .C(n_523), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_68), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_69), .B(n_173), .Y(n_272) );
AND2x2_ASAP7_75t_L g563 ( .A(n_70), .B(n_203), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_71), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_73), .B(n_215), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_74), .A2(n_94), .B1(n_180), .B2(n_182), .Y(n_545) );
INVx2_ASAP7_75t_L g150 ( .A(n_75), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_76), .B(n_268), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_78), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_79), .B(n_226), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_80), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_82), .B(n_156), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_85), .B(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_86), .A2(n_98), .B1(n_152), .B2(n_199), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_87), .B(n_543), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_90), .B(n_226), .Y(n_263) );
INVx1_ASAP7_75t_L g111 ( .A(n_91), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_91), .B(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_92), .B(n_189), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_93), .A2(n_154), .B(n_173), .C(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g202 ( .A(n_95), .B(n_203), .Y(n_202) );
NAND2xp33_ASAP7_75t_L g271 ( .A(n_96), .B(n_198), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_97), .Y(n_532) );
BUFx10_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
BUFx12f_ASAP7_75t_L g855 ( .A(n_101), .Y(n_855) );
NOR2x1p5_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_103), .B(n_104), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g120 ( .A(n_107), .Y(n_120) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g498 ( .A(n_111), .Y(n_498) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_123), .Y(n_114) );
INVxp67_ASAP7_75t_L g843 ( .A(n_115), .Y(n_843) );
NOR2x1_ASAP7_75t_R g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
CKINVDCx8_ASAP7_75t_R g839 ( .A(n_118), .Y(n_839) );
AND2x6_ASAP7_75t_SL g118 ( .A(n_119), .B(n_121), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_121), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NOR2x1_ASAP7_75t_L g853 ( .A(n_122), .B(n_130), .Y(n_853) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_131), .B(n_834), .Y(n_123) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x6_ASAP7_75t_SL g125 ( .A(n_126), .B(n_128), .Y(n_125) );
BUFx3_ASAP7_75t_L g845 ( .A(n_126), .Y(n_845) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_127), .B(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AOI22x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_496), .B1(n_499), .B2(n_833), .Y(n_132) );
INVx2_ASAP7_75t_L g841 ( .A(n_133), .Y(n_841) );
NOR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_410), .Y(n_133) );
NAND4xp75_ASAP7_75t_L g134 ( .A(n_135), .B(n_315), .C(n_357), .D(n_381), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI211xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_204), .B(n_252), .C(n_294), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g401 ( .A(n_139), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g495 ( .A(n_139), .B(n_432), .Y(n_495) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_165), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g310 ( .A(n_141), .B(n_262), .Y(n_310) );
AND2x2_ASAP7_75t_L g351 ( .A(n_141), .B(n_312), .Y(n_351) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g258 ( .A(n_142), .B(n_187), .Y(n_258) );
OR2x2_ASAP7_75t_L g276 ( .A(n_142), .B(n_187), .Y(n_276) );
INVx2_ASAP7_75t_L g302 ( .A(n_142), .Y(n_302) );
AND2x2_ASAP7_75t_L g332 ( .A(n_142), .B(n_262), .Y(n_332) );
AND2x2_ASAP7_75t_L g361 ( .A(n_142), .B(n_186), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_142), .B(n_313), .Y(n_397) );
AO31x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_155), .A3(n_159), .B(n_162), .Y(n_142) );
OAI22x1_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_148), .B1(n_151), .B2(n_153), .Y(n_143) );
INVx4_ASAP7_75t_L g147 ( .A(n_145), .Y(n_147) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVx1_ASAP7_75t_L g173 ( .A(n_146), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_146), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_146), .Y(n_199) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_146), .Y(n_215) );
INVx1_ASAP7_75t_L g217 ( .A(n_146), .Y(n_217) );
INVx2_ASAP7_75t_L g224 ( .A(n_146), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_147), .A2(n_266), .B(n_267), .C(n_268), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_148), .A2(n_169), .B1(n_232), .B2(n_233), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_148), .A2(n_153), .B1(n_285), .B2(n_287), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_148), .A2(n_149), .B1(n_509), .B2(n_510), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_148), .A2(n_542), .B1(n_544), .B2(n_545), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_148), .A2(n_169), .B1(n_567), .B2(n_569), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_148), .A2(n_587), .B(n_588), .Y(n_586) );
INVx6_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_149), .B(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_149), .A2(n_271), .B(n_272), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_149), .A2(n_168), .B(n_178), .C(n_184), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_149), .A2(n_518), .B(n_519), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_149), .A2(n_219), .B1(n_576), .B2(n_577), .Y(n_575) );
BUFx8_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g154 ( .A(n_150), .Y(n_154) );
INVx2_ASAP7_75t_L g171 ( .A(n_150), .Y(n_171) );
INVx1_ASAP7_75t_L g220 ( .A(n_150), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_152), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g288 ( .A(n_152), .Y(n_288) );
INVx2_ASAP7_75t_L g521 ( .A(n_152), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_153), .B(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_SL g544 ( .A(n_154), .Y(n_544) );
INVx1_ASAP7_75t_L g559 ( .A(n_154), .Y(n_559) );
INVx2_ASAP7_75t_L g515 ( .A(n_155), .Y(n_515) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g164 ( .A(n_156), .Y(n_164) );
OAI21xp33_ASAP7_75t_L g184 ( .A1(n_156), .A2(n_176), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_157), .Y(n_227) );
INVx2_ASAP7_75t_L g201 ( .A(n_159), .Y(n_201) );
BUFx10_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g185 ( .A(n_160), .Y(n_185) );
BUFx10_ASAP7_75t_L g235 ( .A(n_160), .Y(n_235) );
INVx1_ASAP7_75t_L g291 ( .A(n_160), .Y(n_291) );
AO31x2_ASAP7_75t_L g565 ( .A1(n_160), .A2(n_540), .A3(n_566), .B(n_570), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
INVx2_ASAP7_75t_L g203 ( .A(n_164), .Y(n_203) );
BUFx2_ASAP7_75t_L g210 ( .A(n_164), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_164), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_164), .B(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_164), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g374 ( .A(n_165), .B(n_303), .Y(n_374) );
INVx2_ASAP7_75t_L g469 ( .A(n_165), .Y(n_469) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_186), .Y(n_165) );
INVx2_ASAP7_75t_L g257 ( .A(n_166), .Y(n_257) );
AND2x4_ASAP7_75t_L g300 ( .A(n_166), .B(n_187), .Y(n_300) );
AOI21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_177), .B(n_183), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_176), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_169), .A2(n_249), .B(n_250), .Y(n_248) );
AOI21x1_ASAP7_75t_L g583 ( .A1(n_169), .A2(n_584), .B(n_585), .Y(n_583) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g269 ( .A(n_171), .Y(n_269) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_175), .B(n_194), .Y(n_193) );
INVxp67_ASAP7_75t_SL g179 ( .A(n_180), .Y(n_179) );
INVx3_ASAP7_75t_L g589 ( .A(n_180), .Y(n_589) );
OAI21xp33_ASAP7_75t_SL g243 ( .A1(n_181), .A2(n_244), .B(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_182), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_185), .A2(n_212), .B(n_221), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_185), .A2(n_555), .B(n_560), .Y(n_554) );
AND2x2_ASAP7_75t_L g459 ( .A(n_186), .B(n_257), .Y(n_459) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g323 ( .A(n_187), .Y(n_323) );
AND2x2_ASAP7_75t_L g380 ( .A(n_187), .B(n_262), .Y(n_380) );
AND2x2_ASAP7_75t_L g395 ( .A(n_187), .B(n_303), .Y(n_395) );
AND2x2_ASAP7_75t_L g417 ( .A(n_187), .B(n_257), .Y(n_417) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_191), .B(n_202), .Y(n_187) );
AOI21x1_ASAP7_75t_L g553 ( .A1(n_188), .A2(n_554), .B(n_563), .Y(n_553) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_195), .B(n_201), .Y(n_191) );
OAI22xp33_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B1(n_199), .B2(n_200), .Y(n_196) );
INVx2_ASAP7_75t_L g286 ( .A(n_198), .Y(n_286) );
INVx1_ASAP7_75t_L g536 ( .A(n_199), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_199), .A2(n_215), .B1(n_557), .B2(n_558), .Y(n_556) );
OAI211xp5_ASAP7_75t_SL g464 ( .A1(n_204), .A2(n_465), .B(n_467), .C(n_474), .Y(n_464) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_238), .Y(n_205) );
INVxp67_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g451 ( .A(n_207), .B(n_387), .Y(n_451) );
OR2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_228), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_208), .B(n_240), .Y(n_350) );
INVxp67_ASAP7_75t_L g364 ( .A(n_208), .Y(n_364) );
AND2x2_ASAP7_75t_L g384 ( .A(n_208), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_208), .B(n_297), .Y(n_391) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g280 ( .A(n_209), .Y(n_280) );
AOI21x1_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_225), .Y(n_209) );
AO31x2_ASAP7_75t_L g283 ( .A1(n_210), .A2(n_284), .A3(n_290), .B(n_292), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_216), .B(n_219), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g568 ( .A(n_215), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g289 ( .A(n_217), .Y(n_289) );
O2A1O1Ixp5_ASAP7_75t_L g531 ( .A1(n_219), .A2(n_289), .B(n_532), .C(n_533), .Y(n_531) );
BUFx4f_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_220), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g523 ( .A(n_220), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
INVx2_ASAP7_75t_SL g543 ( .A(n_224), .Y(n_543) );
INVx2_ASAP7_75t_L g234 ( .A(n_226), .Y(n_234) );
NOR2x1_ASAP7_75t_L g273 ( .A(n_226), .B(n_274), .Y(n_273) );
INVx4_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g251 ( .A(n_227), .B(n_235), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_227), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g529 ( .A(n_227), .Y(n_529) );
BUFx3_ASAP7_75t_L g540 ( .A(n_227), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_227), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_SL g581 ( .A(n_227), .Y(n_581) );
OR2x2_ASAP7_75t_L g325 ( .A(n_228), .B(n_307), .Y(n_325) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g373 ( .A(n_229), .B(n_280), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_229), .B(n_283), .Y(n_379) );
INVx2_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g279 ( .A(n_230), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g348 ( .A(n_230), .B(n_283), .Y(n_348) );
BUFx2_ASAP7_75t_L g355 ( .A(n_230), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_230), .B(n_283), .Y(n_435) );
AO31x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_234), .A3(n_235), .B(n_236), .Y(n_230) );
AOI31xp67_ASAP7_75t_L g507 ( .A1(n_234), .A2(n_235), .A3(n_508), .B(n_511), .Y(n_507) );
INVx1_ASAP7_75t_L g274 ( .A(n_235), .Y(n_274) );
OAI21x1_ASAP7_75t_L g516 ( .A1(n_235), .A2(n_517), .B(n_520), .Y(n_516) );
OAI21x1_ASAP7_75t_L g530 ( .A1(n_235), .A2(n_531), .B(n_534), .Y(n_530) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x4_ASAP7_75t_L g365 ( .A(n_239), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g494 ( .A(n_239), .B(n_279), .Y(n_494) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx3_ASAP7_75t_L g297 ( .A(n_240), .Y(n_297) );
AND2x2_ASAP7_75t_L g308 ( .A(n_240), .B(n_283), .Y(n_308) );
AND2x2_ASAP7_75t_L g354 ( .A(n_240), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g387 ( .A(n_240), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_240), .B(n_298), .Y(n_404) );
AND2x2_ASAP7_75t_L g443 ( .A(n_240), .B(n_444), .Y(n_443) );
AND2x4_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_248), .B(n_251), .Y(n_242) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_259), .B(n_277), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_254), .A2(n_422), .B1(n_423), .B2(n_425), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
AND2x2_ASAP7_75t_L g419 ( .A(n_255), .B(n_310), .Y(n_419) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g334 ( .A(n_256), .Y(n_334) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g483 ( .A(n_257), .B(n_303), .Y(n_483) );
AND2x2_ASAP7_75t_L g447 ( .A(n_258), .B(n_342), .Y(n_447) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_275), .Y(n_259) );
OR2x2_ASAP7_75t_L g344 ( .A(n_260), .B(n_321), .Y(n_344) );
OR2x2_ASAP7_75t_L g456 ( .A(n_260), .B(n_276), .Y(n_456) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g319 ( .A(n_261), .Y(n_319) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g303 ( .A(n_262), .Y(n_303) );
BUFx3_ASAP7_75t_L g385 ( .A(n_262), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_270), .B(n_273), .Y(n_264) );
INVx2_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_269), .A2(n_535), .B1(n_536), .B2(n_537), .Y(n_534) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g453 ( .A(n_276), .B(n_312), .Y(n_453) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
AND2x2_ASAP7_75t_L g295 ( .A(n_279), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g336 ( .A(n_279), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g473 ( .A(n_279), .Y(n_473) );
INVx1_ASAP7_75t_L g492 ( .A(n_279), .Y(n_492) );
INVx2_ASAP7_75t_L g307 ( .A(n_280), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_280), .B(n_283), .Y(n_356) );
INVx1_ASAP7_75t_L g420 ( .A(n_281), .Y(n_420) );
BUFx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g481 ( .A(n_282), .Y(n_481) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g298 ( .A(n_283), .Y(n_298) );
INVx1_ASAP7_75t_L g388 ( .A(n_283), .Y(n_388) );
AO31x2_ASAP7_75t_L g539 ( .A1(n_290), .A2(n_540), .A3(n_541), .B(n_546), .Y(n_539) );
INVx2_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_SL g578 ( .A(n_291), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_299), .B1(n_304), .B2(n_309), .Y(n_294) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx2_ASAP7_75t_L g337 ( .A(n_297), .Y(n_337) );
AND2x2_ASAP7_75t_L g339 ( .A(n_297), .B(n_324), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_297), .B(n_307), .Y(n_399) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx3_ASAP7_75t_L g330 ( .A(n_300), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_300), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g424 ( .A(n_300), .B(n_408), .Y(n_424) );
INVx1_ASAP7_75t_L g328 ( .A(n_301), .Y(n_328) );
AOI222xp33_ASAP7_75t_L g338 ( .A1(n_301), .A2(n_339), .B1(n_340), .B2(n_345), .C1(n_351), .C2(n_352), .Y(n_338) );
OAI21xp33_ASAP7_75t_SL g368 ( .A1(n_301), .A2(n_369), .B(n_370), .Y(n_368) );
AND2x2_ASAP7_75t_L g392 ( .A(n_301), .B(n_311), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_301), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
OR2x2_ASAP7_75t_L g321 ( .A(n_302), .B(n_313), .Y(n_321) );
INVx1_ASAP7_75t_L g409 ( .A(n_302), .Y(n_409) );
BUFx2_ASAP7_75t_L g343 ( .A(n_303), .Y(n_343) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_306), .B(n_347), .Y(n_376) );
OR2x2_ASAP7_75t_L g488 ( .A(n_306), .B(n_348), .Y(n_488) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g371 ( .A(n_308), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g486 ( .A(n_308), .Y(n_486) );
OAI31xp33_ASAP7_75t_L g467 ( .A1(n_309), .A2(n_468), .A3(n_470), .B(n_471), .Y(n_467) );
AND2x4_ASAP7_75t_SL g309 ( .A(n_310), .B(n_311), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_310), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_338), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_324), .B(n_326), .Y(n_316) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x6_ASAP7_75t_L g437 ( .A(n_319), .B(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g369 ( .A(n_322), .Y(n_369) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g460 ( .A(n_323), .B(n_397), .Y(n_460) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_325), .A2(n_414), .B1(n_416), .B2(n_418), .Y(n_413) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_325), .A2(n_386), .B(n_448), .C(n_475), .Y(n_474) );
AOI21xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_331), .B(n_335), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND4xp25_ASAP7_75t_L g427 ( .A(n_330), .B(n_428), .C(n_429), .D(n_431), .Y(n_427) );
NAND2x1_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_332), .B(n_334), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_332), .B(n_417), .Y(n_440) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g406 ( .A(n_337), .B(n_366), .Y(n_406) );
NAND2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_344), .A2(n_488), .B1(n_489), .B2(n_491), .Y(n_487) );
AOI221x1_ASAP7_75t_L g426 ( .A1(n_345), .A2(n_427), .B1(n_433), .B2(n_436), .C(n_439), .Y(n_426) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g366 ( .A(n_348), .Y(n_366) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g378 ( .A(n_350), .B(n_379), .Y(n_378) );
NAND2x1p5_ASAP7_75t_L g441 ( .A(n_351), .B(n_432), .Y(n_441) );
O2A1O1Ixp5_ASAP7_75t_L g454 ( .A1(n_352), .A2(n_436), .B(n_455), .C(n_457), .Y(n_454) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx2_ASAP7_75t_L g403 ( .A(n_355), .Y(n_403) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_367), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_362), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g446 ( .A1(n_359), .A2(n_377), .B1(n_447), .B2(n_448), .C(n_450), .Y(n_446) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g383 ( .A(n_361), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_361), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g482 ( .A(n_361), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
NAND2x1_ASAP7_75t_L g461 ( .A(n_364), .B(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g485 ( .A(n_364), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g425 ( .A(n_365), .Y(n_425) );
AOI222xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .B1(n_374), .B2(n_375), .C1(n_377), .C2(n_380), .Y(n_367) );
INVx1_ASAP7_75t_L g452 ( .A(n_371), .Y(n_452) );
INVx1_ASAP7_75t_L g415 ( .A(n_372), .Y(n_415) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g449 ( .A(n_373), .Y(n_449) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g390 ( .A(n_379), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g444 ( .A(n_379), .Y(n_444) );
AND2x2_ASAP7_75t_L g407 ( .A(n_380), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_400), .Y(n_381) );
AOI222xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .B1(n_389), .B2(n_392), .C1(n_393), .C2(n_398), .Y(n_382) );
INVx3_ASAP7_75t_L g432 ( .A(n_385), .Y(n_432) );
BUFx2_ASAP7_75t_L g490 ( .A(n_385), .Y(n_490) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g462 ( .A(n_387), .Y(n_462) );
OR2x2_ASAP7_75t_L g472 ( .A(n_387), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx2_ASAP7_75t_SL g430 ( .A(n_395), .Y(n_430) );
AND2x2_ASAP7_75t_L g475 ( .A(n_396), .B(n_432), .Y(n_475) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g434 ( .A(n_399), .B(n_435), .Y(n_434) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_401), .B(n_405), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
OR2x2_ASAP7_75t_L g491 ( .A(n_404), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g422 ( .A(n_406), .Y(n_422) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g429 ( .A(n_409), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g479 ( .A(n_409), .Y(n_479) );
NAND4xp75_ASAP7_75t_L g410 ( .A(n_411), .B(n_445), .C(n_463), .D(n_476), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_426), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_420), .B(n_421), .Y(n_412) );
INVxp33_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_415), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g438 ( .A(n_417), .Y(n_438) );
AND2x2_ASAP7_75t_L g478 ( .A(n_417), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g448 ( .A(n_420), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g466 ( .A(n_431), .Y(n_466) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI22xp33_ASAP7_75t_SL g457 ( .A1(n_434), .A2(n_458), .B1(n_460), .B2(n_461), .Y(n_457) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI21xp33_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_441), .B(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g470 ( .A(n_441), .Y(n_470) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_454), .Y(n_445) );
AOI21xp5_ASAP7_75t_SL g450 ( .A1(n_451), .A2(n_452), .B(n_453), .Y(n_450) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_493), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_480), .B1(n_482), .B2(n_484), .C(n_487), .Y(n_477) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx4_ASAP7_75t_L g833 ( .A(n_496), .Y(n_833) );
BUFx12f_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g852 ( .A(n_498), .B(n_853), .Y(n_852) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_734), .Y(n_499) );
AND4x1_ASAP7_75t_L g500 ( .A(n_501), .B(n_656), .C(n_689), .D(n_720), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_623), .Y(n_501) );
OAI221xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_548), .B1(n_591), .B2(n_601), .C(n_610), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g728 ( .A1(n_503), .A2(n_713), .B(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_526), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
INVx2_ASAP7_75t_L g609 ( .A(n_506), .Y(n_609) );
AND2x2_ASAP7_75t_L g619 ( .A(n_506), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g655 ( .A(n_506), .B(n_539), .Y(n_655) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g644 ( .A(n_507), .Y(n_644) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g630 ( .A(n_514), .B(n_620), .Y(n_630) );
OR2x2_ASAP7_75t_L g739 ( .A(n_514), .B(n_528), .Y(n_739) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_525), .Y(n_514) );
OAI21x1_ASAP7_75t_L g608 ( .A1(n_515), .A2(n_516), .B(n_525), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_524), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_526), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
INVx1_ASAP7_75t_L g604 ( .A(n_528), .Y(n_604) );
INVx2_ASAP7_75t_SL g681 ( .A(n_528), .Y(n_681) );
BUFx2_ASAP7_75t_L g711 ( .A(n_528), .Y(n_711) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_538), .Y(n_528) );
OA21x2_ASAP7_75t_L g620 ( .A1(n_529), .A2(n_530), .B(n_538), .Y(n_620) );
AND2x2_ASAP7_75t_L g603 ( .A(n_539), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g622 ( .A(n_539), .Y(n_622) );
OR2x2_ASAP7_75t_L g642 ( .A(n_539), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g683 ( .A(n_539), .Y(n_683) );
INVx1_ASAP7_75t_L g694 ( .A(n_539), .Y(n_694) );
AND2x2_ASAP7_75t_L g701 ( .A(n_539), .B(n_643), .Y(n_701) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g549 ( .A(n_550), .B(n_572), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_564), .Y(n_550) );
INVx1_ASAP7_75t_L g615 ( .A(n_551), .Y(n_615) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_552), .Y(n_627) );
INVx1_ASAP7_75t_L g636 ( .A(n_552), .Y(n_636) );
INVx1_ASAP7_75t_L g675 ( .A(n_552), .Y(n_675) );
AND2x2_ASAP7_75t_L g705 ( .A(n_552), .B(n_565), .Y(n_705) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g599 ( .A(n_553), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_556), .B(n_559), .Y(n_555) );
INVx1_ASAP7_75t_L g611 ( .A(n_564), .Y(n_611) );
AND2x4_ASAP7_75t_L g660 ( .A(n_564), .B(n_574), .Y(n_660) );
AND2x2_ASAP7_75t_L g670 ( .A(n_564), .B(n_599), .Y(n_670) );
INVx1_ASAP7_75t_L g731 ( .A(n_564), .Y(n_731) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g617 ( .A(n_565), .B(n_596), .Y(n_617) );
AND2x2_ASAP7_75t_L g635 ( .A(n_565), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g651 ( .A(n_565), .B(n_596), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_565), .B(n_579), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_572), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_579), .Y(n_572) );
OR2x2_ASAP7_75t_L g777 ( .A(n_573), .B(n_579), .Y(n_777) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g724 ( .A(n_574), .Y(n_724) );
AND2x2_ASAP7_75t_L g749 ( .A(n_574), .B(n_579), .Y(n_749) );
OAI21x1_ASAP7_75t_L g582 ( .A1(n_578), .A2(n_583), .B(n_586), .Y(n_582) );
INVx3_ASAP7_75t_L g600 ( .A(n_579), .Y(n_600) );
AND2x2_ASAP7_75t_L g626 ( .A(n_579), .B(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g648 ( .A(n_579), .Y(n_648) );
INVx1_ASAP7_75t_L g662 ( .A(n_579), .Y(n_662) );
INVx1_ASAP7_75t_L g672 ( .A(n_579), .Y(n_672) );
BUFx2_ASAP7_75t_L g767 ( .A(n_579), .Y(n_767) );
OR2x2_ASAP7_75t_L g795 ( .A(n_579), .B(n_599), .Y(n_795) );
INVxp67_ASAP7_75t_L g812 ( .A(n_579), .Y(n_812) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B(n_590), .Y(n_580) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_597), .Y(n_592) );
AND2x4_ASAP7_75t_L g625 ( .A(n_593), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_593), .B(n_705), .Y(n_786) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g613 ( .A(n_595), .B(n_600), .Y(n_613) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_595), .Y(n_637) );
INVx1_ASAP7_75t_L g761 ( .A(n_595), .Y(n_761) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g674 ( .A(n_596), .Y(n_674) );
AND2x2_ASAP7_75t_L g688 ( .A(n_597), .B(n_651), .Y(n_688) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g650 ( .A(n_599), .Y(n_650) );
OR2x2_ASAP7_75t_L g708 ( .A(n_599), .B(n_674), .Y(n_708) );
INVx1_ASAP7_75t_L g771 ( .A(n_599), .Y(n_771) );
AND2x2_ASAP7_75t_L g714 ( .A(n_600), .B(n_660), .Y(n_714) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x4_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
AND2x2_ASAP7_75t_L g717 ( .A(n_603), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
AND2x2_ASAP7_75t_L g621 ( .A(n_606), .B(n_622), .Y(n_621) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_606), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g640 ( .A(n_607), .Y(n_640) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g719 ( .A(n_608), .B(n_644), .Y(n_719) );
AND2x2_ASAP7_75t_L g682 ( .A(n_609), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g753 ( .A(n_609), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B(n_614), .C(n_618), .Y(n_610) );
INVx1_ASAP7_75t_L g745 ( .A(n_612), .Y(n_745) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_L g741 ( .A(n_613), .B(n_705), .Y(n_741) );
INVx1_ASAP7_75t_L g832 ( .A(n_613), .Y(n_832) );
INVx1_ASAP7_75t_L g797 ( .A(n_614), .Y(n_797) );
AND2x4_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g830 ( .A(n_615), .B(n_749), .Y(n_830) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g647 ( .A(n_617), .B(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g802 ( .A(n_617), .B(n_767), .Y(n_802) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVxp67_ASAP7_75t_L g692 ( .A(n_619), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_619), .B(n_654), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_619), .B(n_621), .Y(n_784) );
INVx1_ASAP7_75t_L g667 ( .A(n_620), .Y(n_667) );
INVx2_ASAP7_75t_SL g632 ( .A(n_622), .Y(n_632) );
OR2x2_ASAP7_75t_L g661 ( .A(n_622), .B(n_662), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_628), .B1(n_633), .B2(n_638), .C(n_645), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR2xp33_ASAP7_75t_SL g669 ( .A(n_625), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g697 ( .A(n_627), .Y(n_697) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g754 ( .A(n_630), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_630), .B(n_632), .Y(n_792) );
OR2x2_ASAP7_75t_L g774 ( .A(n_631), .B(n_764), .Y(n_774) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g743 ( .A(n_632), .B(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g790 ( .A(n_632), .B(n_719), .Y(n_790) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
AND2x2_ASAP7_75t_L g725 ( .A(n_635), .B(n_648), .Y(n_725) );
BUFx2_ASAP7_75t_L g751 ( .A(n_635), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_639), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g654 ( .A(n_640), .Y(n_654) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g727 ( .A(n_642), .Y(n_727) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_649), .B(n_652), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g704 ( .A(n_648), .Y(n_704) );
INVxp67_ASAP7_75t_SL g707 ( .A(n_648), .Y(n_707) );
OR2x2_ASAP7_75t_L g817 ( .A(n_648), .B(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g778 ( .A(n_649), .Y(n_778) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g686 ( .A(n_650), .Y(n_686) );
AND2x2_ASAP7_75t_L g813 ( .A(n_651), .B(n_686), .Y(n_813) );
INVx2_ASAP7_75t_SL g818 ( .A(n_651), .Y(n_818) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx2_ASAP7_75t_L g700 ( .A(n_654), .Y(n_700) );
AND2x4_ASAP7_75t_L g676 ( .A(n_655), .B(n_665), .Y(n_676) );
INVx2_ASAP7_75t_L g740 ( .A(n_655), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_655), .B(n_681), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_655), .B(n_711), .Y(n_827) );
AOI221x1_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_663), .B1(n_668), .B2(n_676), .C(n_677), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVx2_ASAP7_75t_L g796 ( .A(n_659), .Y(n_796) );
AOI21xp33_ASAP7_75t_L g803 ( .A1(n_659), .A2(n_804), .B(n_806), .Y(n_803) );
INVx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g685 ( .A(n_660), .B(n_686), .Y(n_685) );
BUFx2_ASAP7_75t_L g716 ( .A(n_660), .Y(n_716) );
AND2x4_ASAP7_75t_L g770 ( .A(n_660), .B(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g730 ( .A(n_662), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI32xp33_ASAP7_75t_L g775 ( .A1(n_664), .A2(n_773), .A3(n_776), .B1(n_778), .B2(n_779), .Y(n_775) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_665), .B(n_682), .Y(n_798) );
AND2x2_ASAP7_75t_L g814 ( .A(n_665), .B(n_694), .Y(n_814) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_669), .B(n_671), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_670), .B(n_812), .Y(n_811) );
O2A1O1Ixp33_ASAP7_75t_L g746 ( .A1(n_671), .A2(n_747), .B(n_750), .C(n_752), .Y(n_746) );
NAND2x1p5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g695 ( .A(n_673), .Y(n_695) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
OAI21xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_684), .B(n_687), .Y(n_677) );
OAI21xp33_ASAP7_75t_L g712 ( .A1(n_678), .A2(n_713), .B(n_715), .Y(n_712) );
INVx2_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_681), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_685), .A2(n_758), .B1(n_762), .B2(n_763), .Y(n_757) );
AND2x2_ASAP7_75t_L g824 ( .A(n_685), .B(n_812), .Y(n_824) );
NOR2xp33_ASAP7_75t_SL g689 ( .A(n_690), .B(n_712), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_695), .B1(n_696), .B2(n_698), .C(n_702), .Y(n_690) );
AOI21xp33_ASAP7_75t_L g800 ( .A1(n_691), .A2(n_801), .B(n_802), .Y(n_800) );
OR2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
AND2x2_ASAP7_75t_L g783 ( .A(n_697), .B(n_749), .Y(n_783) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
AOI31xp33_ASAP7_75t_L g720 ( .A1(n_700), .A2(n_721), .A3(n_726), .B(n_728), .Y(n_720) );
AND2x2_ASAP7_75t_L g820 ( .A(n_700), .B(n_727), .Y(n_820) );
AND2x2_ASAP7_75t_L g709 ( .A(n_701), .B(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_701), .Y(n_773) );
INVx1_ASAP7_75t_L g807 ( .A(n_701), .Y(n_807) );
OAI21xp33_ASAP7_75t_SL g702 ( .A1(n_703), .A2(n_706), .B(n_709), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx2_ASAP7_75t_L g733 ( .A(n_705), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_705), .B(n_832), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g788 ( .A1(n_706), .A2(n_789), .B(n_791), .Y(n_788) );
NOR2x1p5_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
O2A1O1Ixp33_ASAP7_75t_L g729 ( .A1(n_708), .A2(n_723), .B(n_730), .C(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g742 ( .A(n_711), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g762 ( .A(n_711), .B(n_718), .Y(n_762) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g744 ( .A(n_719), .Y(n_744) );
INVx1_ASAP7_75t_L g780 ( .A(n_719), .Y(n_780) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_725), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_725), .A2(n_742), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g801 ( .A(n_725), .Y(n_801) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NOR2x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_787), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_755), .C(n_765), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_741), .B1(n_742), .B2(n_745), .C(n_746), .Y(n_736) );
INVx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_743), .A2(n_810), .B1(n_813), .B2(n_814), .Y(n_809) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
BUFx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OR2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
OR2x2_ASAP7_75t_L g806 ( .A(n_754), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g805 ( .A(n_760), .Y(n_805) );
INVx2_ASAP7_75t_L g785 ( .A(n_762), .Y(n_785) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AOI211xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_768), .B(n_775), .C(n_781), .Y(n_765) );
BUFx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI21xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_772), .B(n_774), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OR2x2_ASAP7_75t_L g776 ( .A(n_771), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g819 ( .A(n_776), .Y(n_819) );
OAI22xp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NAND4xp75_ASAP7_75t_L g787 ( .A(n_788), .B(n_799), .C(n_808), .D(n_821), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OAI22xp33_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B1(n_797), .B2(n_798), .Y(n_791) );
NAND2x1_ASAP7_75t_SL g793 ( .A(n_794), .B(n_796), .Y(n_793) );
INVx3_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_803), .Y(n_799) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_815), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI21xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_819), .B(n_820), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_824), .B1(n_825), .B2(n_828), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVxp67_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_831), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
A2O1A1O1Ixp25_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_840), .B(n_842), .C(n_844), .D(n_846), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
INVx4_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx3_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
INVx6_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
BUFx10_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
CKINVDCx11_ASAP7_75t_R g854 ( .A(n_855), .Y(n_854) );
endmodule