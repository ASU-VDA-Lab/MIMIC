module fake_ariane_2430_n_960 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_960);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_960;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_936;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_515;
wire n_379;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_857;
wire n_898;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_903;
wire n_871;
wire n_315;
wire n_754;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_218;
wire n_839;
wire n_770;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_458;
wire n_361;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_847;
wire n_939;
wire n_772;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_852;
wire n_793;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_856;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_155),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_96),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_26),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_48),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_55),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_78),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_115),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_40),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_104),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_0),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_72),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_138),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_183),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_142),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_81),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_83),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_118),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_60),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_37),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_38),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_126),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_80),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_85),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_53),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_73),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_26),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_39),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_112),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_128),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_101),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_35),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_141),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_144),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_88),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_56),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_25),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_90),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_109),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_140),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_82),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_15),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_31),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_15),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_166),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_32),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_23),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_70),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_120),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_79),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_135),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_108),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_44),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_92),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_2),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_130),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_10),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_162),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_170),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_134),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_36),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_204),
.Y(n_255)
);

INVxp33_ASAP7_75t_SL g256 ( 
.A(n_189),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_211),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_187),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_211),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_200),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_248),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_187),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_200),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_202),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_185),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_191),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_202),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_193),
.Y(n_279)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_234),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_230),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_194),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_195),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_230),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_237),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_206),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_216),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_217),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_222),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_223),
.Y(n_292)
);

INVxp33_ASAP7_75t_SL g293 ( 
.A(n_227),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_237),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_225),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_244),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_261),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_253),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_273),
.A2(n_244),
.B1(n_238),
.B2(n_240),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_264),
.Y(n_306)
);

OA21x2_ASAP7_75t_L g307 ( 
.A1(n_264),
.A2(n_236),
.B(n_220),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_272),
.B(n_250),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_256),
.A2(n_207),
.B1(n_214),
.B2(n_252),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_258),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_286),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_286),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

BUFx8_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_269),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_260),
.B(n_221),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_272),
.B(n_221),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_256),
.A2(n_251),
.B1(n_247),
.B2(n_245),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_270),
.B(n_0),
.Y(n_325)
);

CKINVDCx8_ASAP7_75t_R g326 ( 
.A(n_274),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_295),
.Y(n_327)
);

AND2x4_ASAP7_75t_L g328 ( 
.A(n_272),
.B(n_221),
.Y(n_328)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

BUFx8_ASAP7_75t_L g330 ( 
.A(n_276),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_259),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_263),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_184),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_255),
.A2(n_243),
.B1(n_242),
.B2(n_186),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_257),
.B(n_192),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_279),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_294),
.B(n_221),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_257),
.B(n_196),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_282),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_241),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_255),
.A2(n_218),
.B1(n_239),
.B2(n_233),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_284),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_287),
.Y(n_346)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_288),
.A2(n_198),
.B(n_197),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_289),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_268),
.B(n_201),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_336),
.B(n_262),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_334),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_334),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_334),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_300),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_322),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_322),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_300),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_300),
.Y(n_362)
);

AO21x2_ASAP7_75t_L g363 ( 
.A1(n_338),
.A2(n_324),
.B(n_341),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_305),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_314),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_306),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_314),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

CKINVDCx6p67_ASAP7_75t_R g369 ( 
.A(n_311),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_344),
.B(n_262),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_323),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_306),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_350),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_312),
.A2(n_293),
.B1(n_290),
.B2(n_292),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_333),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_310),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_310),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_308),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_335),
.B(n_290),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_332),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_308),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_350),
.B(n_293),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_332),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_338),
.B(n_271),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_315),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_315),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_331),
.Y(n_392)
);

AO22x2_ASAP7_75t_L g393 ( 
.A1(n_325),
.A2(n_291),
.B1(n_297),
.B2(n_281),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_331),
.Y(n_394)
);

AOI21x1_ASAP7_75t_L g395 ( 
.A1(n_307),
.A2(n_267),
.B(n_241),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_318),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_302),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_L g400 ( 
.A(n_320),
.B(n_203),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_303),
.B(n_285),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_340),
.B(n_209),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_340),
.B(n_210),
.Y(n_404)
);

AO21x2_ASAP7_75t_L g405 ( 
.A1(n_327),
.A2(n_215),
.B(n_213),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_325),
.B(n_278),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_302),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_298),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_329),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_313),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_337),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_298),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_299),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_307),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_299),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_345),
.Y(n_417)
);

NAND2xp33_ASAP7_75t_L g418 ( 
.A(n_345),
.B(n_219),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_345),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_380),
.Y(n_420)
);

AND2x2_ASAP7_75t_SL g421 ( 
.A(n_388),
.B(n_323),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_359),
.B(n_349),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g423 ( 
.A(n_406),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_376),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_358),
.B(n_342),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_384),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_309),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_369),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_385),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_369),
.B(n_326),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_401),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_390),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_317),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_390),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_363),
.B(n_309),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_363),
.B(n_309),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_374),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_391),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_375),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_393),
.B(n_317),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_406),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_375),
.B(n_346),
.Y(n_442)
);

INVxp33_ASAP7_75t_SL g443 ( 
.A(n_381),
.Y(n_443)
);

BUFx6f_ASAP7_75t_SL g444 ( 
.A(n_374),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_363),
.B(n_374),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_351),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_374),
.B(n_321),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_357),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_387),
.B(n_323),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_357),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_364),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_366),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_402),
.B(n_329),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_372),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_358),
.B(n_321),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_372),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_377),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_377),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_360),
.B(n_330),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_399),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_360),
.B(n_321),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_399),
.B(n_321),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_393),
.B(n_301),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_378),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_399),
.B(n_329),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_412),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_412),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_413),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_411),
.A2(n_347),
.B(n_328),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_393),
.B(n_304),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_403),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_393),
.B(n_328),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_403),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_407),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_370),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_371),
.B(n_328),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_411),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_407),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_405),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_408),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_407),
.Y(n_484)
);

AND2x2_ASAP7_75t_SL g485 ( 
.A(n_416),
.B(n_347),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_396),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_371),
.B(n_339),
.Y(n_487)
);

AND2x2_ASAP7_75t_SL g488 ( 
.A(n_416),
.B(n_347),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_408),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_387),
.B(n_348),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_421),
.A2(n_400),
.B1(n_404),
.B2(n_405),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_480),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_437),
.B(n_387),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_421),
.B(n_410),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_424),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_487),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_424),
.B(n_387),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_445),
.B(n_387),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_441),
.B(n_410),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_422),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_439),
.A2(n_394),
.B1(n_392),
.B2(n_405),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_486),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_445),
.A2(n_353),
.B1(n_355),
.B2(n_354),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_435),
.A2(n_394),
.B1(n_392),
.B2(n_396),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_423),
.B(n_353),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_423),
.B(n_353),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_435),
.A2(n_397),
.B1(n_398),
.B2(n_307),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_442),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_425),
.B(n_415),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_425),
.B(n_415),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_420),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_481),
.B(n_417),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_481),
.B(n_417),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_428),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_427),
.B(n_343),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_479),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_443),
.B(n_417),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_427),
.B(n_343),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_430),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_465),
.B(n_419),
.Y(n_520)
);

NAND2x1p5_ASAP7_75t_L g521 ( 
.A(n_449),
.B(n_461),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_426),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_436),
.A2(n_397),
.B1(n_398),
.B2(n_419),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_447),
.A2(n_414),
.B(n_354),
.Y(n_524)
);

AO22x1_ASAP7_75t_L g525 ( 
.A1(n_431),
.A2(n_330),
.B1(n_352),
.B2(n_354),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_447),
.B(n_353),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_436),
.B(n_354),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_483),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_456),
.B(n_355),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_456),
.B(n_355),
.Y(n_530)
);

NAND3xp33_ASAP7_75t_SL g531 ( 
.A(n_478),
.B(n_226),
.C(n_224),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_462),
.B(n_355),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_462),
.B(n_356),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_448),
.B(n_450),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_429),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_R g536 ( 
.A(n_444),
.B(n_330),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_477),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_489),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_482),
.A2(n_356),
.B1(n_365),
.B2(n_383),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_444),
.B(n_356),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_473),
.B(n_356),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_475),
.B(n_433),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_482),
.B(n_365),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_460),
.B(n_365),
.Y(n_544)
);

INVx8_ASAP7_75t_L g545 ( 
.A(n_446),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g546 ( 
.A(n_432),
.B(n_352),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_484),
.B(n_383),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_434),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_478),
.B(n_383),
.Y(n_549)
);

NOR2x1p5_ASAP7_75t_L g550 ( 
.A(n_451),
.B(n_383),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_494),
.A2(n_449),
.B1(n_454),
.B2(n_452),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_495),
.B(n_508),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_521),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_545),
.Y(n_554)
);

CKINVDCx11_ASAP7_75t_R g555 ( 
.A(n_514),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_521),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_495),
.B(n_438),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_508),
.B(n_440),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_494),
.A2(n_491),
.B1(n_500),
.B2(n_505),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_499),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_546),
.A2(n_524),
.B(n_529),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_545),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_516),
.B(n_455),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_492),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_500),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_549),
.B(n_464),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_505),
.A2(n_457),
.B1(n_459),
.B2(n_458),
.Y(n_567)
);

NAND3xp33_ASAP7_75t_SL g568 ( 
.A(n_536),
.B(n_540),
.C(n_501),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_545),
.Y(n_569)
);

OR2x4_ASAP7_75t_L g570 ( 
.A(n_531),
.B(n_468),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_541),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_496),
.B(n_519),
.Y(n_572)
);

AND2x2_ASAP7_75t_SL g573 ( 
.A(n_542),
.B(n_485),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_511),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_550),
.B(n_464),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_516),
.B(n_463),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_522),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_515),
.B(n_466),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_506),
.A2(n_474),
.B1(n_476),
.B2(n_488),
.Y(n_579)
);

A2O1A1Ixp33_ASAP7_75t_L g580 ( 
.A1(n_518),
.A2(n_472),
.B(n_469),
.C(n_471),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_506),
.B(n_470),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_528),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_527),
.B(n_382),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_517),
.B(n_382),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_540),
.B(n_382),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_538),
.Y(n_586)
);

NOR3xp33_ASAP7_75t_SL g587 ( 
.A(n_493),
.B(n_231),
.C(n_229),
.Y(n_587)
);

NOR3xp33_ASAP7_75t_L g588 ( 
.A(n_525),
.B(n_534),
.C(n_544),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_535),
.Y(n_589)
);

OAI221xp5_ASAP7_75t_L g590 ( 
.A1(n_501),
.A2(n_490),
.B1(n_379),
.B2(n_361),
.C(n_362),
.Y(n_590)
);

BUFx4_ASAP7_75t_SL g591 ( 
.A(n_548),
.Y(n_591)
);

NOR3xp33_ASAP7_75t_SL g592 ( 
.A(n_543),
.B(n_490),
.C(n_1),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_537),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_502),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_539),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_520),
.B(n_509),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_510),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_504),
.B(n_367),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_503),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_497),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_547),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_512),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_498),
.B(n_368),
.Y(n_603)
);

A2O1A1Ixp33_ASAP7_75t_L g604 ( 
.A1(n_559),
.A2(n_551),
.B(n_567),
.C(n_592),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_560),
.B(n_523),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_560),
.B(n_523),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g607 ( 
.A1(n_561),
.A2(n_532),
.B(n_530),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_559),
.A2(n_533),
.B1(n_513),
.B2(n_526),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_580),
.A2(n_507),
.B(n_453),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_564),
.Y(n_610)
);

OAI222xp33_ASAP7_75t_L g611 ( 
.A1(n_558),
.A2(n_507),
.B1(n_395),
.B2(n_389),
.C1(n_379),
.C2(n_414),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_571),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_578),
.A2(n_583),
.B(n_567),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_566),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_574),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_552),
.B(n_389),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_565),
.B(n_329),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_557),
.B(n_418),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_593),
.B(n_1),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_579),
.A2(n_551),
.B(n_581),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_563),
.B(n_414),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_579),
.A2(n_467),
.B(n_409),
.Y(n_622)
);

OAI221xp5_ASAP7_75t_L g623 ( 
.A1(n_588),
.A2(n_395),
.B1(n_241),
.B2(n_373),
.C(n_409),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_553),
.A2(n_409),
.B(n_373),
.Y(n_624)
);

AO31x2_ASAP7_75t_L g625 ( 
.A1(n_598),
.A2(n_373),
.A3(n_241),
.B(n_87),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_598),
.A2(n_2),
.B(n_3),
.Y(n_626)
);

A2O1A1Ixp33_ASAP7_75t_L g627 ( 
.A1(n_599),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_553),
.A2(n_34),
.B(n_33),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_596),
.B(n_4),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_555),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_589),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_631)
);

OAI21x1_ASAP7_75t_L g632 ( 
.A1(n_603),
.A2(n_602),
.B(n_601),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_576),
.B(n_6),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_589),
.A2(n_7),
.B(n_8),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_597),
.B(n_8),
.Y(n_635)
);

CKINVDCx8_ASAP7_75t_R g636 ( 
.A(n_569),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_554),
.B(n_41),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_SL g638 ( 
.A(n_595),
.B(n_9),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_586),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_572),
.B(n_9),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_571),
.B(n_10),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_582),
.A2(n_43),
.B(n_42),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_577),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_554),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_571),
.B(n_11),
.Y(n_645)
);

AOI21x1_ASAP7_75t_L g646 ( 
.A1(n_600),
.A2(n_46),
.B(n_45),
.Y(n_646)
);

AND3x4_ASAP7_75t_L g647 ( 
.A(n_591),
.B(n_12),
.C(n_13),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_590),
.A2(n_12),
.B(n_13),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_607),
.A2(n_582),
.B(n_594),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_638),
.B(n_562),
.Y(n_650)
);

AO32x2_ASAP7_75t_L g651 ( 
.A1(n_620),
.A2(n_562),
.A3(n_568),
.B1(n_570),
.B2(n_573),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_609),
.A2(n_556),
.B(n_570),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_604),
.A2(n_587),
.B(n_575),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_610),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_613),
.A2(n_575),
.B(n_556),
.Y(n_655)
);

NOR3xp33_ASAP7_75t_SL g656 ( 
.A(n_631),
.B(n_14),
.C(n_16),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_620),
.A2(n_556),
.B(n_585),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_648),
.A2(n_584),
.B(n_16),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_622),
.A2(n_14),
.B(n_17),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_621),
.A2(n_18),
.B(n_19),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_615),
.Y(n_661)
);

AO31x2_ASAP7_75t_L g662 ( 
.A1(n_643),
.A2(n_107),
.A3(n_181),
.B(n_180),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_612),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_639),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_644),
.Y(n_665)
);

AO22x2_ASAP7_75t_L g666 ( 
.A1(n_605),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_612),
.B(n_20),
.Y(n_667)
);

BUFx6f_ASAP7_75t_SL g668 ( 
.A(n_630),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_612),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_636),
.Y(n_670)
);

BUFx12f_ASAP7_75t_L g671 ( 
.A(n_630),
.Y(n_671)
);

AOI221x1_ASAP7_75t_L g672 ( 
.A1(n_627),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.C(n_24),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_626),
.A2(n_618),
.B(n_634),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_626),
.A2(n_22),
.B(n_24),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_623),
.A2(n_27),
.B(n_28),
.Y(n_675)
);

NOR2x1_ASAP7_75t_L g676 ( 
.A(n_633),
.B(n_27),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_638),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_634),
.A2(n_608),
.B(n_616),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_608),
.A2(n_29),
.B(n_30),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_606),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_611),
.A2(n_182),
.B(n_47),
.Y(n_681)
);

O2A1O1Ixp33_ASAP7_75t_SL g682 ( 
.A1(n_640),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_637),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_619),
.B(n_179),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_642),
.A2(n_617),
.B(n_628),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_629),
.B(n_52),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_635),
.B(n_178),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_641),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_645),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_632),
.A2(n_54),
.B(n_57),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_625),
.B(n_58),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_625),
.Y(n_692)
);

AO32x2_ASAP7_75t_L g693 ( 
.A1(n_625),
.A2(n_59),
.A3(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_647),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_646),
.B(n_624),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_613),
.A2(n_67),
.B(n_68),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_614),
.B(n_69),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_604),
.B(n_71),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_636),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_614),
.B(n_74),
.Y(n_700)
);

BUFx2_ASAP7_75t_SL g701 ( 
.A(n_699),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_679),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_670),
.Y(n_703)
);

CKINVDCx6p67_ASAP7_75t_R g704 ( 
.A(n_668),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_654),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_669),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_683),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_665),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_670),
.Y(n_709)
);

INVx6_ASAP7_75t_L g710 ( 
.A(n_663),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_653),
.A2(n_84),
.B1(n_86),
.B2(n_89),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_663),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_671),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_666),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_650),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_666),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_688),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_689),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_661),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_680),
.B(n_99),
.Y(n_720)
);

BUFx4f_ASAP7_75t_L g721 ( 
.A(n_697),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_664),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_678),
.B(n_177),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_658),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_667),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_649),
.Y(n_726)
);

BUFx6f_ASAP7_75t_SL g727 ( 
.A(n_697),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_700),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_SL g729 ( 
.A1(n_673),
.A2(n_674),
.B1(n_700),
.B2(n_692),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_677),
.A2(n_105),
.B1(n_110),
.B2(n_111),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_672),
.A2(n_113),
.B1(n_114),
.B2(n_116),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_SL g732 ( 
.A1(n_691),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_732)
);

BUFx12f_ASAP7_75t_L g733 ( 
.A(n_695),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_SL g734 ( 
.A1(n_681),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_734)
);

BUFx8_ASAP7_75t_L g735 ( 
.A(n_651),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_651),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_693),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_656),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_652),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_676),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_662),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_698),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_662),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_684),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_662),
.Y(n_745)
);

BUFx12f_ASAP7_75t_L g746 ( 
.A(n_695),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_693),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_657),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_655),
.B(n_176),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_705),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_733),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_746),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_719),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_722),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_726),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_737),
.B(n_693),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_739),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_706),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_748),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_741),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_747),
.B(n_659),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_721),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_743),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_708),
.Y(n_764)
);

AO21x2_ASAP7_75t_L g765 ( 
.A1(n_745),
.A2(n_685),
.B(n_690),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_702),
.A2(n_694),
.B1(n_660),
.B2(n_687),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_731),
.A2(n_675),
.B1(n_686),
.B2(n_696),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_708),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_707),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_707),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_736),
.Y(n_771)
);

OAI21x1_ASAP7_75t_L g772 ( 
.A1(n_723),
.A2(n_682),
.B(n_143),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_717),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_718),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_720),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_702),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_721),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_720),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_740),
.Y(n_779)
);

AOI222xp33_ASAP7_75t_L g780 ( 
.A1(n_735),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.C1(n_154),
.C2(n_156),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_725),
.B(n_158),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_735),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_712),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_749),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_750),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_755),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_SL g787 ( 
.A(n_777),
.B(n_704),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_773),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_750),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_753),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_755),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_777),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_753),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_758),
.B(n_744),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_760),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_755),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_764),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_755),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_758),
.B(n_728),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_756),
.B(n_729),
.Y(n_800)
);

NOR2x1_ASAP7_75t_SL g801 ( 
.A(n_777),
.B(n_701),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_768),
.Y(n_802)
);

AO21x2_ASAP7_75t_L g803 ( 
.A1(n_765),
.A2(n_731),
.B(n_738),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_757),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_779),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_775),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_756),
.B(n_729),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_771),
.B(n_712),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_760),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_763),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_765),
.A2(n_738),
.B(n_711),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_759),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_771),
.B(n_712),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_812),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_797),
.B(n_802),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_805),
.B(n_773),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_812),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_812),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_795),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_SL g820 ( 
.A(n_794),
.B(n_751),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_804),
.Y(n_821)
);

AO21x2_ASAP7_75t_L g822 ( 
.A1(n_803),
.A2(n_811),
.B(n_775),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_794),
.B(n_774),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_786),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_795),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_800),
.A2(n_780),
.B1(n_766),
.B2(n_727),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_809),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_809),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_806),
.B(n_778),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_810),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_786),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_800),
.B(n_774),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_807),
.B(n_783),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_807),
.B(n_783),
.Y(n_834)
);

NOR2x1_ASAP7_75t_R g835 ( 
.A(n_792),
.B(n_709),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_824),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_815),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_817),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_816),
.B(n_788),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_815),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_816),
.B(n_788),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_827),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_829),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_827),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_822),
.B(n_799),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_824),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_822),
.B(n_785),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_817),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_833),
.B(n_808),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_834),
.B(n_813),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_843),
.B(n_837),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_840),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_844),
.B(n_822),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_849),
.B(n_821),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_849),
.B(n_823),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_842),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_850),
.B(n_823),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_842),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_838),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_850),
.B(n_839),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_855),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_856),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_860),
.B(n_839),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_851),
.B(n_845),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_852),
.B(n_845),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_853),
.A2(n_826),
.B(n_820),
.C(n_847),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_858),
.B(n_830),
.Y(n_867)
);

NOR2x1_ASAP7_75t_L g868 ( 
.A(n_862),
.B(n_713),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_861),
.B(n_863),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_865),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_864),
.B(n_860),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_867),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_870),
.B(n_855),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_868),
.B(n_871),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_869),
.B(n_857),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_872),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_870),
.A2(n_866),
.B1(n_803),
.B2(n_811),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_868),
.B(n_854),
.Y(n_878)
);

INVx3_ASAP7_75t_SL g879 ( 
.A(n_868),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_872),
.Y(n_880)
);

AOI321xp33_ASAP7_75t_L g881 ( 
.A1(n_877),
.A2(n_716),
.A3(n_714),
.B1(n_767),
.B2(n_859),
.C(n_724),
.Y(n_881)
);

NOR3xp33_ASAP7_75t_L g882 ( 
.A(n_874),
.B(n_703),
.C(n_859),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_SL g883 ( 
.A1(n_878),
.A2(n_854),
.B(n_751),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_879),
.Y(n_884)
);

NOR2xp67_ASAP7_75t_L g885 ( 
.A(n_873),
.B(n_875),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_876),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_884),
.A2(n_803),
.B1(n_876),
.B2(n_880),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_882),
.A2(n_811),
.B1(n_787),
.B2(n_715),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_885),
.A2(n_767),
.B(n_776),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_883),
.B(n_841),
.Y(n_890)
);

OAI31xp33_ASAP7_75t_L g891 ( 
.A1(n_886),
.A2(n_730),
.A3(n_832),
.B(n_724),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_881),
.B(n_836),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_890),
.Y(n_893)
);

AOI221xp5_ASAP7_75t_L g894 ( 
.A1(n_887),
.A2(n_778),
.B1(n_730),
.B2(n_848),
.C(n_761),
.Y(n_894)
);

AOI322xp5_ASAP7_75t_L g895 ( 
.A1(n_892),
.A2(n_761),
.A3(n_782),
.B1(n_784),
.B2(n_734),
.C1(n_817),
.C2(n_846),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_889),
.B(n_836),
.Y(n_896)
);

NAND4xp25_ASAP7_75t_L g897 ( 
.A(n_888),
.B(n_792),
.C(n_751),
.D(n_752),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_896),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_893),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_895),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_897),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_894),
.B(n_891),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_896),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_896),
.Y(n_904)
);

NOR3x1_ASAP7_75t_L g905 ( 
.A(n_904),
.B(n_799),
.C(n_835),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_899),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_899),
.B(n_846),
.Y(n_907)
);

NAND3xp33_ASAP7_75t_L g908 ( 
.A(n_898),
.B(n_732),
.C(n_734),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_903),
.Y(n_909)
);

OA22x2_ASAP7_75t_L g910 ( 
.A1(n_901),
.A2(n_752),
.B1(n_792),
.B2(n_831),
.Y(n_910)
);

NOR3x1_ASAP7_75t_L g911 ( 
.A(n_902),
.B(n_835),
.C(n_781),
.Y(n_911)
);

NOR2x1p5_ASAP7_75t_L g912 ( 
.A(n_909),
.B(n_900),
.Y(n_912)
);

NOR2x1_ASAP7_75t_L g913 ( 
.A(n_906),
.B(n_752),
.Y(n_913)
);

OAI211xp5_ASAP7_75t_L g914 ( 
.A1(n_907),
.A2(n_792),
.B(n_752),
.C(n_742),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_911),
.Y(n_915)
);

AND4x1_ASAP7_75t_L g916 ( 
.A(n_913),
.B(n_905),
.C(n_908),
.D(n_910),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_915),
.B(n_831),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_SL g918 ( 
.A(n_912),
.B(n_777),
.C(n_818),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_915),
.B(n_710),
.Y(n_919)
);

NOR5xp2_ASAP7_75t_L g920 ( 
.A(n_914),
.B(n_790),
.C(n_789),
.D(n_785),
.E(n_793),
.Y(n_920)
);

OAI211xp5_ASAP7_75t_L g921 ( 
.A1(n_918),
.A2(n_828),
.B(n_825),
.C(n_819),
.Y(n_921)
);

NAND4xp75_ASAP7_75t_L g922 ( 
.A(n_919),
.B(n_814),
.C(n_819),
.D(n_789),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_917),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_916),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_920),
.Y(n_925)
);

NAND3x1_ASAP7_75t_L g926 ( 
.A(n_916),
.B(n_804),
.C(n_769),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_924),
.B(n_925),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_923),
.B(n_754),
.Y(n_928)
);

AND3x1_ASAP7_75t_L g929 ( 
.A(n_926),
.B(n_770),
.C(n_769),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_922),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_921),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_924),
.Y(n_932)
);

XNOR2xp5_ASAP7_75t_L g933 ( 
.A(n_924),
.B(n_782),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_924),
.B(n_801),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_924),
.Y(n_935)
);

NAND2x1_ASAP7_75t_SL g936 ( 
.A(n_932),
.B(n_798),
.Y(n_936)
);

AO22x2_ASAP7_75t_L g937 ( 
.A1(n_935),
.A2(n_927),
.B1(n_930),
.B2(n_934),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_933),
.B(n_798),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_928),
.Y(n_939)
);

AOI222xp33_ASAP7_75t_SL g940 ( 
.A1(n_931),
.A2(n_798),
.B1(n_796),
.B2(n_791),
.C1(n_786),
.C2(n_757),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_SL g941 ( 
.A1(n_929),
.A2(n_762),
.B1(n_757),
.B2(n_791),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_936),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_937),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_939),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_938),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_941),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_943),
.A2(n_940),
.B(n_772),
.Y(n_947)
);

OAI22x1_ASAP7_75t_SL g948 ( 
.A1(n_942),
.A2(n_757),
.B1(n_159),
.B2(n_160),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_944),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_949),
.A2(n_946),
.B(n_945),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_950),
.Y(n_951)
);

INVxp67_ASAP7_75t_SL g952 ( 
.A(n_951),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_952),
.A2(n_947),
.B1(n_948),
.B2(n_762),
.Y(n_953)
);

OAI22xp33_ASAP7_75t_L g954 ( 
.A1(n_952),
.A2(n_762),
.B1(n_796),
.B2(n_791),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_953),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_954),
.A2(n_161),
.B(n_163),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_955),
.A2(n_164),
.B(n_165),
.Y(n_957)
);

AOI21xp33_ASAP7_75t_SL g958 ( 
.A1(n_956),
.A2(n_168),
.B(n_169),
.Y(n_958)
);

AO22x2_ASAP7_75t_L g959 ( 
.A1(n_957),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_959)
);

AOI211xp5_ASAP7_75t_L g960 ( 
.A1(n_959),
.A2(n_958),
.B(n_174),
.C(n_175),
.Y(n_960)
);


endmodule