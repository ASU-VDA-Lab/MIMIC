module fake_jpeg_3339_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_48),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx2_ASAP7_75t_SL g69 ( 
.A(n_54),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_23),
.B(n_9),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_60),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_61),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_63),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_28),
.Y(n_91)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_65),
.B(n_0),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_28),
.B1(n_37),
.B2(n_19),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_66),
.A2(n_86),
.B(n_100),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_17),
.B1(n_21),
.B2(n_31),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_71),
.B1(n_103),
.B2(n_109),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_17),
.B1(n_21),
.B2(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_73),
.B(n_81),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_32),
.B1(n_26),
.B2(n_37),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_10),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_29),
.B1(n_22),
.B2(n_34),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_99),
.B1(n_5),
.B2(n_9),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_34),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_84),
.B(n_93),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_28),
.B1(n_33),
.B2(n_18),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_33),
.C(n_26),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_15),
.C(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_92),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_108),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_38),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_98),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_24),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_29),
.B1(n_18),
.B2(n_31),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_41),
.A2(n_31),
.B1(n_21),
.B2(n_18),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_44),
.A2(n_30),
.B(n_31),
.C(n_18),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_102),
.B(n_104),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_41),
.A2(n_18),
.B1(n_30),
.B2(n_3),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_44),
.B(n_10),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_50),
.A2(n_18),
.B1(n_30),
.B2(n_3),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_106),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_41),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_110),
.B(n_112),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_116),
.A2(n_126),
.B1(n_130),
.B2(n_71),
.Y(n_172)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_135),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_67),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_92),
.B1(n_94),
.B2(n_108),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_131),
.B(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_91),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_138),
.Y(n_160)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_96),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_136),
.B(n_144),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_95),
.C(n_70),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_15),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_142),
.B(n_146),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_96),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_105),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_86),
.B(n_15),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_101),
.B(n_78),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_147),
.A2(n_113),
.B(n_135),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_70),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_148),
.B(n_151),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_88),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_156),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_95),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_154),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_85),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_126),
.C(n_140),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_157),
.B(n_181),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_105),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_171),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_123),
.B1(n_145),
.B2(n_127),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_128),
.B1(n_125),
.B2(n_97),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_165),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_106),
.B1(n_89),
.B2(n_77),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_112),
.B1(n_132),
.B2(n_138),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_169),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_86),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_172),
.B(n_116),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_74),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_97),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_114),
.B(n_82),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_89),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_74),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_110),
.B(n_77),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_117),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_175),
.A2(n_146),
.B1(n_142),
.B2(n_122),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_183),
.A2(n_190),
.B(n_192),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_158),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_195),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_185),
.B(n_180),
.Y(n_230)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_150),
.A2(n_129),
.B1(n_144),
.B2(n_136),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_191),
.A2(n_209),
.B1(n_212),
.B2(n_207),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_139),
.Y(n_192)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_124),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_196),
.B(n_208),
.Y(n_225)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_210),
.B(n_192),
.Y(n_239)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_180),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_152),
.B1(n_174),
.B2(n_156),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_203),
.A2(n_179),
.B1(n_174),
.B2(n_165),
.Y(n_220)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_205),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_214),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_207),
.A2(n_202),
.B1(n_194),
.B2(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_148),
.B(n_75),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_75),
.B1(n_111),
.B2(n_97),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_147),
.A2(n_97),
.B(n_173),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_154),
.B(n_157),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_211),
.B(n_213),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_168),
.A2(n_179),
.B1(n_159),
.B2(n_174),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_166),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_223),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_149),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_222),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_179),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_149),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_224),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_167),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_227),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_183),
.A2(n_153),
.B1(n_163),
.B2(n_170),
.Y(n_227)
);

A2O1A1O1Ixp25_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_153),
.B(n_180),
.C(n_164),
.D(n_176),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_229),
.B(n_232),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_231),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_163),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_164),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_210),
.B(n_199),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_193),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_245),
.C(n_259),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_212),
.B1(n_188),
.B2(n_185),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_256),
.B1(n_225),
.B2(n_223),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_193),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_255),
.Y(n_264)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_191),
.B(n_203),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_230),
.A2(n_188),
.B1(n_208),
.B2(n_209),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_198),
.C(n_197),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_225),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_258),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_217),
.A3(n_216),
.B1(n_228),
.B2(n_221),
.C1(n_236),
.C2(n_226),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_263),
.B(n_242),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_236),
.C(n_216),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_272),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_218),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_249),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_247),
.A2(n_217),
.B1(n_222),
.B2(n_238),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_254),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_227),
.B1(n_218),
.B2(n_224),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_255),
.A2(n_190),
.B1(n_219),
.B2(n_229),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_231),
.C(n_219),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_246),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_276),
.A2(n_258),
.B1(n_261),
.B2(n_273),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_257),
.B(n_253),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_278),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_284),
.B1(n_272),
.B2(n_243),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_244),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_283),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_257),
.B1(n_251),
.B2(n_256),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_284),
.A2(n_270),
.B1(n_251),
.B2(n_269),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_294),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_SL g290 ( 
.A(n_281),
.B(n_274),
.C(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_293),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_262),
.C(n_260),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_289),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_277),
.B(n_276),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_282),
.B(n_288),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_292),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_295),
.A2(n_287),
.B(n_293),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_301),
.C(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_306),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_299),
.B(n_300),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_299),
.Y(n_310)
);


endmodule