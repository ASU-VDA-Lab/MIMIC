module fake_jpeg_500_n_619 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_619);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_619;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx6f_ASAP7_75t_SL g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_58),
.Y(n_163)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g133 ( 
.A(n_63),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_68),
.B(n_110),
.Y(n_149)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_70),
.Y(n_168)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_71),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_72),
.B(n_116),
.Y(n_145)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_76),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_77),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_48),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_80),
.B(n_101),
.Y(n_210)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_81),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_82),
.Y(n_200)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_85),
.Y(n_205)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_87),
.Y(n_207)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_90),
.Y(n_223)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_50),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_93),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_94),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_97),
.Y(n_222)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_99),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_42),
.B(n_3),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_54),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_103),
.A2(n_32),
.B1(n_37),
.B2(n_49),
.Y(n_174)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_24),
.B(n_18),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_118),
.Y(n_146)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_47),
.B(n_3),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_120),
.Y(n_217)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_17),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_122),
.B(n_3),
.Y(n_186)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_123),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_44),
.Y(n_125)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_125),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_44),
.Y(n_126)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_126),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_44),
.Y(n_128)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_47),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_129),
.B(n_157),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_70),
.A2(n_54),
.B1(n_28),
.B2(n_38),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_131),
.A2(n_153),
.B1(n_171),
.B2(n_198),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_63),
.A2(n_54),
.B1(n_53),
.B2(n_28),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_132),
.A2(n_131),
.B1(n_171),
.B2(n_170),
.Y(n_240)
);

NAND2x1_ASAP7_75t_L g147 ( 
.A(n_80),
.B(n_21),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_L g287 ( 
.A(n_147),
.B(n_10),
.C(n_11),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_76),
.A2(n_128),
.B1(n_127),
.B2(n_126),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_56),
.B(n_55),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_154),
.B(n_13),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_64),
.B(n_55),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_91),
.B(n_29),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_160),
.B(n_166),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_64),
.B(n_29),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_77),
.A2(n_20),
.B1(n_52),
.B2(n_49),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_60),
.B(n_32),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_172),
.B(n_175),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_174),
.A2(n_216),
.B1(n_20),
.B2(n_34),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_61),
.B(n_37),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_57),
.B(n_19),
.C(n_52),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_213),
.C(n_33),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_84),
.B(n_16),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_185),
.B(n_193),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_186),
.B(n_203),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_107),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_71),
.A2(n_19),
.B(n_52),
.Y(n_195)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_195),
.B(n_15),
.CI(n_13),
.CON(n_302),
.SN(n_302)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_58),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_197),
.B(n_204),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_66),
.A2(n_19),
.B1(n_49),
.B2(n_45),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_82),
.B(n_45),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_86),
.B(n_45),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_88),
.B(n_39),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_209),
.B(n_211),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_94),
.B(n_39),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_85),
.B(n_39),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_212),
.B(n_12),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_78),
.B(n_38),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_119),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_87),
.A2(n_53),
.B1(n_38),
.B2(n_34),
.Y(n_216)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_224),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_226),
.A2(n_241),
.B1(n_267),
.B2(n_282),
.Y(n_307)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_156),
.Y(n_227)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_227),
.Y(n_311)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_228),
.Y(n_346)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_230),
.Y(n_320)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_158),
.Y(n_232)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_232),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_153),
.A2(n_108),
.B1(n_100),
.B2(n_99),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_233),
.A2(n_245),
.B1(n_253),
.B2(n_263),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_147),
.B(n_78),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_235),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_236),
.B(n_258),
.Y(n_325)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_136),
.Y(n_238)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_238),
.Y(n_322)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_159),
.Y(n_239)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_239),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_240),
.A2(n_244),
.B1(n_303),
.B2(n_151),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_182),
.A2(n_125),
.B1(n_97),
.B2(n_95),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_162),
.Y(n_242)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_242),
.Y(n_339)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_141),
.Y(n_243)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

INVx11_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_173),
.A2(n_34),
.B1(n_33),
.B2(n_28),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_150),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_246),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_133),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_247),
.B(n_248),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_133),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_144),
.Y(n_249)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_249),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_164),
.B(n_33),
.C(n_21),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_250),
.B(n_161),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_137),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_252),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_184),
.A2(n_21),
.B1(n_20),
.B2(n_5),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_143),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_254),
.B(n_281),
.Y(n_306)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_255),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_143),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_256),
.B(n_295),
.Y(n_323)
);

BUFx2_ASAP7_75t_SL g257 ( 
.A(n_167),
.Y(n_257)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_257),
.Y(n_330)
);

OA22x2_ASAP7_75t_L g258 ( 
.A1(n_132),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_258)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_150),
.Y(n_259)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_259),
.Y(n_335)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_261),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_188),
.Y(n_262)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_262),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_210),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_263)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_265),
.Y(n_338)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_183),
.Y(n_266)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_266),
.Y(n_341)
);

AOI22x1_ASAP7_75t_L g267 ( 
.A1(n_146),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_188),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_268),
.B(n_287),
.Y(n_328)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_135),
.Y(n_269)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_269),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_191),
.Y(n_270)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_270),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_163),
.Y(n_271)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_178),
.Y(n_272)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_272),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_196),
.Y(n_273)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_273),
.Y(n_350)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_148),
.Y(n_275)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_179),
.Y(n_276)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_276),
.Y(n_359)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_278),
.Y(n_358)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_136),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_280),
.Y(n_316)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_152),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_142),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_194),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_163),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_283),
.B(n_284),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_165),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_130),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_286),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_167),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_139),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_288),
.B(n_289),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_165),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_217),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_290),
.B(n_297),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_291),
.B(n_292),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_213),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_187),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_293),
.B(n_294),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_149),
.B(n_12),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_140),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_152),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_177),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_298),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_L g361 ( 
.A(n_299),
.B(n_302),
.Y(n_361)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_168),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_300),
.B(n_301),
.Y(n_344)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_168),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_138),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_145),
.B(n_15),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_304),
.A2(n_305),
.B(n_140),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_201),
.B(n_206),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_310),
.B(n_225),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_235),
.A2(n_221),
.B1(n_220),
.B2(n_207),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_312),
.A2(n_314),
.B1(n_254),
.B2(n_286),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_296),
.A2(n_241),
.B1(n_237),
.B2(n_292),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_233),
.A2(n_219),
.B1(n_214),
.B2(n_190),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_324),
.A2(n_327),
.B1(n_348),
.B2(n_259),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_240),
.A2(n_219),
.B1(n_189),
.B2(n_205),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_277),
.A2(n_146),
.B(n_176),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_333),
.B(n_301),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_264),
.A2(n_169),
.B1(n_222),
.B2(n_223),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_334),
.A2(n_222),
.B1(n_332),
.B2(n_312),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_342),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_251),
.A2(n_151),
.B1(n_176),
.B2(n_161),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_357),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_253),
.A2(n_200),
.B1(n_189),
.B2(n_190),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_234),
.A2(n_274),
.B1(n_302),
.B2(n_240),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_155),
.Y(n_402)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_363),
.Y(n_364)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_364),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_327),
.A2(n_267),
.B1(n_282),
.B2(n_304),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_365),
.A2(n_378),
.B1(n_382),
.B2(n_398),
.Y(n_415)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_353),
.Y(n_366)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_366),
.Y(n_412)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_316),
.Y(n_367)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_367),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_350),
.Y(n_368)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_368),
.Y(n_437)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_377),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_287),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_371),
.B(n_373),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_325),
.A2(n_258),
.B(n_298),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_372),
.A2(n_407),
.B(n_345),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_245),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_307),
.A2(n_272),
.B1(n_231),
.B2(n_229),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_375),
.A2(n_390),
.B1(n_395),
.B2(n_408),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_230),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_376),
.B(n_391),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_306),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_347),
.B(n_224),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_379),
.B(n_399),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_383),
.Y(n_418)
);

FAx1_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_258),
.CI(n_303),
.CON(n_381),
.SN(n_381)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_381),
.B(n_344),
.Y(n_417)
);

OAI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_318),
.A2(n_297),
.B1(n_271),
.B2(n_283),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_331),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_331),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_384),
.B(n_387),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_268),
.C(n_262),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_385),
.B(n_402),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_314),
.A2(n_355),
.B1(n_353),
.B2(n_346),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_386),
.Y(n_438)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_328),
.A2(n_244),
.B(n_223),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_388),
.A2(n_396),
.B(n_330),
.Y(n_423)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_354),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_389),
.B(n_393),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_318),
.A2(n_200),
.B1(n_205),
.B2(n_284),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_335),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_346),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_405),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_324),
.A2(n_246),
.B1(n_289),
.B2(n_178),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_328),
.A2(n_155),
.B(n_270),
.Y(n_396)
);

NOR2x1_ASAP7_75t_L g397 ( 
.A(n_328),
.B(n_252),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_397),
.Y(n_441)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_311),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_R g420 ( 
.A(n_400),
.B(n_406),
.Y(n_420)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_313),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_401),
.B(n_403),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_343),
.B(n_300),
.Y(n_403)
);

BUFx24_ASAP7_75t_L g404 ( 
.A(n_321),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_404),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_315),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_352),
.B(n_207),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_351),
.A2(n_322),
.B1(n_320),
.B2(n_335),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_319),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_409),
.Y(n_414)
);

OAI21xp33_ASAP7_75t_SL g449 ( 
.A1(n_413),
.A2(n_423),
.B(n_447),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_381),
.A2(n_361),
.B1(n_344),
.B2(n_309),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_416),
.A2(n_419),
.B1(n_439),
.B2(n_441),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_417),
.A2(n_426),
.B(n_428),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_381),
.A2(n_344),
.B1(n_322),
.B2(n_317),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_424),
.A2(n_439),
.B1(n_365),
.B2(n_406),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_329),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_425),
.B(n_442),
.C(n_385),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_392),
.A2(n_319),
.B(n_330),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_374),
.A2(n_336),
.B(n_320),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_427),
.A2(n_388),
.B(n_396),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_392),
.A2(n_336),
.B(n_358),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_377),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_431),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_380),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_383),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_392),
.A2(n_358),
.B(n_359),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_381),
.A2(n_390),
.B1(n_373),
.B2(n_364),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_402),
.B(n_338),
.Y(n_442)
);

OAI32xp33_ASAP7_75t_L g445 ( 
.A1(n_367),
.A2(n_341),
.A3(n_313),
.B1(n_356),
.B2(n_337),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_445),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_372),
.A2(n_337),
.B(n_339),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_411),
.B(n_405),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_448),
.B(n_451),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_425),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_369),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_411),
.B(n_371),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_452),
.B(n_459),
.Y(n_505)
);

A2O1A1Ixp33_ASAP7_75t_SL g453 ( 
.A1(n_417),
.A2(n_374),
.B(n_376),
.C(n_397),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_453),
.A2(n_447),
.B(n_413),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_454),
.A2(n_468),
.B1(n_479),
.B2(n_410),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_457),
.A2(n_423),
.B(n_427),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_387),
.Y(n_459)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_424),
.A2(n_378),
.B1(n_407),
.B2(n_384),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_461),
.A2(n_464),
.B1(n_440),
.B2(n_444),
.Y(n_513)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_436),
.Y(n_462)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_462),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_419),
.B(n_389),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_463),
.B(n_470),
.Y(n_488)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_465),
.Y(n_514)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_430),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_467),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_430),
.B(n_409),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_416),
.A2(n_395),
.B1(n_394),
.B2(n_391),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_421),
.B(n_404),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_437),
.Y(n_471)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_471),
.Y(n_499)
);

BUFx5_ASAP7_75t_L g472 ( 
.A(n_437),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_472),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_421),
.B(n_401),
.C(n_399),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_432),
.C(n_433),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_435),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_474),
.Y(n_494)
);

INVxp33_ASAP7_75t_L g475 ( 
.A(n_435),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_475),
.B(n_476),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_422),
.B(n_393),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_445),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_477),
.B(n_480),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_421),
.B(n_404),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_442),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_415),
.A2(n_391),
.B1(n_404),
.B2(n_366),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_422),
.B(n_339),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_410),
.B(n_326),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_481),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_440),
.B(n_340),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_482),
.Y(n_508)
);

XOR2x2_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_425),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_484),
.B(n_497),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_491),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_492),
.B(n_493),
.C(n_498),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_473),
.B(n_418),
.C(n_446),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_454),
.A2(n_415),
.B1(n_417),
.B2(n_446),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_495),
.A2(n_500),
.B1(n_461),
.B2(n_458),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_478),
.B(n_418),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_450),
.B(n_429),
.C(n_426),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_501),
.A2(n_506),
.B(n_512),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_463),
.B(n_443),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_502),
.B(n_503),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_466),
.B(n_443),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_460),
.B(n_429),
.C(n_428),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_504),
.B(n_475),
.C(n_456),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_455),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_509),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_467),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_510),
.A2(n_513),
.B1(n_458),
.B2(n_468),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_469),
.A2(n_438),
.B(n_420),
.Y(n_512)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_487),
.Y(n_515)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_515),
.Y(n_557)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_487),
.Y(n_516)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_516),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_502),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_518),
.B(n_521),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_494),
.B(n_465),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_514),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_522),
.B(n_524),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_523),
.A2(n_535),
.B1(n_511),
.B2(n_504),
.Y(n_544)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_514),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_483),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_525),
.A2(n_533),
.B1(n_537),
.B2(n_540),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_526),
.B(n_538),
.Y(n_555)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_507),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_527),
.B(n_530),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_486),
.B(n_456),
.C(n_469),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_528),
.B(n_532),
.C(n_492),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_529),
.A2(n_495),
.B1(n_511),
.B2(n_506),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_501),
.A2(n_457),
.B(n_453),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_498),
.B(n_476),
.C(n_449),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_507),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_513),
.A2(n_479),
.B1(n_420),
.B2(n_482),
.Y(n_535)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_485),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_493),
.B(n_453),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_485),
.B(n_489),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_539),
.Y(n_552)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_489),
.Y(n_540)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_531),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_541),
.B(n_559),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_532),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_542),
.B(n_545),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_544),
.A2(n_526),
.B1(n_539),
.B2(n_538),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_517),
.B(n_488),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_546),
.A2(n_515),
.B1(n_537),
.B2(n_540),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_519),
.B(n_497),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_547),
.B(n_519),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_528),
.B(n_488),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_550),
.B(n_551),
.C(n_560),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_484),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_523),
.A2(n_490),
.B1(n_505),
.B2(n_496),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_553),
.B(n_554),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_536),
.B(n_512),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_520),
.B(n_491),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_561),
.A2(n_573),
.B1(n_414),
.B2(n_551),
.Y(n_578)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_556),
.Y(n_562)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_562),
.Y(n_583)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_549),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_564),
.A2(n_575),
.B1(n_483),
.B2(n_412),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_548),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_565),
.B(n_412),
.Y(n_585)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_543),
.Y(n_566)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_566),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_567),
.A2(n_542),
.B1(n_550),
.B2(n_545),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_552),
.A2(n_557),
.B1(n_558),
.B2(n_521),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_568),
.A2(n_569),
.B1(n_499),
.B2(n_480),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_559),
.A2(n_508),
.B1(n_503),
.B2(n_530),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_555),
.A2(n_534),
.B(n_453),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_570),
.A2(n_577),
.B(n_569),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_572),
.B(n_340),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_554),
.A2(n_534),
.B1(n_453),
.B2(n_525),
.Y(n_573)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_555),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_547),
.A2(n_414),
.B(n_520),
.Y(n_577)
);

XNOR2x1_ASAP7_75t_L g593 ( 
.A(n_578),
.B(n_580),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_579),
.B(n_582),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_581),
.B(n_590),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_568),
.A2(n_560),
.B1(n_499),
.B2(n_444),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_584),
.B(n_586),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_585),
.A2(n_574),
.B(n_563),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_573),
.B(n_360),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_567),
.B(n_360),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_588),
.B(n_589),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_566),
.A2(n_412),
.B1(n_308),
.B2(n_472),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_565),
.B(n_308),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_591),
.B(n_561),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_583),
.B(n_562),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_594),
.B(n_597),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_598),
.B(n_599),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_587),
.B(n_575),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_585),
.B(n_576),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_601),
.B(n_578),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_595),
.B(n_588),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_602),
.B(n_606),
.C(n_607),
.Y(n_609)
);

AND2x2_ASAP7_75t_SL g612 ( 
.A(n_604),
.B(n_589),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_592),
.B(n_580),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_593),
.B(n_596),
.Y(n_607)
);

NOR2x1_ASAP7_75t_L g608 ( 
.A(n_593),
.B(n_586),
.Y(n_608)
);

AOI21x1_ASAP7_75t_L g610 ( 
.A1(n_608),
.A2(n_581),
.B(n_570),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_610),
.A2(n_612),
.B(n_608),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_603),
.A2(n_577),
.B(n_600),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_611),
.A2(n_605),
.B(n_572),
.Y(n_614)
);

AO21x1_ASAP7_75t_L g615 ( 
.A1(n_613),
.A2(n_614),
.B(n_609),
.Y(n_615)
);

AOI31xp33_ASAP7_75t_L g616 ( 
.A1(n_615),
.A2(n_576),
.A3(n_595),
.B(n_602),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_616),
.A2(n_571),
.B(n_590),
.Y(n_617)
);

O2A1O1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_617),
.A2(n_571),
.B(n_326),
.C(n_356),
.Y(n_618)
);

BUFx24_ASAP7_75t_SL g619 ( 
.A(n_618),
.Y(n_619)
);


endmodule