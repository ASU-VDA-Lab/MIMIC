module real_jpeg_7140_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_1),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_2),
.A2(n_45),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_2),
.A2(n_45),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_2),
.A2(n_45),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_3),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_3),
.A2(n_92),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_3),
.A2(n_92),
.B1(n_180),
.B2(n_183),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_3),
.B(n_25),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_3),
.A2(n_331),
.B(n_333),
.C(n_339),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_3),
.B(n_71),
.C(n_174),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_3),
.B(n_148),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_3),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_3),
.B(n_75),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_4),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_4),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_4),
.A2(n_233),
.B1(n_249),
.B2(n_252),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_4),
.A2(n_233),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_4),
.A2(n_233),
.B1(n_367),
.B2(n_369),
.Y(n_366)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_5),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_6),
.Y(n_176)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_6),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_6),
.Y(n_384)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_7),
.Y(n_260)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_9),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_10),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_11),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_11),
.A2(n_27),
.B1(n_41),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_11),
.A2(n_41),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_11),
.A2(n_41),
.B1(n_174),
.B2(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_12),
.Y(n_430)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_426),
.B(n_428),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_200),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_199),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_149),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_19),
.B(n_149),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_140),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_132),
.B2(n_133),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_60),
.B1(n_61),
.B2(n_131),
.Y(n_22)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_23),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_35),
.B(n_42),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_24),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_25),
.B(n_43),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_25),
.B(n_136),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_25),
.B(n_231),
.Y(n_243)
);

AO22x1_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_30),
.B2(n_32),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g262 ( 
.A(n_26),
.B(n_123),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_27),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_29),
.Y(n_111)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_29),
.Y(n_115)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_29),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_29),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_37),
.A2(n_92),
.B(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g256 ( 
.A1(n_40),
.A2(n_257),
.A3(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_42),
.B(n_243),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_49),
.B(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_49),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_49),
.B(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_56),
.B2(n_58),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_94),
.B1(n_95),
.B2(n_130),
.Y(n_61)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_62),
.A2(n_130),
.B1(n_141),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_62),
.A2(n_130),
.B1(n_245),
.B2(n_253),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_62),
.B(n_242),
.C(n_245),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_85),
.B(n_86),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_63),
.A2(n_188),
.B(n_194),
.Y(n_187)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_64),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_64),
.B(n_87),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_64),
.B(n_345),
.Y(n_344)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_75),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_68),
.Y(n_346)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_69),
.Y(n_338)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_73),
.Y(n_190)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_75),
.B(n_160),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_75),
.B(n_345),
.Y(n_361)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_81),
.B2(n_83),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_78),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_79),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_82),
.Y(n_174)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_82),
.Y(n_370)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_85),
.B(n_86),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_85),
.A2(n_159),
.B(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_92),
.B(n_138),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g333 ( 
.A1(n_92),
.A2(n_334),
.B(n_336),
.Y(n_333)
);

INVx4_ASAP7_75t_SL g193 ( 
.A(n_93),
.Y(n_193)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_116),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_96),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_108),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_100),
.Y(n_335)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_104),
.Y(n_349)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_109),
.B(n_142),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_109),
.A2(n_142),
.B(n_148),
.Y(n_301)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_110),
.Y(n_252)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_111),
.Y(n_251)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_116),
.A2(n_143),
.B(n_148),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_116),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_124),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_120),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_129),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_133),
.C(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_133),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_134),
.B(n_230),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_135),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_137),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_138),
.Y(n_234)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B(n_146),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_142),
.B(n_248),
.Y(n_271)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_147),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_147),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_148),
.B(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.C(n_167),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_150),
.A2(n_154),
.B1(n_155),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_155),
.A2(n_156),
.B(n_166),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_166),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_157),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_159),
.B(n_361),
.Y(n_405)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_195),
.B(n_196),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_169),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_187),
.Y(n_169)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_195),
.B1(n_196),
.B2(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_170),
.A2(n_187),
.B1(n_195),
.B2(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_170),
.B(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_170),
.A2(n_195),
.B1(n_330),
.B2(n_408),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_177),
.B(n_179),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_171),
.B(n_179),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_171),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_171),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_217),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_183),
.Y(n_265)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_187),
.Y(n_313)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g285 ( 
.A(n_194),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_194),
.B(n_344),
.Y(n_372)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_235),
.B(n_425),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_202),
.B(n_205),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.C(n_212),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_206),
.A2(n_210),
.B1(n_211),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_206),
.Y(n_317)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_212),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_226),
.C(n_228),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_213),
.A2(n_214),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_225),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_215),
.B(n_225),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_216),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_218),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_219),
.A2(n_264),
.B(n_266),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx8_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_224),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_226),
.B(n_228),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_227),
.B(n_247),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_417),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_306),
.C(n_320),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_293),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_279),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_240),
.B(n_279),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_254),
.C(n_269),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_241),
.B(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_254),
.A2(n_255),
.B1(n_269),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_263),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_256),
.B(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_276),
.B(n_284),
.Y(n_283)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_268),
.Y(n_392)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_269),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.C(n_274),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_274),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_275),
.B(n_382),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_276),
.B(n_365),
.Y(n_395)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_287),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_282),
.C(n_287),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_285),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_286),
.B(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_290),
.C(n_291),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_293),
.A2(n_420),
.B(n_421),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_305),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_294),
.B(n_305),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_302),
.C(n_303),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_318),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_307),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_315),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_308),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_308),
.B(n_319),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_308),
.B(n_315),
.Y(n_424)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_312),
.CI(n_314),
.CON(n_308),
.SN(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_318),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_350),
.B(n_416),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_322),
.B(n_325),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.C(n_341),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_326),
.B(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_329),
.A2(n_341),
.B1(n_342),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_329),
.Y(n_413)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

INVx8_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_338),
.Y(n_358)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_410),
.B(n_415),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_400),
.B(n_409),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_376),
.B(n_399),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_362),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_362),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_360),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_355),
.A2(n_356),
.B1(n_360),
.B2(n_379),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_360),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_371),
.Y(n_362)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_363),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_383),
.Y(n_382)
);

INVx6_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx6_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_373),
.B1(n_374),
.B2(n_375),
.Y(n_371)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_372),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_373),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_374),
.C(n_402),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_385),
.B(n_398),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_380),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_380),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_394),
.B(n_397),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_393),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_395),
.B(n_396),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_403),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_401),
.B(n_403),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_407),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_406),
.C(n_407),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_414),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_411),
.B(n_414),
.Y(n_415)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_419),
.B(n_422),
.C(n_423),
.D(n_424),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_426),
.Y(n_429)
);

INVx13_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);


endmodule