module fake_jpeg_3608_n_431 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_431);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_431;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_54),
.B(n_58),
.Y(n_132)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g165 ( 
.A(n_55),
.Y(n_165)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_16),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_59),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_60),
.Y(n_176)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_27),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_64),
.B(n_72),
.Y(n_120)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_16),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_73),
.B(n_85),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

INVx2_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_105),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_77),
.B(n_78),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_12),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_79),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_33),
.B(n_0),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_86),
.Y(n_177)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_87),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_19),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_93),
.Y(n_173)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_25),
.B(n_0),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_97),
.Y(n_142)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_100),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_26),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_106),
.Y(n_144)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_43),
.B(n_8),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_107),
.B(n_111),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_26),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_109),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_26),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_38),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_112),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_113),
.B(n_89),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_69),
.A2(n_38),
.B1(n_47),
.B2(n_50),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_115),
.A2(n_116),
.B1(n_122),
.B2(n_127),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_47),
.B1(n_42),
.B2(n_50),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_62),
.A2(n_51),
.B1(n_49),
.B2(n_47),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_117),
.A2(n_150),
.B1(n_157),
.B2(n_158),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_83),
.B1(n_79),
.B2(n_99),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_65),
.A2(n_36),
.B1(n_40),
.B2(n_46),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g190 ( 
.A(n_124),
.B(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_76),
.B(n_40),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_125),
.B(n_162),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_61),
.A2(n_49),
.B1(n_36),
.B2(n_46),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_34),
.B1(n_44),
.B2(n_42),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_131),
.A2(n_143),
.B1(n_175),
.B2(n_157),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_86),
.A2(n_44),
.B1(n_34),
.B2(n_43),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_SL g149 ( 
.A1(n_96),
.A2(n_29),
.B(n_39),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_149),
.A2(n_138),
.B(n_150),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_105),
.A2(n_49),
.B1(n_29),
.B2(n_39),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_35),
.B1(n_53),
.B2(n_4),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_170),
.B1(n_178),
.B2(n_185),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_71),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_80),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_92),
.B(n_2),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_66),
.B(n_2),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_182),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_112),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_102),
.A2(n_7),
.B1(n_8),
.B2(n_81),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_93),
.A2(n_7),
.B1(n_8),
.B2(n_104),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_90),
.A2(n_59),
.B1(n_67),
.B2(n_82),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_66),
.B(n_89),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_138),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_59),
.B(n_55),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_165),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_97),
.A2(n_60),
.B1(n_74),
.B2(n_58),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_186),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_97),
.B1(n_115),
.B2(n_163),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_187),
.A2(n_229),
.B1(n_193),
.B2(n_234),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_165),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_188),
.B(n_201),
.Y(n_254)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_189),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_191),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_194),
.A2(n_199),
.B(n_236),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_142),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_195),
.B(n_205),
.Y(n_260)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_196),
.Y(n_259)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_200),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_144),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_203),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_120),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_204),
.B(n_214),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_148),
.B(n_146),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_128),
.B(n_132),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_206),
.B(n_210),
.Y(n_272)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_135),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_140),
.B(n_147),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_145),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_165),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_215),
.Y(n_256)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_121),
.B(n_136),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_118),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_143),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_217),
.B(n_219),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_118),
.B(n_156),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_218),
.B(n_223),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_131),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_220),
.B(n_226),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_156),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_221),
.Y(n_274)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_167),
.B(n_133),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_227),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_126),
.B(n_141),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_225),
.B(n_237),
.Y(n_291)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_152),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_230),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_126),
.A2(n_116),
.B1(n_155),
.B2(n_135),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_167),
.B(n_129),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_129),
.B(n_152),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_231),
.B(n_235),
.Y(n_277)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_232),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_117),
.B(n_158),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_234),
.C(n_198),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_153),
.B(n_178),
.C(n_175),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_153),
.B(n_134),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_114),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_141),
.B(n_173),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_134),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_240),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_222),
.B1(n_193),
.B2(n_229),
.Y(n_257)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVx13_ASAP7_75t_L g247 ( 
.A(n_241),
.Y(n_247)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_138),
.B(n_76),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_243),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_142),
.B(n_160),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_246),
.B1(n_243),
.B2(n_245),
.Y(n_263)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_154),
.Y(n_245)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_142),
.B(n_160),
.Y(n_246)
);

OAI32xp33_ASAP7_75t_L g248 ( 
.A1(n_206),
.A2(n_195),
.A3(n_217),
.B1(n_194),
.B2(n_219),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_248),
.B(n_269),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_249),
.A2(n_276),
.B1(n_270),
.B2(n_286),
.Y(n_323)
);

AND2x6_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_194),
.Y(n_250)
);

BUFx12_ASAP7_75t_L g313 ( 
.A(n_250),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_205),
.B(n_216),
.CI(n_192),
.CON(n_253),
.SN(n_253)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_263),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_257),
.A2(n_290),
.B1(n_249),
.B2(n_274),
.Y(n_303)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_197),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_233),
.A2(n_225),
.B1(n_239),
.B2(n_198),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_271),
.A2(n_282),
.B1(n_257),
.B2(n_291),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g279 ( 
.A(n_190),
.B(n_243),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_264),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_221),
.A2(n_198),
.B1(n_226),
.B2(n_236),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_237),
.A2(n_210),
.B1(n_220),
.B2(n_190),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_198),
.B(n_240),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_293),
.A2(n_297),
.B(n_318),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_252),
.B(n_186),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_294),
.B(n_309),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_221),
.C(n_203),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_295),
.B(n_296),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_221),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_242),
.B(n_208),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_213),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_304),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g300 ( 
.A(n_260),
.B(n_241),
.C(n_207),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_316),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_191),
.C(n_232),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_301),
.B(n_308),
.Y(n_342)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_255),
.Y(n_302)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_303),
.A2(n_305),
.B1(n_307),
.B2(n_312),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_275),
.A2(n_248),
.B1(n_274),
.B2(n_280),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_275),
.A2(n_250),
.B1(n_279),
.B2(n_277),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_264),
.B(n_260),
.C(n_268),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_252),
.B(n_283),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_266),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_319),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_311),
.B(n_314),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_273),
.A2(n_255),
.B1(n_259),
.B2(n_261),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_259),
.B(n_261),
.C(n_283),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_288),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_288),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_321),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_256),
.A2(n_284),
.B(n_288),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_253),
.B(n_273),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_253),
.B(n_278),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_325),
.Y(n_334)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_251),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_278),
.A2(n_270),
.B(n_254),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_258),
.B(n_265),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_281),
.B(n_287),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_285),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_281),
.B(n_251),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_322),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_328),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_325),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_293),
.A2(n_286),
.B(n_287),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_330),
.A2(n_333),
.B(n_337),
.Y(n_357)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_307),
.B(n_258),
.CI(n_265),
.CON(n_335),
.SN(n_335)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_335),
.B(n_336),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g336 ( 
.A(n_326),
.B(n_267),
.CI(n_247),
.CON(n_336),
.SN(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_304),
.A2(n_247),
.B(n_285),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_352),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_315),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_312),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_306),
.A2(n_276),
.B(n_247),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_346),
.A2(n_349),
.B(n_301),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_305),
.A2(n_276),
.B1(n_297),
.B2(n_326),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_347),
.A2(n_303),
.B1(n_329),
.B2(n_349),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_306),
.A2(n_326),
.B(n_317),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_299),
.B(n_319),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_308),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_362),
.C(n_368),
.Y(n_375)
);

OAI321xp33_ASAP7_75t_L g355 ( 
.A1(n_352),
.A2(n_332),
.A3(n_334),
.B1(n_331),
.B2(n_320),
.C(n_329),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_355),
.A2(n_356),
.B1(n_358),
.B2(n_370),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_347),
.A2(n_296),
.B1(n_292),
.B2(n_295),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_341),
.Y(n_360)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_360),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_314),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_361),
.B(n_365),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_318),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_350),
.A2(n_313),
.B1(n_316),
.B2(n_310),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_364),
.A2(n_347),
.B1(n_331),
.B2(n_349),
.Y(n_377)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_321),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_367),
.Y(n_382)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_343),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_313),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_339),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_344),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_338),
.A2(n_298),
.B1(n_302),
.B2(n_313),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_371),
.A2(n_329),
.B(n_330),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_372),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_373),
.A2(n_363),
.B(n_330),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_353),
.B(n_332),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_376),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_362),
.B(n_342),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_359),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_356),
.A2(n_350),
.B1(n_338),
.B2(n_348),
.Y(n_381)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_381),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_342),
.C(n_351),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_375),
.C(n_376),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_385),
.Y(n_397)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_350),
.Y(n_386)
);

OAI21xp33_ASAP7_75t_L g390 ( 
.A1(n_386),
.A2(n_387),
.B(n_364),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_361),
.B(n_334),
.Y(n_387)
);

NAND2x1_ASAP7_75t_SL g389 ( 
.A(n_383),
.B(n_357),
.Y(n_389)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_389),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_394),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_373),
.A2(n_357),
.B(n_371),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_395),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_382),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_393),
.A2(n_400),
.B1(n_363),
.B2(n_327),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_346),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_396),
.B(n_375),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_380),
.B(n_359),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_398),
.B(n_401),
.Y(n_409)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_388),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_383),
.B(n_369),
.Y(n_401)
);

FAx1_ASAP7_75t_SL g402 ( 
.A(n_392),
.B(n_355),
.CI(n_384),
.CON(n_402),
.SN(n_402)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_402),
.B(n_407),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_397),
.Y(n_404)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_404),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_397),
.A2(n_379),
.B1(n_378),
.B2(n_381),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_405),
.A2(n_412),
.B1(n_377),
.B2(n_400),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_406),
.B(n_411),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_391),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_396),
.B(n_351),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_414),
.A2(n_403),
.B1(n_354),
.B2(n_402),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_409),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_408),
.A2(n_395),
.B1(n_354),
.B2(n_389),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_386),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_410),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_420),
.A2(n_423),
.B1(n_417),
.B2(n_402),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_387),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_421),
.B(n_374),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_422),
.A2(n_415),
.B1(n_418),
.B2(n_419),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_416),
.A2(n_403),
.B1(n_372),
.B2(n_389),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_425),
.C(n_426),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_427),
.Y(n_428)
);

CKINVDCx14_ASAP7_75t_R g429 ( 
.A(n_428),
.Y(n_429)
);

OAI21xp33_ASAP7_75t_SL g430 ( 
.A1(n_429),
.A2(n_425),
.B(n_399),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_399),
.Y(n_431)
);


endmodule