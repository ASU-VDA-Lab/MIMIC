module fake_ariane_601_n_1052 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1052);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1052;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_913;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_183;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_515;
wire n_379;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_958;
wire n_945;
wire n_207;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_779;
wire n_731;
wire n_903;
wire n_315;
wire n_871;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_928;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1045;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_612;
wire n_333;
wire n_449;
wire n_388;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_998;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_1044;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_124),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_18),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_65),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_18),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_38),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_44),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_168),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_160),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_69),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_48),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_145),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_100),
.Y(n_196)
);

BUFx8_ASAP7_75t_SL g197 ( 
.A(n_143),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_9),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_63),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_117),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_29),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_64),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_87),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_32),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_68),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_139),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_135),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_0),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_33),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_119),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_159),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_57),
.Y(n_219)
);

CKINVDCx12_ASAP7_75t_R g220 ( 
.A(n_45),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_23),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_6),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_130),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_114),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_111),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_169),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_54),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_115),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_155),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_179),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_131),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_137),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_138),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_83),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_36),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_80),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_104),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_12),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_14),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_144),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_15),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_73),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_60),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_150),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_116),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_51),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_108),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_89),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_161),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_17),
.Y(n_251)
);

INVxp33_ASAP7_75t_SL g252 ( 
.A(n_185),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

INVxp33_ASAP7_75t_SL g255 ( 
.A(n_181),
.Y(n_255)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_240),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_186),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_191),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_202),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_251),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_214),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_234),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_182),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_197),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_247),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_250),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_199),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_228),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_204),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_198),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_207),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_213),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_200),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_220),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_221),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_239),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_183),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_242),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_232),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_235),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_236),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_184),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_241),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_246),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_225),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_252),
.A2(n_195),
.B1(n_206),
.B2(n_187),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_245),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_270),
.A2(n_216),
.B1(n_248),
.B2(n_243),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_262),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_227),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_288),
.A2(n_249),
.B1(n_238),
.B2(n_233),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_278),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_189),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_267),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_227),
.Y(n_317)
);

BUFx8_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_256),
.B(n_266),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_276),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

AND2x6_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_227),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_270),
.A2(n_231),
.B1(n_230),
.B2(n_229),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_190),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_289),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_259),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_271),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_279),
.B(n_192),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_292),
.B(n_193),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_272),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_277),
.A2(n_268),
.B1(n_260),
.B2(n_255),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_281),
.B(n_196),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_201),
.Y(n_343)
);

OAI21x1_ASAP7_75t_L g344 ( 
.A1(n_284),
.A2(n_298),
.B(n_290),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_253),
.B(n_227),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_263),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_263),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_278),
.A2(n_226),
.B1(n_224),
.B2(n_223),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_258),
.B(n_203),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_264),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_259),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_277),
.B(n_205),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_297),
.B(n_208),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_313),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_316),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_330),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_305),
.Y(n_363)
);

AOI21x1_ASAP7_75t_L g364 ( 
.A1(n_307),
.A2(n_188),
.B(n_257),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_351),
.B(n_260),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_307),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_305),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_317),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_310),
.B(n_268),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_308),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_305),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_308),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_309),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_351),
.B(n_287),
.Y(n_374)
);

CKINVDCx6p67_ASAP7_75t_R g375 ( 
.A(n_332),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_309),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_301),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_301),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_301),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_351),
.B(n_275),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_301),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_351),
.B(n_280),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_301),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_314),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_314),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_317),
.B(n_280),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

NOR2x1p5_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_210),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_319),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

INVxp33_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_312),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_324),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_312),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_348),
.B(n_211),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_302),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_351),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_322),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_322),
.Y(n_403)
);

AND3x2_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_0),
.C(n_1),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_327),
.B(n_212),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_323),
.Y(n_407)
);

NOR3xp33_ASAP7_75t_L g408 ( 
.A(n_303),
.B(n_218),
.C(n_215),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_323),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_325),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_325),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_334),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_333),
.B(n_188),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_339),
.Y(n_415)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_354),
.B(n_1),
.C(n_2),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_333),
.B(n_353),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_339),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_320),
.B(n_188),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_342),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_310),
.B(n_188),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_342),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_335),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_354),
.B(n_2),
.C(n_3),
.Y(n_425)
);

NOR2x1p5_ASAP7_75t_L g426 ( 
.A(n_353),
.B(n_3),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_346),
.B(n_4),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_349),
.B(n_188),
.Y(n_429)
);

AND2x2_ASAP7_75t_SL g430 ( 
.A(n_399),
.B(n_408),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_373),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_373),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_406),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_406),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_424),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_366),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g438 ( 
.A(n_392),
.B(n_340),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_377),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_367),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_367),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_371),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_371),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_400),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_385),
.B(n_311),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_357),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_386),
.B(n_346),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_410),
.Y(n_450)
);

OR2x6_ASAP7_75t_L g451 ( 
.A(n_387),
.B(n_355),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_369),
.B(n_338),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_395),
.B(n_355),
.Y(n_453)
);

BUFx2_ASAP7_75t_R g454 ( 
.A(n_374),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_375),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_R g457 ( 
.A(n_387),
.B(n_347),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_357),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_375),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_415),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_377),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_366),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_405),
.B(n_347),
.Y(n_466)
);

XNOR2x2_ASAP7_75t_L g467 ( 
.A(n_416),
.B(n_306),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_420),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_420),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_419),
.B(n_310),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_382),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_403),
.Y(n_472)
);

XOR2x2_ASAP7_75t_L g473 ( 
.A(n_383),
.B(n_326),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_368),
.B(n_352),
.Y(n_474)
);

NOR2xp67_ASAP7_75t_L g475 ( 
.A(n_401),
.B(n_350),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_366),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_403),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_365),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_427),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_380),
.B(n_349),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_418),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_405),
.B(n_350),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_419),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_418),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_368),
.B(n_320),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_422),
.Y(n_486)
);

NAND2x1p5_ASAP7_75t_L g487 ( 
.A(n_397),
.B(n_330),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_390),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_422),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_423),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_423),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_407),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_370),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_370),
.B(n_304),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_407),
.Y(n_496)
);

NOR2xp67_ASAP7_75t_L g497 ( 
.A(n_401),
.B(n_315),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_382),
.A2(n_341),
.B(n_336),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_357),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_409),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

BUFx8_ASAP7_75t_L g502 ( 
.A(n_427),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_409),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_411),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_404),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_426),
.B(n_349),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_411),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_417),
.B(n_429),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_377),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_370),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_360),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_463),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_470),
.B(n_372),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_431),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_470),
.B(n_483),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_449),
.B(n_337),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_432),
.B(n_372),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_433),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_474),
.B(n_318),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_457),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_452),
.B(n_304),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_506),
.B(n_390),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_434),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_448),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_459),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_490),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_491),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_452),
.B(n_304),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_474),
.B(n_402),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_430),
.A2(n_426),
.B1(n_329),
.B2(n_402),
.Y(n_533)
);

NOR3xp33_ASAP7_75t_L g534 ( 
.A(n_438),
.B(n_425),
.C(n_343),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_453),
.B(n_318),
.Y(n_535)
);

A2O1A1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_509),
.A2(n_376),
.B(n_372),
.C(n_402),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_485),
.B(n_402),
.Y(n_537)
);

NOR2xp67_ASAP7_75t_L g538 ( 
.A(n_456),
.B(n_421),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_466),
.B(n_412),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_430),
.B(n_330),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_473),
.A2(n_414),
.B1(n_389),
.B2(n_393),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_451),
.B(n_318),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_451),
.A2(n_412),
.B1(n_356),
.B2(n_362),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_457),
.A2(n_389),
.B1(n_393),
.B2(n_376),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_445),
.B(n_376),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_446),
.B(n_356),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_463),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_440),
.B(n_397),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_482),
.B(n_362),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_459),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_451),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_499),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_499),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_L g554 ( 
.A(n_488),
.B(n_391),
.Y(n_554)
);

AND2x6_ASAP7_75t_SL g555 ( 
.A(n_447),
.B(n_345),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_463),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_436),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_479),
.B(n_345),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_502),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_502),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_461),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_479),
.B(n_345),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_494),
.B(n_463),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_439),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_494),
.B(n_358),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_461),
.B(n_397),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_440),
.B(n_397),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_441),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_497),
.B(n_358),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_475),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_467),
.A2(n_360),
.B1(n_361),
.B2(n_331),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_442),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_450),
.B(n_360),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_443),
.B(n_361),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_455),
.B(n_361),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_510),
.B(n_509),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_471),
.A2(n_391),
.B1(n_393),
.B2(n_389),
.Y(n_577)
);

AND2x6_ASAP7_75t_SL g578 ( 
.A(n_458),
.B(n_4),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_510),
.B(n_331),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_510),
.B(n_331),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_518),
.B(n_480),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_526),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_527),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_523),
.B(n_460),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_567),
.Y(n_585)
);

NOR3xp33_ASAP7_75t_SL g586 ( 
.A(n_521),
.B(n_498),
.C(n_444),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_558),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_562),
.B(n_505),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_567),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_566),
.B(n_478),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_529),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_R g592 ( 
.A(n_566),
.B(n_559),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_530),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_563),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_547),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_R g596 ( 
.A(n_560),
.B(n_478),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_563),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_531),
.B(n_524),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_522),
.B(n_462),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_517),
.B(n_464),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_516),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_561),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_520),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_577),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_542),
.B(n_454),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_528),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_555),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_L g608 ( 
.A(n_535),
.B(n_435),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_SL g609 ( 
.A(n_534),
.B(n_498),
.C(n_469),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_547),
.Y(n_610)
);

AOI22x1_ASAP7_75t_L g611 ( 
.A1(n_557),
.A2(n_471),
.B1(n_435),
.B2(n_465),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_525),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_547),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_563),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_517),
.B(n_454),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_564),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_551),
.B(n_468),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_568),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_539),
.A2(n_476),
.B1(n_493),
.B2(n_511),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_549),
.B(n_437),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_524),
.B(n_572),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_SL g622 ( 
.A(n_577),
.B(n_495),
.C(n_492),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_554),
.A2(n_510),
.B1(n_331),
.B2(n_393),
.Y(n_623)
);

BUFx2_ASAP7_75t_SL g624 ( 
.A(n_538),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_532),
.B(n_513),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_541),
.B(n_331),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_514),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_515),
.B(n_513),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_580),
.Y(n_629)
);

AND3x1_ASAP7_75t_SL g630 ( 
.A(n_578),
.B(n_5),
.C(n_6),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_537),
.B(n_472),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_550),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_548),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_570),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_580),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_R g636 ( 
.A(n_514),
.B(n_364),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_515),
.B(n_477),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_556),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_552),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_533),
.B(n_487),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_556),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_543),
.B(n_481),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_580),
.B(n_424),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_546),
.A2(n_512),
.B1(n_508),
.B2(n_507),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_611),
.A2(n_519),
.B(n_574),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_596),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_582),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_591),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_602),
.Y(n_649)
);

OAI22x1_ASAP7_75t_L g650 ( 
.A1(n_615),
.A2(n_581),
.B1(n_590),
.B2(n_598),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_587),
.B(n_546),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_586),
.B(n_544),
.Y(n_652)
);

AO31x2_ASAP7_75t_L g653 ( 
.A1(n_628),
.A2(n_536),
.A3(n_625),
.B(n_637),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_593),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_600),
.B(n_545),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_644),
.A2(n_519),
.B(n_545),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_584),
.B(n_565),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_583),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_621),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_588),
.B(n_540),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_626),
.A2(n_574),
.B(n_576),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_609),
.A2(n_575),
.B(n_573),
.Y(n_662)
);

AOI21x1_ASAP7_75t_L g663 ( 
.A1(n_640),
.A2(n_364),
.B(n_579),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_601),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_644),
.A2(n_569),
.B(n_548),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_603),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_615),
.B(n_389),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_612),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_604),
.B(n_553),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_604),
.A2(n_500),
.B(n_496),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_609),
.A2(n_571),
.B(n_503),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_620),
.A2(n_504),
.B(n_501),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_586),
.A2(n_384),
.B(n_381),
.C(n_378),
.Y(n_673)
);

O2A1O1Ixp5_ASAP7_75t_L g674 ( 
.A1(n_627),
.A2(n_424),
.B(n_428),
.C(n_378),
.Y(n_674)
);

A2O1A1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_622),
.A2(n_384),
.B(n_381),
.C(n_378),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_596),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_633),
.A2(n_486),
.B(n_484),
.Y(n_677)
);

AND2x6_ASAP7_75t_L g678 ( 
.A(n_614),
.B(n_489),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_622),
.A2(n_424),
.B1(n_428),
.B2(n_388),
.Y(n_679)
);

AOI21x1_ASAP7_75t_L g680 ( 
.A1(n_594),
.A2(n_384),
.B(n_381),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_643),
.A2(n_487),
.B(n_359),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_617),
.B(n_428),
.Y(n_682)
);

OAI21x1_ASAP7_75t_L g683 ( 
.A1(n_633),
.A2(n_396),
.B(n_388),
.Y(n_683)
);

NAND2x1p5_ASAP7_75t_L g684 ( 
.A(n_629),
.B(n_428),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_634),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_L g686 ( 
.A1(n_619),
.A2(n_396),
.B(n_388),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_617),
.A2(n_396),
.B(n_398),
.C(n_379),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_643),
.A2(n_398),
.B(n_379),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_629),
.A2(n_394),
.B(n_35),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_619),
.A2(n_324),
.B(n_394),
.Y(n_690)
);

AO21x1_ASAP7_75t_L g691 ( 
.A1(n_599),
.A2(n_188),
.B(n_324),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_623),
.A2(n_37),
.B(n_34),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_605),
.B(n_616),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_610),
.A2(n_631),
.B(n_606),
.Y(n_694)
);

INVx5_ASAP7_75t_L g695 ( 
.A(n_635),
.Y(n_695)
);

AOI21xp33_ASAP7_75t_L g696 ( 
.A1(n_642),
.A2(n_597),
.B(n_594),
.Y(n_696)
);

AOI21x1_ASAP7_75t_L g697 ( 
.A1(n_597),
.A2(n_324),
.B(n_394),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_624),
.B(n_614),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_618),
.A2(n_639),
.B(n_632),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_610),
.Y(n_700)
);

AOI21x1_ASAP7_75t_SL g701 ( 
.A1(n_630),
.A2(n_638),
.B(n_627),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_585),
.A2(n_40),
.B(n_39),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_635),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_608),
.B(n_592),
.Y(n_704)
);

OAI22x1_ASAP7_75t_L g705 ( 
.A1(n_693),
.A2(n_630),
.B1(n_607),
.B2(n_629),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_698),
.B(n_614),
.Y(n_706)
);

O2A1O1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_652),
.A2(n_585),
.B(n_589),
.C(n_592),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_651),
.B(n_589),
.Y(n_708)
);

AO31x2_ASAP7_75t_L g709 ( 
.A1(n_691),
.A2(n_641),
.A3(n_638),
.B(n_595),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_656),
.A2(n_629),
.B(n_641),
.Y(n_710)
);

NAND3x1_ASAP7_75t_L g711 ( 
.A(n_667),
.B(n_5),
.C(n_7),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_L g712 ( 
.A(n_676),
.B(n_613),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_645),
.A2(n_636),
.B(n_635),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_655),
.A2(n_613),
.B(n_635),
.Y(n_714)
);

O2A1O1Ixp33_ASAP7_75t_SL g715 ( 
.A1(n_682),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_663),
.A2(n_636),
.B(n_613),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_665),
.A2(n_613),
.B(n_595),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_675),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_657),
.A2(n_614),
.B(n_394),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_650),
.A2(n_324),
.B1(n_394),
.B2(n_12),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_657),
.A2(n_394),
.B(n_10),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_659),
.B(n_11),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_SL g723 ( 
.A1(n_673),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_685),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_671),
.A2(n_13),
.B(n_16),
.Y(n_725)
);

OR2x6_ASAP7_75t_L g726 ( 
.A(n_698),
.B(n_41),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_661),
.A2(n_43),
.B(n_42),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_646),
.A2(n_649),
.B1(n_669),
.B2(n_704),
.Y(n_728)
);

AO31x2_ASAP7_75t_L g729 ( 
.A1(n_670),
.A2(n_121),
.A3(n_177),
.B(n_176),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_669),
.A2(n_690),
.B(n_671),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_662),
.A2(n_674),
.B(n_679),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_648),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_695),
.B(n_16),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_660),
.B(n_654),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_695),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_664),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_666),
.B(n_19),
.Y(n_737)
);

AO31x2_ASAP7_75t_L g738 ( 
.A1(n_672),
.A2(n_679),
.A3(n_687),
.B(n_647),
.Y(n_738)
);

AO31x2_ASAP7_75t_L g739 ( 
.A1(n_658),
.A2(n_120),
.A3(n_175),
.B(n_173),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_668),
.B(n_19),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_678),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_699),
.B(n_695),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_700),
.Y(n_743)
);

O2A1O1Ixp33_ASAP7_75t_SL g744 ( 
.A1(n_701),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_699),
.B(n_23),
.Y(n_745)
);

OAI22x1_ASAP7_75t_L g746 ( 
.A1(n_703),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_690),
.A2(n_681),
.B(n_686),
.Y(n_747)
);

AO31x2_ASAP7_75t_L g748 ( 
.A1(n_689),
.A2(n_126),
.A3(n_172),
.B(n_167),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_696),
.B(n_24),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_678),
.B(n_25),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_696),
.B(n_26),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_694),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_678),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_684),
.A2(n_688),
.B1(n_686),
.B2(n_680),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_684),
.B(n_27),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_692),
.A2(n_27),
.B(n_28),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_702),
.A2(n_28),
.B(n_29),
.Y(n_757)
);

O2A1O1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_653),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_758)
);

AO31x2_ASAP7_75t_L g759 ( 
.A1(n_653),
.A2(n_129),
.A3(n_165),
.B(n_46),
.Y(n_759)
);

OAI21x1_ASAP7_75t_L g760 ( 
.A1(n_683),
.A2(n_132),
.B(n_163),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_678),
.B(n_30),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_677),
.B(n_31),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_653),
.A2(n_47),
.B(n_49),
.C(n_50),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_697),
.B(n_52),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_667),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_645),
.A2(n_58),
.B(n_59),
.Y(n_766)
);

AOI31xp67_ASAP7_75t_L g767 ( 
.A1(n_652),
.A2(n_61),
.A3(n_62),
.B(n_66),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_667),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_648),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_656),
.A2(n_178),
.B(n_74),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_656),
.A2(n_162),
.B(n_75),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_743),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_732),
.Y(n_773)
);

CKINVDCx6p67_ASAP7_75t_R g774 ( 
.A(n_705),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_734),
.B(n_72),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_725),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_724),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_SL g778 ( 
.A1(n_761),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_722),
.Y(n_779)
);

INVx4_ASAP7_75t_SL g780 ( 
.A(n_726),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_735),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_736),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_SL g783 ( 
.A1(n_741),
.A2(n_85),
.B(n_86),
.Y(n_783)
);

CKINVDCx6p67_ASAP7_75t_R g784 ( 
.A(n_726),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_742),
.Y(n_785)
);

CKINVDCx11_ASAP7_75t_R g786 ( 
.A(n_753),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_755),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_728),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_753),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_769),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_737),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_751),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_708),
.Y(n_793)
);

CKINVDCx11_ASAP7_75t_R g794 ( 
.A(n_706),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_749),
.Y(n_795)
);

INVx6_ASAP7_75t_L g796 ( 
.A(n_706),
.Y(n_796)
);

INVx6_ASAP7_75t_L g797 ( 
.A(n_712),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_711),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_798)
);

INVx4_ASAP7_75t_L g799 ( 
.A(n_752),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_740),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_716),
.Y(n_801)
);

OAI22xp33_ASAP7_75t_L g802 ( 
.A1(n_750),
.A2(n_720),
.B1(n_768),
.B2(n_765),
.Y(n_802)
);

INVx3_ASAP7_75t_SL g803 ( 
.A(n_733),
.Y(n_803)
);

CKINVDCx6p67_ASAP7_75t_R g804 ( 
.A(n_746),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_745),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_709),
.Y(n_806)
);

BUFx10_ASAP7_75t_L g807 ( 
.A(n_762),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_713),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_730),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_SL g810 ( 
.A1(n_770),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_714),
.Y(n_811)
);

BUFx4f_ASAP7_75t_SL g812 ( 
.A(n_764),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_758),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_759),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_739),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_719),
.Y(n_816)
);

CKINVDCx11_ASAP7_75t_R g817 ( 
.A(n_754),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_715),
.A2(n_106),
.B1(n_107),
.B2(n_110),
.Y(n_818)
);

CKINVDCx8_ASAP7_75t_R g819 ( 
.A(n_707),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_717),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_721),
.A2(n_112),
.B1(n_113),
.B2(n_118),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_710),
.B(n_125),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_739),
.Y(n_823)
);

CKINVDCx11_ASAP7_75t_R g824 ( 
.A(n_744),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_727),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_747),
.B(n_127),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_738),
.Y(n_827)
);

BUFx12f_ASAP7_75t_L g828 ( 
.A(n_723),
.Y(n_828)
);

CKINVDCx8_ASAP7_75t_R g829 ( 
.A(n_767),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_772),
.Y(n_830)
);

NAND2x1p5_ASAP7_75t_L g831 ( 
.A(n_820),
.B(n_766),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_773),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_782),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_790),
.Y(n_834)
);

OR2x6_ASAP7_75t_L g835 ( 
.A(n_815),
.B(n_823),
.Y(n_835)
);

BUFx2_ASAP7_75t_R g836 ( 
.A(n_777),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_814),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_779),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_799),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_801),
.A2(n_731),
.B(n_771),
.Y(n_840)
);

INVxp67_ASAP7_75t_R g841 ( 
.A(n_809),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_785),
.B(n_738),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_806),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_795),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_801),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_793),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_827),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_793),
.B(n_763),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_800),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_808),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_808),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_820),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_826),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_811),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_791),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_813),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_783),
.A2(n_718),
.B(n_757),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_781),
.B(n_128),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_789),
.Y(n_859)
);

AOI21x1_ASAP7_75t_L g860 ( 
.A1(n_822),
.A2(n_809),
.B(n_756),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_788),
.B(n_709),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_807),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_804),
.A2(n_760),
.B1(n_729),
.B2(n_748),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_807),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_825),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_825),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_825),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_787),
.B(n_729),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_797),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_787),
.B(n_748),
.Y(n_870)
);

AOI21x1_ASAP7_75t_L g871 ( 
.A1(n_798),
.A2(n_133),
.B(n_136),
.Y(n_871)
);

AO21x1_ASAP7_75t_SL g872 ( 
.A1(n_853),
.A2(n_818),
.B(n_817),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_845),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_862),
.Y(n_874)
);

CKINVDCx10_ASAP7_75t_R g875 ( 
.A(n_836),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_834),
.B(n_774),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_847),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_847),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_832),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_837),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_844),
.B(n_786),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_832),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_837),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_851),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_833),
.Y(n_885)
);

OAI21x1_ASAP7_75t_L g886 ( 
.A1(n_840),
.A2(n_798),
.B(n_818),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_844),
.B(n_780),
.Y(n_887)
);

AO21x2_ASAP7_75t_L g888 ( 
.A1(n_868),
.A2(n_802),
.B(n_783),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_869),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_862),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_833),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_834),
.B(n_784),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_851),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_838),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_846),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_849),
.Y(n_896)
);

INVx4_ASAP7_75t_SL g897 ( 
.A(n_842),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_845),
.B(n_780),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_843),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_852),
.B(n_829),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_852),
.B(n_816),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_859),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_843),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_875),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_884),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_884),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_899),
.B(n_856),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_899),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_898),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_897),
.B(n_869),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_897),
.B(n_881),
.Y(n_911)
);

OA21x2_ASAP7_75t_L g912 ( 
.A1(n_886),
.A2(n_850),
.B(n_861),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_903),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_895),
.B(n_842),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_898),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_884),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_903),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_893),
.Y(n_918)
);

OAI211xp5_ASAP7_75t_L g919 ( 
.A1(n_876),
.A2(n_824),
.B(n_857),
.C(n_864),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_879),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_897),
.B(n_881),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_897),
.B(n_889),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_893),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_879),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_912),
.Y(n_925)
);

OR2x6_ASAP7_75t_L g926 ( 
.A(n_911),
.B(n_886),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_911),
.B(n_889),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_922),
.B(n_897),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_922),
.B(n_889),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_921),
.B(n_864),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_921),
.B(n_874),
.Y(n_931)
);

INVx1_ASAP7_75t_SL g932 ( 
.A(n_904),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_912),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_909),
.B(n_874),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_909),
.B(n_890),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_909),
.B(n_890),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_915),
.B(n_876),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_905),
.Y(n_938)
);

INVxp67_ASAP7_75t_SL g939 ( 
.A(n_925),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_932),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_937),
.B(n_907),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_928),
.B(n_915),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_938),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_928),
.B(n_915),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_930),
.B(n_910),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_930),
.Y(n_946)
);

NAND3xp33_ASAP7_75t_L g947 ( 
.A(n_933),
.B(n_912),
.C(n_919),
.Y(n_947)
);

OAI21xp33_ASAP7_75t_L g948 ( 
.A1(n_947),
.A2(n_926),
.B(n_892),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_941),
.B(n_914),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_939),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_940),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_939),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_943),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_948),
.A2(n_888),
.B1(n_926),
.B2(n_854),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_951),
.B(n_875),
.Y(n_955)
);

NAND2xp33_ASAP7_75t_SL g956 ( 
.A(n_950),
.B(n_942),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_952),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_949),
.B(n_946),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_958),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_955),
.B(n_942),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_956),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_954),
.B(n_944),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_957),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_958),
.Y(n_964)
);

INVxp67_ASAP7_75t_SL g965 ( 
.A(n_954),
.Y(n_965)
);

INVxp67_ASAP7_75t_L g966 ( 
.A(n_955),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_960),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_966),
.A2(n_945),
.B1(n_953),
.B2(n_841),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_964),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_965),
.A2(n_871),
.B(n_776),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_959),
.Y(n_971)
);

XNOR2x1_ASAP7_75t_L g972 ( 
.A(n_963),
.B(n_871),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_966),
.B(n_894),
.Y(n_973)
);

OAI21xp33_ASAP7_75t_L g974 ( 
.A1(n_967),
.A2(n_962),
.B(n_961),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_R g975 ( 
.A(n_969),
.B(n_902),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_971),
.B(n_855),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_970),
.A2(n_888),
.B(n_929),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_973),
.B(n_934),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_972),
.B(n_935),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_968),
.B(n_936),
.Y(n_980)
);

OAI22xp33_ASAP7_75t_SL g981 ( 
.A1(n_979),
.A2(n_970),
.B1(n_803),
.B2(n_938),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_976),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_975),
.B(n_929),
.Y(n_983)
);

AOI221xp5_ASAP7_75t_L g984 ( 
.A1(n_977),
.A2(n_863),
.B1(n_900),
.B2(n_848),
.C(n_896),
.Y(n_984)
);

AOI221xp5_ASAP7_75t_L g985 ( 
.A1(n_974),
.A2(n_900),
.B1(n_896),
.B2(n_858),
.C(n_821),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_980),
.A2(n_931),
.B(n_927),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_983),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_986),
.B(n_978),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_985),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_981),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_984),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_982),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_982),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_988),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_992),
.B(n_908),
.Y(n_995)
);

NAND3xp33_ASAP7_75t_SL g996 ( 
.A(n_990),
.B(n_778),
.C(n_810),
.Y(n_996)
);

NOR3xp33_ASAP7_75t_L g997 ( 
.A(n_993),
.B(n_775),
.C(n_794),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_987),
.A2(n_913),
.B(n_917),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_989),
.B(n_913),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_994),
.A2(n_991),
.B(n_917),
.Y(n_1000)
);

OAI211xp5_ASAP7_75t_L g1001 ( 
.A1(n_995),
.A2(n_792),
.B(n_805),
.C(n_920),
.Y(n_1001)
);

OAI221xp5_ASAP7_75t_L g1002 ( 
.A1(n_997),
.A2(n_870),
.B1(n_819),
.B2(n_797),
.C(n_860),
.Y(n_1002)
);

NAND3xp33_ASAP7_75t_SL g1003 ( 
.A(n_999),
.B(n_887),
.C(n_901),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_998),
.Y(n_1004)
);

NAND4xp25_ASAP7_75t_L g1005 ( 
.A(n_996),
.B(n_898),
.C(n_887),
.D(n_873),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_1004),
.B(n_924),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_1005),
.A2(n_812),
.B1(n_828),
.B2(n_916),
.Y(n_1007)
);

AO22x2_ASAP7_75t_L g1008 ( 
.A1(n_1003),
.A2(n_923),
.B1(n_918),
.B2(n_916),
.Y(n_1008)
);

OAI221xp5_ASAP7_75t_L g1009 ( 
.A1(n_1002),
.A2(n_860),
.B1(n_831),
.B2(n_916),
.C(n_906),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_1001),
.B(n_905),
.Y(n_1010)
);

AND4x1_ASAP7_75t_L g1011 ( 
.A(n_1000),
.B(n_872),
.C(n_885),
.D(n_882),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_1006),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_1010),
.A2(n_867),
.B1(n_865),
.B2(n_866),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1007),
.A2(n_1009),
.B1(n_1008),
.B2(n_1011),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1006),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1006),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1006),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_1011),
.B(n_873),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_1012),
.B(n_882),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_1015),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1016),
.B(n_891),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_1017),
.B(n_839),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_L g1023 ( 
.A(n_1014),
.B(n_867),
.C(n_865),
.Y(n_1023)
);

NAND4xp75_ASAP7_75t_L g1024 ( 
.A(n_1018),
.B(n_923),
.C(n_918),
.D(n_906),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_1013),
.B(n_866),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_1012),
.B(n_893),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1012),
.B(n_831),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_L g1028 ( 
.A(n_1012),
.B(n_883),
.C(n_880),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_1020),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1026),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1019),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_1022),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_1024),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_1021),
.Y(n_1034)
);

AO22x2_ASAP7_75t_L g1035 ( 
.A1(n_1029),
.A2(n_1023),
.B1(n_1027),
.B2(n_1028),
.Y(n_1035)
);

OAI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_1031),
.A2(n_1025),
.B1(n_796),
.B2(n_880),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_1032),
.B(n_883),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1034),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_1033),
.A2(n_878),
.B1(n_877),
.B2(n_830),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_1034),
.A2(n_878),
.B1(n_877),
.B2(n_830),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1030),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1041),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_1038),
.Y(n_1043)
);

NOR2x1_ASAP7_75t_L g1044 ( 
.A(n_1037),
.B(n_1036),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1043),
.A2(n_1035),
.B1(n_1039),
.B2(n_1040),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_1045),
.Y(n_1046)
);

AO21x2_ASAP7_75t_L g1047 ( 
.A1(n_1046),
.A2(n_1042),
.B(n_1044),
.Y(n_1047)
);

OAI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_1047),
.A2(n_878),
.B1(n_877),
.B2(n_835),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1048),
.A2(n_141),
.B(n_142),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_1049),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_1050)
);

AOI221xp5_ASAP7_75t_L g1051 ( 
.A1(n_1050),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_1051)
);

AOI211xp5_ASAP7_75t_L g1052 ( 
.A1(n_1051),
.A2(n_156),
.B(n_157),
.C(n_158),
.Y(n_1052)
);


endmodule