module fake_jpeg_13218_n_100 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_22),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_10),
.B(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_2),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_4),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_69),
.Y(n_72)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_68),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_49),
.B1(n_27),
.B2(n_50),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

AOI22x1_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_46),
.B1(n_45),
.B2(n_41),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_44),
.B(n_61),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_33),
.C(n_35),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_52),
.C(n_45),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_79),
.B(n_36),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_59),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_77),
.B1(n_80),
.B2(n_73),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_83),
.B1(n_4),
.B2(n_5),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_27),
.B1(n_66),
.B2(n_65),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_33),
.B1(n_64),
.B2(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_86),
.Y(n_89)
);

AOI21x1_ASAP7_75t_SL g92 ( 
.A1(n_88),
.A2(n_84),
.B(n_87),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_17),
.C(n_21),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_81),
.Y(n_94)
);

OA21x2_ASAP7_75t_SL g93 ( 
.A1(n_91),
.A2(n_85),
.B(n_89),
.Y(n_93)
);

A2O1A1O1Ixp25_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_94),
.B(n_14),
.C(n_19),
.D(n_18),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_11),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_25),
.Y(n_97)
);

AOI21x1_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_8),
.B(n_6),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_7),
.Y(n_100)
);


endmodule