module fake_aes_609_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_8), .B(n_6), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_9), .B(n_3), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_2), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_2), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_0), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
BUFx3_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_18), .A2(n_17), .B1(n_13), .B2(n_14), .Y(n_23) );
AOI21xp33_ASAP7_75t_L g24 ( .A1(n_18), .A2(n_13), .B(n_11), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_13), .B1(n_12), .B2(n_11), .Y(n_25) );
BUFx4f_ASAP7_75t_L g26 ( .A(n_19), .Y(n_26) );
INVxp67_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
AOI21xp5_ASAP7_75t_L g28 ( .A1(n_23), .A2(n_22), .B(n_21), .Y(n_28) );
NAND2x1_ASAP7_75t_L g29 ( .A(n_25), .B(n_15), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_16), .Y(n_30) );
AOI33xp33_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_12), .A3(n_16), .B1(n_19), .B2(n_4), .B3(n_5), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_30), .B(n_28), .Y(n_32) );
NAND2xp33_ASAP7_75t_R g33 ( .A(n_30), .B(n_0), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
XOR2xp5_ASAP7_75t_L g35 ( .A(n_33), .B(n_1), .Y(n_35) );
OAI22xp5_ASAP7_75t_L g36 ( .A1(n_32), .A2(n_19), .B1(n_31), .B2(n_15), .Y(n_36) );
NOR2xp33_ASAP7_75t_L g37 ( .A(n_35), .B(n_3), .Y(n_37) );
NOR3x1_ASAP7_75t_L g38 ( .A(n_36), .B(n_4), .C(n_5), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_38), .Y(n_39) );
NAND4xp25_ASAP7_75t_L g40 ( .A(n_37), .B(n_15), .C(n_34), .D(n_6), .Y(n_40) );
AOI22xp33_ASAP7_75t_L g41 ( .A1(n_39), .A2(n_15), .B1(n_26), .B2(n_40), .Y(n_41) );
endmodule