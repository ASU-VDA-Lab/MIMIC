module fake_netlist_6_2546_n_45 (n_7, n_6, n_12, n_4, n_2, n_15, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_10, n_45);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_10;

output n_45;

wire n_41;
wire n_16;
wire n_34;
wire n_42;
wire n_18;
wire n_21;
wire n_24;
wire n_37;
wire n_33;
wire n_27;
wire n_38;
wire n_39;
wire n_32;
wire n_36;
wire n_22;
wire n_26;
wire n_35;
wire n_28;
wire n_17;
wire n_23;
wire n_20;
wire n_30;
wire n_43;
wire n_19;
wire n_29;
wire n_31;
wire n_25;
wire n_40;
wire n_44;

BUFx2_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

AND2x4_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_0),
.Y(n_17)
);

OAI21x1_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_0),
.B(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVxp33_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_17),
.B(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_22),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_17),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OR2x6_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_29),
.Y(n_33)
);

OAI21x1_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_18),
.B(n_22),
.Y(n_34)
);

OAI21x1_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_22),
.B(n_20),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_28),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_32),
.B(n_25),
.Y(n_38)
);

NAND5xp2_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_19),
.C(n_23),
.D(n_21),
.E(n_16),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_32),
.B(n_20),
.C(n_26),
.Y(n_40)
);

OAI221xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_38),
.B1(n_24),
.B2(n_34),
.C(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);


endmodule