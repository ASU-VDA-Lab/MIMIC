module fake_jpeg_17198_n_24 (n_3, n_2, n_1, n_0, n_4, n_5, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_SL g6 ( 
.A(n_4),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

AOI21xp33_ASAP7_75t_L g8 ( 
.A1(n_2),
.A2(n_0),
.B(n_4),
.Y(n_8)
);

AND2x2_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_5),
.Y(n_9)
);

HB1xp67_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_9),
.B(n_1),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_14),
.C(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_15),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_9),
.C(n_7),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g15 ( 
.A1(n_6),
.A2(n_3),
.B1(n_5),
.B2(n_10),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_18),
.C(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_22),
.Y(n_23)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_23),
.B(n_21),
.Y(n_24)
);


endmodule