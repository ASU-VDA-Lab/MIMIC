module fake_jpeg_5460_n_258 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_31;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_34),
.A2(n_37),
.B1(n_39),
.B2(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_15),
.Y(n_48)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_29),
.B1(n_16),
.B2(n_17),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_27),
.B1(n_15),
.B2(n_20),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_52),
.Y(n_74)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_63),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_22),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_20),
.B1(n_30),
.B2(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_18),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_36),
.C(n_39),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_79),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_37),
.B1(n_34),
.B2(n_16),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_72),
.B1(n_84),
.B2(n_55),
.Y(n_91)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_66),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_85),
.B(n_74),
.C(n_19),
.Y(n_106)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_36),
.C(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_37),
.B1(n_34),
.B2(n_39),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_37),
.B1(n_34),
.B2(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_97),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_89),
.B(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_105),
.B1(n_107),
.B2(n_109),
.Y(n_119)
);

AO22x1_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_60),
.B1(n_46),
.B2(n_58),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_100),
.B(n_27),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_52),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_74),
.B(n_60),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_44),
.B(n_15),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_68),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_42),
.B1(n_56),
.B2(n_34),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_106),
.B1(n_86),
.B2(n_25),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_74),
.B(n_48),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_70),
.A2(n_37),
.B1(n_61),
.B2(n_42),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_35),
.B1(n_41),
.B2(n_33),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_67),
.A2(n_35),
.B1(n_41),
.B2(n_33),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_82),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_69),
.A3(n_46),
.B1(n_18),
.B2(n_27),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_115),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_113),
.A2(n_132),
.B(n_25),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_121),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_76),
.CI(n_43),
.CON(n_117),
.SN(n_117)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_117),
.B(n_124),
.Y(n_141)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_78),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_92),
.A2(n_81),
.B1(n_86),
.B2(n_68),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_133),
.B1(n_99),
.B2(n_108),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_30),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_25),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_109),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_25),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_105),
.C(n_107),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_81),
.B1(n_35),
.B2(n_33),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_101),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_41),
.B1(n_35),
.B2(n_33),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_131),
.A2(n_119),
.B1(n_132),
.B2(n_127),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_132)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_147),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_92),
.B1(n_99),
.B2(n_108),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_151),
.B1(n_47),
.B2(n_57),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_94),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_154),
.B(n_113),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_153),
.C(n_119),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_144),
.B(n_155),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_106),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_89),
.B1(n_93),
.B2(n_103),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_149),
.A2(n_122),
.B1(n_124),
.B2(n_117),
.Y(n_170)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_57),
.B1(n_43),
.B2(n_24),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_25),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_57),
.C(n_43),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_167),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_154),
.B(n_141),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_146),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_173),
.B(n_140),
.C(n_137),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_171),
.C(n_143),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

OA21x2_ASAP7_75t_SL g165 ( 
.A1(n_150),
.A2(n_117),
.B(n_115),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_170),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_120),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_144),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_83),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_176),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_83),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_184),
.C(n_190),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_170),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_163),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_159),
.A2(n_147),
.B(n_155),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_181),
.A2(n_187),
.B(n_162),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_140),
.C(n_153),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_191),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_158),
.B(n_24),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_41),
.C(n_35),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_194),
.C(n_157),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_41),
.C(n_47),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_203),
.B(n_208),
.Y(n_214)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_200),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_186),
.B(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_194),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_204),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_160),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_166),
.C(n_176),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_207),
.A2(n_177),
.B(n_187),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_160),
.B(n_174),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_178),
.B(n_174),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_175),
.C(n_24),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_23),
.B(n_1),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_186),
.B1(n_180),
.B2(n_179),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_11),
.B1(n_14),
.B2(n_2),
.Y(n_226)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_196),
.A2(n_187),
.B1(n_185),
.B2(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_192),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_217),
.B(n_202),
.Y(n_224)
);

AO22x1_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_195),
.B1(n_204),
.B2(n_207),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_197),
.A2(n_206),
.B1(n_209),
.B2(n_205),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_1),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_226),
.Y(n_234)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_219),
.Y(n_225)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_225),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_228),
.B(n_1),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_0),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_212),
.B1(n_213),
.B2(n_221),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_229),
.A2(n_216),
.B1(n_220),
.B2(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_215),
.B(n_217),
.Y(n_235)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_236),
.A3(n_239),
.B1(n_2),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_228),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_231),
.A2(n_28),
.B1(n_31),
.B2(n_5),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_SL g239 ( 
.A1(n_231),
.A2(n_24),
.B(n_3),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_230),
.B1(n_227),
.B2(n_225),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_242),
.B(n_244),
.C(n_9),
.Y(n_249)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_223),
.A3(n_21),
.B1(n_31),
.B2(n_10),
.C1(n_11),
.C2(n_5),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_7),
.C(n_9),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_232),
.C(n_21),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_246),
.A2(n_247),
.B(n_249),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_31),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_SL g251 ( 
.A1(n_248),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

NAND2x1p5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_12),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_254),
.A2(n_255),
.B1(n_12),
.B2(n_13),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_31),
.B(n_13),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_253),
.B1(n_13),
.B2(n_14),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_12),
.Y(n_258)
);


endmodule