module fake_jpeg_18566_n_229 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_14),
.B(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_15),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_21),
.B1(n_16),
.B2(n_17),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_24),
.B1(n_27),
.B2(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_14),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_22),
.Y(n_74)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_21),
.B1(n_18),
.B2(n_23),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_38),
.B1(n_21),
.B2(n_28),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_64),
.B1(n_44),
.B2(n_47),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_38),
.B(n_19),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_22),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_45),
.B(n_52),
.C(n_42),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_85),
.B(n_60),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_62),
.B1(n_66),
.B2(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_23),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_91),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_70),
.B1(n_69),
.B2(n_64),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_66),
.C(n_71),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_85),
.C(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_111),
.Y(n_113)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_26),
.B1(n_19),
.B2(n_17),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_52),
.A3(n_18),
.B1(n_23),
.B2(n_75),
.C1(n_65),
.C2(n_31),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_102),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_52),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_109),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_76),
.Y(n_103)
);

XNOR2x2_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_108),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_110),
.B(n_17),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_72),
.B1(n_58),
.B2(n_60),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_59),
.B1(n_50),
.B2(n_51),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_58),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_75),
.B(n_65),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_59),
.B1(n_31),
.B2(n_28),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_90),
.B1(n_80),
.B2(n_59),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_117),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_0),
.B(n_1),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_11),
.C(n_13),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_129),
.B1(n_96),
.B2(n_107),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_79),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_123),
.B1(n_127),
.B2(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_11),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_83),
.B1(n_18),
.B2(n_19),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_109),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_0),
.B(n_3),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_94),
.B(n_11),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_11),
.B1(n_15),
.B2(n_20),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_13),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_135),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_108),
.B(n_107),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_148),
.B(n_152),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_147),
.B1(n_123),
.B2(n_120),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_132),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_0),
.Y(n_150)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_0),
.Y(n_153)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_122),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_163),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_166),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_172),
.B1(n_151),
.B2(n_116),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_155),
.B(n_153),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_140),
.Y(n_168)
);

BUFx4f_ASAP7_75t_SL g177 ( 
.A(n_168),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_132),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_133),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_113),
.B1(n_135),
.B2(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_173),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_155),
.B(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_180),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_147),
.B1(n_159),
.B2(n_138),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_148),
.B(n_143),
.C(n_152),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_129),
.B(n_151),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_158),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_184),
.B(n_176),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_171),
.Y(n_192)
);

AND2x4_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_172),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_174),
.A2(n_154),
.B1(n_167),
.B2(n_169),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_145),
.B1(n_177),
.B2(n_181),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_156),
.B1(n_136),
.B2(n_139),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_194),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_192),
.B(n_186),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_196),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_183),
.C(n_163),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_203),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_187),
.A2(n_156),
.B(n_180),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_177),
.B(n_121),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_3),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_177),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_5),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_183),
.C(n_193),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_9),
.C(n_4),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_212),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_210),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_3),
.B(n_4),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_5),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_213),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_5),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_206),
.A2(n_200),
.B1(n_205),
.B2(n_6),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

OA21x2_ASAP7_75t_SL g219 ( 
.A1(n_209),
.A2(n_6),
.B(n_7),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_217),
.A2(n_216),
.B(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_222),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_218),
.B(n_6),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_215),
.B(n_219),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_221),
.C(n_7),
.Y(n_226)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_225),
.B(n_7),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_7),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);


endmodule