module fake_jpeg_29738_n_58 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx4_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_30),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_19),
.B1(n_23),
.B2(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_0),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_24),
.B1(n_19),
.B2(n_20),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_36),
.B1(n_27),
.B2(n_12),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_29),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_20),
.C(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_43),
.B1(n_3),
.B2(n_4),
.Y(n_46)
);

AO22x1_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_27),
.B1(n_16),
.B2(n_15),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_35),
.B(n_37),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_4),
.C(n_5),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_46),
.B1(n_7),
.B2(n_9),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_49),
.C(n_6),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_5),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_6),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_11),
.C(n_7),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_41),
.B1(n_38),
.B2(n_8),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_53),
.B1(n_10),
.B2(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_52),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_44),
.C(n_50),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_54),
.C(n_55),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_55),
.C(n_10),
.Y(n_58)
);


endmodule