module fake_jpeg_33_n_538 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_538);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_538;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_54),
.B(n_56),
.Y(n_115)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_68),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_62),
.B(n_63),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_20),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_67),
.B(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_29),
.B(n_17),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_84),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_33),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_73),
.B(n_74),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_0),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_86),
.A2(n_38),
.B(n_37),
.C(n_28),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g125 ( 
.A(n_87),
.Y(n_125)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_19),
.B(n_16),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_93),
.Y(n_164)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_35),
.A2(n_48),
.B1(n_45),
.B2(n_47),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_22),
.B1(n_51),
.B2(n_38),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_35),
.B(n_0),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_52),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_43),
.B1(n_40),
.B2(n_39),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_114),
.A2(n_120),
.B1(n_135),
.B2(n_146),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_93),
.A2(n_43),
.B1(n_40),
.B2(n_39),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_69),
.A2(n_48),
.B1(n_45),
.B2(n_43),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_121),
.A2(n_124),
.B1(n_130),
.B2(n_24),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_53),
.A2(n_41),
.B1(n_25),
.B2(n_40),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_126),
.B(n_131),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_86),
.A2(n_52),
.B1(n_51),
.B2(n_22),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_64),
.A2(n_41),
.B1(n_40),
.B2(n_43),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_86),
.A2(n_81),
.B1(n_75),
.B2(n_88),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_132),
.B(n_6),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_80),
.A2(n_83),
.B1(n_96),
.B2(n_97),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_SL g138 ( 
.A(n_72),
.Y(n_138)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g139 ( 
.A1(n_65),
.A2(n_40),
.B1(n_43),
.B2(n_41),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_98),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_151),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_77),
.B(n_92),
.C(n_78),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_101),
.A2(n_37),
.B1(n_28),
.B2(n_26),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_85),
.B(n_26),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_70),
.B(n_23),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_159),
.B(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_91),
.B(n_23),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_125),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_166),
.B(n_168),
.Y(n_272)
);

INVx3_ASAP7_75t_SL g167 ( 
.A(n_106),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_118),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_157),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_169),
.B(n_195),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_170),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_171),
.B(n_174),
.Y(n_251)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_24),
.B(n_94),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_179),
.A2(n_182),
.B1(n_208),
.B2(n_212),
.Y(n_246)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_180),
.Y(n_244)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_116),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_77),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_203),
.C(n_213),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_113),
.B(n_95),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_184),
.B(n_198),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_186),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_188),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_189),
.B(n_193),
.Y(n_257)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_190),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_146),
.A2(n_82),
.B1(n_76),
.B2(n_61),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_164),
.B1(n_156),
.B2(n_136),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_141),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx4_ASAP7_75t_SL g241 ( 
.A(n_194),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_154),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_119),
.A2(n_77),
.B(n_102),
.C(n_59),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_196),
.B(n_202),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_108),
.B(n_59),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_197),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_115),
.B(n_79),
.Y(n_198)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_106),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_200),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_114),
.A2(n_66),
.B1(n_105),
.B2(n_99),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_128),
.B1(n_158),
.B2(n_123),
.Y(n_231)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_139),
.A2(n_103),
.B(n_3),
.C(n_4),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_143),
.B(n_1),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_126),
.A2(n_1),
.B(n_4),
.C(n_5),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_220),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_109),
.Y(n_205)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_138),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_206),
.B(n_207),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_1),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_126),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_209),
.B(n_211),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

INVx13_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_107),
.B(n_5),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_131),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_143),
.B(n_134),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_215),
.B1(n_221),
.B2(n_222),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_120),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_128),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_218),
.Y(n_239)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_219),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_112),
.B(n_7),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_131),
.A2(n_150),
.B1(n_163),
.B2(n_152),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_136),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_148),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_140),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_147),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_225),
.B(n_243),
.C(n_245),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_227),
.A2(n_235),
.B1(n_252),
.B2(n_255),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_231),
.A2(n_234),
.B1(n_171),
.B2(n_230),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_217),
.A2(n_135),
.B1(n_155),
.B2(n_153),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_174),
.A2(n_158),
.B1(n_165),
.B2(n_155),
.Y(n_235)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_238),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_187),
.B(n_149),
.C(n_140),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_177),
.B(n_149),
.C(n_153),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_179),
.B(n_149),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_260),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_182),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_171),
.A2(n_12),
.B1(n_14),
.B2(n_202),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_256),
.A2(n_222),
.B1(n_168),
.B2(n_169),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_180),
.B(n_14),
.C(n_190),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_258),
.B(n_260),
.C(n_170),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_203),
.B(n_14),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_203),
.B(n_189),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_186),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_213),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_270),
.B(n_214),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_273),
.A2(n_312),
.B1(n_252),
.B2(n_262),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_263),
.A2(n_192),
.B(n_214),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_274),
.A2(n_284),
.B(n_287),
.Y(n_336)
);

XNOR2x1_ASAP7_75t_L g276 ( 
.A(n_225),
.B(n_196),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_276),
.B(n_301),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_277),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_195),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_279),
.B(n_289),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_285),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_272),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_291),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_242),
.B(n_178),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_302),
.C(n_314),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_251),
.A2(n_166),
.B(n_215),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_251),
.A2(n_197),
.B1(n_201),
.B2(n_204),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_286),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_251),
.A2(n_213),
.B(n_197),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_236),
.Y(n_288)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_288),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_272),
.B(n_240),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_186),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_290),
.A2(n_296),
.B(n_298),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_244),
.Y(n_292)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

OAI32xp33_ASAP7_75t_L g294 ( 
.A1(n_249),
.A2(n_205),
.A3(n_223),
.B1(n_209),
.B2(n_219),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_294),
.B(n_297),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_229),
.Y(n_295)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_257),
.A2(n_216),
.B1(n_194),
.B2(n_193),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_257),
.A2(n_218),
.B1(n_181),
.B2(n_185),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g298 ( 
.A1(n_259),
.A2(n_167),
.B(n_199),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_248),
.Y(n_299)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_226),
.A2(n_185),
.B1(n_200),
.B2(n_176),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_304),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_242),
.B(n_188),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_247),
.A2(n_246),
.B1(n_234),
.B2(n_226),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_303),
.A2(n_315),
.B(n_250),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_261),
.B(n_172),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_306),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_259),
.A2(n_206),
.B(n_199),
.C(n_167),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_232),
.B(n_200),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_307),
.B(n_316),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_269),
.B(n_188),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_308),
.Y(n_355)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_244),
.Y(n_309)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_264),
.B(n_173),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_266),
.C(n_228),
.Y(n_338)
);

AOI22x1_ASAP7_75t_L g312 ( 
.A1(n_256),
.A2(n_175),
.B1(n_210),
.B2(n_231),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_238),
.Y(n_313)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_313),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_243),
.B(n_210),
.C(n_175),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_232),
.A2(n_239),
.B1(n_224),
.B2(n_241),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_245),
.B(n_210),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_299),
.A2(n_241),
.B1(n_239),
.B2(n_262),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_321),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_322),
.A2(n_327),
.B1(n_341),
.B2(n_297),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_267),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_328),
.C(n_345),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_303),
.A2(n_265),
.B1(n_267),
.B2(n_253),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_283),
.B(n_258),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_307),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_329),
.B(n_352),
.Y(n_384)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_286),
.Y(n_332)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_281),
.A2(n_289),
.B1(n_293),
.B2(n_273),
.Y(n_337)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_337),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_275),
.A2(n_265),
.B1(n_253),
.B2(n_237),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_298),
.A2(n_284),
.B(n_274),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_344),
.A2(n_285),
.B(n_316),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_283),
.B(n_233),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_282),
.B(n_233),
.C(n_266),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_356),
.C(n_305),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_293),
.A2(n_237),
.B1(n_241),
.B2(n_268),
.Y(n_349)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_349),
.Y(n_382)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_350),
.Y(n_361)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_292),
.Y(n_351)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_290),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_353),
.A2(n_287),
.B(n_315),
.Y(n_364)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_276),
.B(n_250),
.C(n_228),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_301),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_367),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_344),
.A2(n_306),
.B(n_296),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_358),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_290),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_362),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g396 ( 
.A(n_364),
.Y(n_396)
);

BUFx24_ASAP7_75t_SL g365 ( 
.A(n_348),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_365),
.B(n_371),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_366),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_275),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_378),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_345),
.B(n_314),
.C(n_313),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_379),
.C(n_385),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_333),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_341),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_372),
.B(n_373),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_354),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_374),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_304),
.Y(n_375)
);

NAND3xp33_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_376),
.C(n_383),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_340),
.B(n_280),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_351),
.Y(n_377)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_377),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_353),
.A2(n_294),
.B(n_310),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_300),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_381),
.B(n_386),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_347),
.B(n_309),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_278),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_342),
.A2(n_312),
.B(n_278),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_323),
.B(n_268),
.C(n_254),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_346),
.C(n_336),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_336),
.A2(n_312),
.B(n_254),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_388),
.B(n_324),
.Y(n_414)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_320),
.Y(n_390)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_390),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_318),
.A2(n_334),
.B1(n_343),
.B2(n_346),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_391),
.A2(n_380),
.B1(n_318),
.B2(n_379),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_360),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_393),
.B(n_402),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_403),
.C(n_409),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_400),
.A2(n_412),
.B1(n_376),
.B2(n_362),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_366),
.A2(n_343),
.B1(n_327),
.B2(n_326),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_362),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_360),
.B(n_317),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_317),
.Y(n_403)
);

FAx1_ASAP7_75t_SL g407 ( 
.A(n_389),
.B(n_356),
.CI(n_326),
.CON(n_407),
.SN(n_407)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_402),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_342),
.C(n_338),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_391),
.A2(n_350),
.B1(n_339),
.B2(n_320),
.Y(n_412)
);

NAND3xp33_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_319),
.C(n_330),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_422),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_414),
.A2(n_378),
.B(n_364),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_387),
.B(n_324),
.C(n_331),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_416),
.C(n_421),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_368),
.B(n_331),
.C(n_339),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_361),
.Y(n_419)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_419),
.Y(n_428)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_361),
.Y(n_420)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_420),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_358),
.B(n_325),
.C(n_330),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_384),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_424),
.A2(n_398),
.B1(n_400),
.B2(n_418),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_449),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_377),
.Y(n_427)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_427),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_410),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_429),
.A2(n_433),
.B1(n_434),
.B2(n_439),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_440),
.Y(n_456)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_394),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_408),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_370),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_435),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_397),
.B(n_370),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_442),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_399),
.B(n_388),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_417),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_404),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_409),
.B(n_407),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_406),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_412),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_446),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_392),
.B(n_393),
.C(n_395),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_444),
.B(n_448),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_405),
.B(n_325),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_445),
.B(n_447),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_396),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_390),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_392),
.B(n_386),
.C(n_374),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_395),
.B(n_381),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_446),
.A2(n_363),
.B1(n_411),
.B2(n_382),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_451),
.A2(n_465),
.B1(n_438),
.B2(n_426),
.Y(n_483)
);

FAx1_ASAP7_75t_SL g454 ( 
.A(n_424),
.B(n_401),
.CI(n_407),
.CON(n_454),
.SN(n_454)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_454),
.B(n_468),
.Y(n_481)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_425),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_441),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_403),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_461),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_462),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_463),
.B(n_450),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_443),
.A2(n_411),
.B1(n_418),
.B2(n_363),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_433),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_466),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_427),
.Y(n_467)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_467),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_435),
.Y(n_468)
);

OA21x2_ASAP7_75t_SL g470 ( 
.A1(n_440),
.A2(n_421),
.B(n_359),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_470),
.Y(n_474)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_472),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_441),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_473),
.B(n_476),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_448),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_478),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_430),
.C(n_449),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_430),
.C(n_437),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_471),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_437),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_485),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_431),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_482),
.B(n_467),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_483),
.B(n_459),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_438),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_490),
.B(n_503),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_465),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_491),
.B(n_478),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_474),
.A2(n_456),
.B(n_469),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_492),
.A2(n_494),
.B(n_497),
.Y(n_516)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_493),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_488),
.A2(n_459),
.B(n_471),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_488),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_496),
.B(n_229),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_SL g498 ( 
.A1(n_480),
.A2(n_453),
.B1(n_462),
.B2(n_436),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_498),
.A2(n_500),
.B1(n_432),
.B2(n_434),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_SL g500 ( 
.A(n_481),
.B(n_452),
.C(n_462),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_485),
.A2(n_453),
.B(n_452),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_501),
.A2(n_487),
.B(n_454),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_486),
.A2(n_454),
.B1(n_466),
.B2(n_442),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_502),
.B(n_486),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_479),
.B(n_484),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_504),
.B(n_477),
.C(n_476),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_505),
.B(n_511),
.Y(n_520)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_506),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_507),
.Y(n_522)
);

AOI21xp33_ASAP7_75t_L g525 ( 
.A1(n_510),
.A2(n_513),
.B(n_515),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_499),
.B(n_428),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_489),
.B(n_428),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_514),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_501),
.A2(n_432),
.B(n_359),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_504),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_517),
.B(n_502),
.Y(n_519)
);

AND2x2_ASAP7_75t_SL g518 ( 
.A(n_508),
.B(n_493),
.Y(n_518)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_518),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_521),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_495),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_505),
.C(n_516),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_527),
.A2(n_525),
.B(n_524),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_522),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_530),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_515),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_526),
.C(n_248),
.Y(n_535)
);

AOI311xp33_ASAP7_75t_L g533 ( 
.A1(n_528),
.A2(n_518),
.A3(n_498),
.B(n_514),
.C(n_495),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_491),
.Y(n_534)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_534),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_532),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_535),
.Y(n_538)
);


endmodule