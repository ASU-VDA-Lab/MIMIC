module fake_jpeg_1500_n_662 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_662);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_662;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_0),
.B(n_1),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_0),
.B(n_10),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_59),
.B(n_60),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_62),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_63),
.B(n_101),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g219 ( 
.A(n_66),
.Y(n_219)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

AND2x4_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_73),
.Y(n_131)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_72),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_79),
.B(n_98),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_80),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_85),
.Y(n_166)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_86),
.Y(n_175)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_87),
.Y(n_174)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_88),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_90),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

BUFx16f_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g130 ( 
.A(n_92),
.Y(n_130)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_93),
.Y(n_188)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_94),
.Y(n_217)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_34),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_99),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_46),
.B(n_17),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_100),
.B(n_104),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_19),
.B(n_17),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_103),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_46),
.B(n_16),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_105),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_57),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_107),
.B(n_110),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_108),
.Y(n_190)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_30),
.B(n_16),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_56),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_111),
.B(n_118),
.Y(n_192)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_25),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_36),
.B(n_2),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_119),
.B(n_124),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_24),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_24),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_24),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_37),
.B(n_2),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_37),
.Y(n_126)
);

BUFx4f_ASAP7_75t_SL g206 ( 
.A(n_126),
.Y(n_206)
);

INVx5_ASAP7_75t_SL g127 ( 
.A(n_25),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_127),
.B(n_55),
.Y(n_207)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_39),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_128),
.B(n_129),
.Y(n_209)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_39),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_92),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_137),
.B(n_139),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_116),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_87),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_140),
.B(n_149),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_61),
.A2(n_30),
.B1(n_27),
.B2(n_23),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_141),
.A2(n_150),
.B1(n_157),
.B2(n_32),
.Y(n_236)
);

INVx6_ASAP7_75t_SL g145 ( 
.A(n_66),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g296 ( 
.A(n_145),
.Y(n_296)
);

BUFx4f_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_148),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_64),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_58),
.B1(n_50),
.B2(n_42),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_110),
.B(n_53),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_156),
.B(n_167),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_30),
.B1(n_23),
.B2(n_27),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_157),
.A2(n_23),
.B1(n_27),
.B2(n_45),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_58),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_158),
.B(n_180),
.Y(n_232)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_160),
.Y(n_237)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_163),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_74),
.B(n_55),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_62),
.B(n_42),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_186),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_72),
.B(n_50),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_203),
.Y(n_235)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_109),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_201),
.B(n_8),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_86),
.B(n_47),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_65),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_97),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_127),
.B(n_40),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_214),
.Y(n_241)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_69),
.Y(n_210)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_210),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_95),
.Y(n_211)
);

INVx11_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_103),
.Y(n_212)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_70),
.B(n_40),
.Y(n_214)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_75),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_77),
.Y(n_220)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_78),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_70),
.B(n_41),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_32),
.Y(n_244)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_80),
.Y(n_223)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_223),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_108),
.B1(n_106),
.B2(n_96),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_224),
.A2(n_254),
.B1(n_285),
.B2(n_133),
.Y(n_315)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_225),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_226),
.B(n_244),
.Y(n_335)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_227),
.Y(n_318)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_132),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_228),
.Y(n_319)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_154),
.Y(n_229)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_229),
.Y(n_349)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_230),
.Y(n_313)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_231),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_99),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_233),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_234),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_236),
.A2(n_171),
.B1(n_173),
.B2(n_138),
.Y(n_333)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_238),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_239),
.B(n_258),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_81),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_243),
.Y(n_343)
);

CKINVDCx12_ASAP7_75t_R g247 ( 
.A(n_219),
.Y(n_247)
);

INVx13_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

AOI21xp33_ASAP7_75t_L g248 ( 
.A1(n_131),
.A2(n_45),
.B(n_25),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_SL g332 ( 
.A(n_248),
.B(n_283),
.Y(n_332)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_249),
.Y(n_346)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_253),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_131),
.A2(n_90),
.B1(n_41),
.B2(n_26),
.Y(n_254)
);

INVx11_ASAP7_75t_L g257 ( 
.A(n_186),
.Y(n_257)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_257),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_209),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_259),
.Y(n_354)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_130),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_261),
.Y(n_356)
);

CKINVDCx12_ASAP7_75t_R g263 ( 
.A(n_130),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_263),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_193),
.B(n_47),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_276),
.Y(n_311)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_159),
.Y(n_267)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_267),
.Y(n_355)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_214),
.A2(n_19),
.B(n_53),
.C(n_26),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_268),
.B(n_282),
.Y(n_320)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_132),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_269),
.Y(n_331)
);

CKINVDCx12_ASAP7_75t_R g270 ( 
.A(n_176),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_270),
.Y(n_308)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_144),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_271),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_192),
.B(n_2),
.Y(n_272)
);

NAND2x1_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_287),
.Y(n_316)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_183),
.Y(n_273)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

OA22x2_ASAP7_75t_L g359 ( 
.A1(n_274),
.A2(n_161),
.B1(n_155),
.B2(n_190),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_193),
.B(n_3),
.Y(n_276)
);

BUFx24_ASAP7_75t_L g277 ( 
.A(n_179),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g339 ( 
.A(n_277),
.Y(n_339)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_168),
.Y(n_278)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_168),
.Y(n_279)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_279),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_153),
.B(n_4),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_289),
.Y(n_326)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_178),
.Y(n_281)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_207),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g283 ( 
.A(n_222),
.B(n_84),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_134),
.Y(n_284)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_284),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_153),
.A2(n_45),
.B1(n_82),
.B2(n_54),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_164),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_286),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_169),
.B(n_146),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_169),
.B(n_4),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_141),
.A2(n_54),
.B1(n_38),
.B2(n_29),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_290),
.A2(n_147),
.B1(n_135),
.B2(n_152),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_177),
.B(n_5),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_295),
.Y(n_329)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_136),
.Y(n_292)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_292),
.Y(n_345)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_211),
.Y(n_293)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_177),
.B(n_5),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_208),
.B(n_5),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_297),
.B(n_218),
.Y(n_344)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_175),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_176),
.Y(n_299)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_178),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_300),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_142),
.B(n_6),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_302),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_194),
.B(n_6),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_179),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_307),
.B(n_344),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_235),
.A2(n_195),
.B1(n_148),
.B2(n_205),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_312),
.A2(n_136),
.B1(n_161),
.B2(n_155),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_315),
.A2(n_359),
.B1(n_362),
.B2(n_234),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_317),
.A2(n_338),
.B1(n_348),
.B2(n_296),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_333),
.A2(n_337),
.B1(n_350),
.B2(n_362),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_264),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_251),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_290),
.A2(n_174),
.B1(n_170),
.B2(n_190),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_254),
.A2(n_174),
.B1(n_170),
.B2(n_143),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_233),
.B(n_217),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_347),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_241),
.A2(n_213),
.B1(n_218),
.B2(n_138),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_243),
.A2(n_185),
.B1(n_165),
.B2(n_182),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_287),
.B(n_188),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_353),
.B(n_245),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_232),
.B(n_204),
.C(n_200),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_357),
.B(n_172),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_226),
.A2(n_272),
.B1(n_283),
.B2(n_248),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_363),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_274),
.A2(n_163),
.B1(n_191),
.B2(n_196),
.Y(n_362)
);

OAI22x1_ASAP7_75t_L g363 ( 
.A1(n_285),
.A2(n_54),
.B1(n_38),
.B2(n_204),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_364),
.Y(n_419)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_314),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_372),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_366),
.B(n_373),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_367),
.Y(n_413)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_318),
.Y(n_368)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

INVx13_ASAP7_75t_L g369 ( 
.A(n_358),
.Y(n_369)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_369),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_340),
.A2(n_256),
.B1(n_224),
.B2(n_189),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_370),
.A2(n_408),
.B1(n_228),
.B2(n_269),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_332),
.A2(n_361),
.B(n_320),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_371),
.A2(n_360),
.B(n_323),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_311),
.B(n_283),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_306),
.B(n_298),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_268),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_374),
.B(n_377),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_304),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_376),
.B(n_396),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_316),
.B(n_227),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_378),
.A2(n_383),
.B1(n_386),
.B2(n_395),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_316),
.B(n_303),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_379),
.B(n_382),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_337),
.A2(n_189),
.B1(n_185),
.B2(n_182),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_380),
.A2(n_409),
.B1(n_410),
.B2(n_305),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_234),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_335),
.B(n_271),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_338),
.A2(n_252),
.B1(n_296),
.B2(n_242),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_328),
.Y(n_385)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_385),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_359),
.A2(n_252),
.B1(n_242),
.B2(n_237),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_313),
.Y(n_387)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_387),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_260),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_326),
.B(n_265),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_390),
.B(n_398),
.Y(n_436)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_325),
.Y(n_392)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_392),
.Y(n_433)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_345),
.Y(n_393)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_393),
.Y(n_445)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_345),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_394),
.Y(n_421)
);

INVx13_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_313),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_329),
.B(n_260),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_397),
.B(n_399),
.Y(n_441)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_322),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_322),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_400),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_335),
.B(n_265),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_401),
.B(n_402),
.Y(n_442)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_317),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_309),
.B(n_246),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_403),
.B(n_404),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_310),
.B(n_246),
.Y(n_404)
);

INVx13_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_356),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_406),
.B(n_363),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_343),
.B(n_284),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_407),
.B(n_342),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_359),
.A2(n_165),
.B1(n_143),
.B2(n_172),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_332),
.A2(n_262),
.B1(n_255),
.B2(n_275),
.Y(n_409)
);

NAND2xp33_ASAP7_75t_SL g484 ( 
.A(n_414),
.B(n_424),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_415),
.B(n_429),
.C(n_434),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_374),
.A2(n_333),
.B1(n_350),
.B2(n_262),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_416),
.B(n_427),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_423),
.B(n_380),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_409),
.A2(n_346),
.B1(n_355),
.B2(n_321),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_308),
.C(n_349),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_342),
.B1(n_319),
.B2(n_331),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_432),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_391),
.A2(n_378),
.B1(n_367),
.B2(n_408),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_360),
.C(n_323),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_435),
.A2(n_443),
.B1(n_389),
.B2(n_385),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_438),
.A2(n_407),
.B(n_382),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_391),
.A2(n_305),
.B(n_351),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_440),
.A2(n_438),
.B(n_442),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_410),
.A2(n_292),
.B1(n_275),
.B2(n_255),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_391),
.A2(n_370),
.B1(n_386),
.B2(n_372),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_449),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_448),
.B(n_401),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_377),
.A2(n_240),
.B1(n_331),
.B2(n_319),
.Y(n_449)
);

INVx13_ASAP7_75t_L g450 ( 
.A(n_446),
.Y(n_450)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_450),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_411),
.B(n_376),
.Y(n_451)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_451),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_412),
.Y(n_453)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_453),
.Y(n_502)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_439),
.Y(n_455)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_455),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_456),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_476),
.Y(n_493)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_418),
.Y(n_458)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_458),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_412),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_459),
.B(n_462),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_460),
.A2(n_466),
.B1(n_383),
.B2(n_327),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_461),
.A2(n_447),
.B1(n_416),
.B2(n_413),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_412),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_414),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_463),
.B(n_467),
.Y(n_509)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_418),
.Y(n_464)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_464),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_SL g466 ( 
.A1(n_432),
.A2(n_385),
.B1(n_381),
.B2(n_327),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_414),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_444),
.B(n_397),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_469),
.B(n_485),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_436),
.B(n_390),
.Y(n_470)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_470),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_421),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_471),
.B(n_473),
.Y(n_512)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_426),
.Y(n_472)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_472),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_446),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_426),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_474),
.B(n_475),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_436),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_445),
.Y(n_476)
);

AND2x2_ASAP7_75t_SL g477 ( 
.A(n_442),
.B(n_379),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_SL g498 ( 
.A1(n_477),
.A2(n_417),
.B(n_448),
.C(n_441),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_478),
.A2(n_484),
.B(n_456),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_422),
.B(n_384),
.C(n_373),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_429),
.C(n_422),
.Y(n_486)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_419),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_483),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_420),
.B(n_404),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_481),
.B(n_482),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_437),
.B(n_403),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_444),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_445),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_486),
.B(n_504),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_488),
.A2(n_511),
.B1(n_508),
.B2(n_461),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_491),
.A2(n_498),
.B(n_511),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_434),
.C(n_417),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_492),
.B(n_497),
.C(n_477),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_468),
.A2(n_413),
.B1(n_423),
.B2(n_443),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_495),
.A2(n_503),
.B1(n_507),
.B2(n_510),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_451),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_496),
.B(n_388),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_479),
.C(n_457),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_483),
.B(n_366),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_499),
.B(n_368),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_468),
.A2(n_440),
.B1(n_415),
.B2(n_427),
.Y(n_503)
);

XOR2x2_ASAP7_75t_SL g504 ( 
.A(n_470),
.B(n_430),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_454),
.A2(n_435),
.B1(n_428),
.B2(n_449),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_454),
.A2(n_428),
.B1(n_430),
.B2(n_431),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_478),
.A2(n_425),
.B(n_424),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_452),
.A2(n_462),
.B1(n_459),
.B2(n_453),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_513),
.A2(n_515),
.B1(n_452),
.B2(n_463),
.Y(n_524)
);

AOI322xp5_ASAP7_75t_SL g514 ( 
.A1(n_469),
.A2(n_375),
.A3(n_365),
.B1(n_399),
.B2(n_395),
.C1(n_369),
.C2(n_437),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_514),
.B(n_395),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_455),
.B(n_375),
.Y(n_518)
);

CKINVDCx14_ASAP7_75t_R g530 ( 
.A(n_518),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_521),
.B(n_533),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_492),
.B(n_477),
.C(n_482),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_523),
.B(n_527),
.C(n_532),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_524),
.A2(n_549),
.B1(n_550),
.B2(n_501),
.Y(n_555)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_509),
.Y(n_525)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_525),
.Y(n_552)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_509),
.Y(n_526)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_526),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_497),
.B(n_477),
.C(n_475),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_512),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_528),
.B(n_512),
.Y(n_553)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_490),
.Y(n_529)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_529),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_486),
.B(n_481),
.C(n_471),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_500),
.B(n_493),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_490),
.Y(n_534)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_534),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_493),
.B(n_484),
.Y(n_535)
);

MAJx2_ASAP7_75t_L g557 ( 
.A(n_535),
.B(n_539),
.C(n_541),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_495),
.A2(n_516),
.B1(n_507),
.B2(n_510),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_536),
.B(n_544),
.Y(n_570)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_538),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_493),
.B(n_472),
.Y(n_539)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_540),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_504),
.B(n_513),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_519),
.Y(n_542)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_542),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_520),
.B(n_474),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_506),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_489),
.B(n_341),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_491),
.A2(n_467),
.B(n_476),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_545),
.A2(n_498),
.B(n_487),
.Y(n_562)
);

NOR3xp33_ASAP7_75t_SL g567 ( 
.A(n_546),
.B(n_369),
.C(n_498),
.Y(n_567)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_519),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_547),
.B(n_548),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_488),
.A2(n_517),
.B1(n_503),
.B2(n_505),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_502),
.A2(n_461),
.B1(n_464),
.B2(n_458),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_520),
.A2(n_461),
.B1(n_485),
.B2(n_460),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_551),
.A2(n_508),
.B1(n_494),
.B2(n_505),
.Y(n_554)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_553),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_554),
.B(n_537),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_555),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_558),
.B(n_574),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_521),
.B(n_473),
.C(n_501),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_560),
.B(n_568),
.C(n_572),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_533),
.B(n_506),
.Y(n_561)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_561),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_562),
.A2(n_545),
.B(n_535),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_524),
.A2(n_498),
.B1(n_487),
.B2(n_480),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_SL g565 ( 
.A(n_541),
.B(n_498),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_565),
.B(n_537),
.Y(n_581)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_567),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_532),
.B(n_433),
.C(n_351),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_522),
.B(n_433),
.C(n_393),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_527),
.B(n_387),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_559),
.B(n_569),
.C(n_560),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_577),
.B(n_579),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_559),
.B(n_522),
.C(n_523),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_581),
.A2(n_583),
.B1(n_563),
.B2(n_552),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_569),
.B(n_528),
.C(n_531),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_582),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_585),
.B(n_554),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_568),
.B(n_543),
.C(n_539),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_595),
.C(n_558),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_562),
.A2(n_530),
.B(n_549),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_587),
.A2(n_590),
.B(n_594),
.Y(n_599)
);

CKINVDCx16_ASAP7_75t_R g588 ( 
.A(n_561),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_588),
.A2(n_576),
.B1(n_567),
.B2(n_334),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_572),
.A2(n_550),
.B(n_419),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_574),
.B(n_394),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_592),
.B(n_593),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_557),
.B(n_364),
.Y(n_593)
);

A2O1A1O1Ixp25_ASAP7_75t_L g594 ( 
.A1(n_565),
.A2(n_450),
.B(n_398),
.C(n_392),
.D(n_405),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_557),
.B(n_324),
.C(n_450),
.Y(n_595)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_598),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_600),
.B(n_605),
.Y(n_617)
);

MAJx2_ASAP7_75t_L g602 ( 
.A(n_583),
.B(n_564),
.C(n_553),
.Y(n_602)
);

MAJx2_ASAP7_75t_L g618 ( 
.A(n_602),
.B(n_608),
.C(n_593),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_580),
.B(n_555),
.C(n_570),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_604),
.A2(n_606),
.B(n_613),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_580),
.B(n_566),
.C(n_556),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_591),
.B(n_571),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_607),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_591),
.B(n_573),
.Y(n_608)
);

INVx11_ASAP7_75t_L g609 ( 
.A(n_594),
.Y(n_609)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_609),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_582),
.B(n_575),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_610),
.B(n_592),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_612),
.B(n_597),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_SL g613 ( 
.A1(n_585),
.A2(n_334),
.B(n_405),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_589),
.A2(n_240),
.B1(n_237),
.B2(n_288),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_614),
.A2(n_596),
.B1(n_597),
.B2(n_589),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_586),
.B(n_324),
.C(n_288),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_615),
.B(n_595),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_618),
.B(n_599),
.Y(n_630)
);

MAJx2_ASAP7_75t_L g621 ( 
.A(n_600),
.B(n_584),
.C(n_578),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_621),
.B(n_598),
.Y(n_637)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_622),
.Y(n_633)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_623),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_624),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_625),
.B(n_608),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_604),
.A2(n_196),
.B1(n_200),
.B2(n_330),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_626),
.A2(n_609),
.B1(n_606),
.B2(n_615),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_601),
.B(n_341),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_628),
.B(n_611),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_605),
.A2(n_294),
.B(n_261),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_629),
.A2(n_294),
.B(n_286),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_630),
.B(n_637),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_SL g631 ( 
.A1(n_620),
.A2(n_602),
.B(n_607),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_631),
.A2(n_638),
.B1(n_640),
.B2(n_250),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_632),
.B(n_639),
.C(n_617),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_SL g644 ( 
.A1(n_634),
.A2(n_619),
.B1(n_618),
.B2(n_621),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_627),
.A2(n_603),
.B(n_611),
.Y(n_638)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_641),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_633),
.B(n_616),
.C(n_617),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_642),
.B(n_643),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_636),
.B(n_619),
.C(n_625),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_644),
.B(n_645),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_635),
.A2(n_257),
.B1(n_250),
.B2(n_191),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_634),
.B(n_330),
.C(n_245),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_646),
.A2(n_647),
.B(n_630),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_648),
.B(n_631),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_649),
.B(n_652),
.Y(n_655)
);

AOI322xp5_ASAP7_75t_L g654 ( 
.A1(n_653),
.A2(n_645),
.A3(n_339),
.B1(n_293),
.B2(n_299),
.C1(n_24),
.C2(n_277),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_654),
.B(n_656),
.C(n_651),
.Y(n_657)
);

AOI322xp5_ASAP7_75t_L g656 ( 
.A1(n_650),
.A2(n_339),
.A3(n_277),
.B1(n_38),
.B2(n_14),
.C1(n_9),
.C2(n_12),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g659 ( 
.A1(n_657),
.A2(n_658),
.B1(n_9),
.B2(n_14),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_655),
.B(n_339),
.C(n_11),
.Y(n_658)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_659),
.B(n_9),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_660),
.B(n_15),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_661),
.A2(n_15),
.B1(n_385),
.B2(n_358),
.Y(n_662)
);


endmodule