module real_jpeg_24162_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_344, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_344;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_2),
.A2(n_33),
.B1(n_36),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_2),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_2),
.A2(n_29),
.B1(n_44),
.B2(n_128),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_2),
.A2(n_52),
.B1(n_53),
.B2(n_128),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_2),
.A2(n_58),
.B1(n_59),
.B2(n_128),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_4),
.A2(n_44),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_4),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_4),
.B(n_32),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g207 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_137),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_4),
.B(n_54),
.C(n_59),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_4),
.B(n_67),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_4),
.A2(n_109),
.B1(n_235),
.B2(n_240),
.Y(n_239)
);

INVx8_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_6),
.A2(n_33),
.B1(n_36),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_6),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_130),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_130),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_6),
.A2(n_25),
.B1(n_43),
.B2(n_130),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_7),
.A2(n_29),
.B1(n_39),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_7),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_7),
.A2(n_33),
.B1(n_36),
.B2(n_140),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_7),
.A2(n_52),
.B1(n_53),
.B2(n_140),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_140),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_8),
.A2(n_27),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_8),
.A2(n_33),
.B1(n_36),
.B2(n_42),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_8),
.A2(n_42),
.B1(n_58),
.B2(n_59),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_8),
.A2(n_42),
.B1(n_52),
.B2(n_53),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_9),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_9),
.A2(n_28),
.B1(n_52),
.B2(n_53),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_9),
.A2(n_28),
.B1(n_58),
.B2(n_59),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_9),
.A2(n_28),
.B1(n_33),
.B2(n_36),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_11),
.A2(n_33),
.B1(n_36),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_74),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_74),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_74),
.Y(n_116)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_14),
.A2(n_33),
.B1(n_36),
.B2(n_62),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_14),
.A2(n_29),
.B1(n_44),
.B2(n_62),
.Y(n_298)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_15),
.Y(n_112)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_15),
.Y(n_221)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_15),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_95),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_93),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_85),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_85),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.C(n_79),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_20),
.A2(n_21),
.B1(n_75),
.B2(n_330),
.Y(n_336)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_46),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_22),
.B(n_48),
.C(n_63),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B1(n_32),
.B2(n_41),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_24),
.A2(n_31),
.B(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_26),
.B(n_137),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_26),
.B(n_35),
.C(n_36),
.Y(n_152)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_30),
.B(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_30),
.A2(n_41),
.B(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_30),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_30),
.A2(n_32),
.B1(n_139),
.B2(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_30),
.A2(n_32),
.B1(n_147),
.B2(n_275),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_30),
.A2(n_275),
.B(n_297),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_30),
.A2(n_89),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_38),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_31),
.B(n_78),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_31),
.A2(n_133),
.B1(n_134),
.B2(n_138),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_31),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_33),
.A2(n_36),
.B1(n_68),
.B2(n_69),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_33),
.A2(n_37),
.B(n_136),
.C(n_152),
.Y(n_151)
);

HAxp5_ASAP7_75t_SL g180 ( 
.A(n_33),
.B(n_137),
.CON(n_180),
.SN(n_180)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_36),
.A2(n_53),
.A3(n_68),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_63),
.B2(n_64),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_75),
.C(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_47),
.A2(n_48),
.B1(n_80),
.B2(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_57),
.B(n_60),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_50),
.B(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_50),
.A2(n_61),
.B(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_50),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_50),
.A2(n_189),
.B(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_50),
.A2(n_188),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_50),
.A2(n_187),
.B1(n_188),
.B2(n_208),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_50),
.A2(n_188),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_50),
.A2(n_124),
.B(n_269),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_53),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_52),
.B(n_69),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_53),
.B(n_210),
.Y(n_209)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_54),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_57),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_57),
.B(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_57),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_57),
.B(n_60),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_57),
.B(n_137),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_58),
.B(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_70),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_65),
.A2(n_126),
.B(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_67),
.B(n_71),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_66),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_67),
.A2(n_71),
.B1(n_171),
.B2(n_180),
.Y(n_185)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_70),
.A2(n_131),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_81),
.B(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_75),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_75),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_79),
.B(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_80),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_82),
.A2(n_126),
.B1(n_131),
.B2(n_301),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_84),
.A2(n_126),
.B(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_92),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI321xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_327),
.A3(n_337),
.B1(n_340),
.B2(n_341),
.C(n_344),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_306),
.B(n_326),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_283),
.B(n_305),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_172),
.B(n_259),
.C(n_282),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_157),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_100),
.B(n_157),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_143),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_121),
.B1(n_141),
.B2(n_142),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_102),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_102),
.B(n_142),
.C(n_143),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_103),
.B(n_108),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_104),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_105),
.B(n_313),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_113),
.B(n_115),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_109),
.A2(n_115),
.B(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_109),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_109),
.A2(n_226),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_109),
.A2(n_183),
.B(n_236),
.Y(n_291)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_110),
.A2(n_114),
.B1(n_119),
.B2(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_110),
.B(n_116),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_110),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_112),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_120),
.Y(n_244)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.C(n_132),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_137),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_150),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_146),
.B(n_148),
.C(n_150),
.Y(n_280)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_153),
.B1(n_154),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_163),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_158),
.B(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_161),
.B(n_163),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.C(n_169),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_167),
.B1(n_168),
.B2(n_194),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_164),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_166),
.B(n_219),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_254),
.B(n_258),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_202),
.B(n_253),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_190),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_177),
.B(n_190),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_185),
.C(n_186),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_178),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_185),
.B(n_186),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_191),
.B(n_198),
.C(n_201),
.Y(n_255)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_197),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_200),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_248),
.B(n_252),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_222),
.B(n_247),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_211),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_205),
.B(n_211),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_209),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_216),
.C(n_217),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_215),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_231),
.B(n_246),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_230),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_238),
.B(n_245),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_250),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_255),
.B(n_256),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_261),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_280),
.B2(n_281),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_271),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_271),
.C(n_281),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_270),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_270),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_267),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_279),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_276),
.C(n_279),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_284),
.B(n_285),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_304),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_292),
.B1(n_302),
.B2(n_303),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_303),
.C(n_304),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_290),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_290),
.A2(n_291),
.B1(n_318),
.B2(n_320),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_290),
.A2(n_320),
.B(n_321),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_296),
.C(n_299),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_299),
.B2(n_300),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_307),
.B(n_308),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_324),
.B2(n_325),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_316),
.B1(n_322),
.B2(n_323),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_311),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_323),
.C(n_325),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_314),
.B(n_315),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_314),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_329),
.C(n_334),
.Y(n_328)
);

FAx1_ASAP7_75t_SL g339 ( 
.A(n_315),
.B(n_329),
.CI(n_334),
.CON(n_339),
.SN(n_339)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_321),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_318),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_335),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_335),
.Y(n_341)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_338),
.B(n_339),
.Y(n_340)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_339),
.Y(n_342)
);


endmodule