module fake_netlist_6_280_n_105 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_10, n_105);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_10;

output n_105;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_18;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_17;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_97;
wire n_94;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVxp67_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_22),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_26),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

OR2x6_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

OAI221xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_19),
.B1(n_18),
.B2(n_27),
.C(n_29),
.Y(n_52)
);

AO22x2_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AND2x6_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

AOI221xp5_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_27),
.B1(n_35),
.B2(n_38),
.C(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_54),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_60),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_61),
.B(n_63),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_48),
.B(n_33),
.C(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_71),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_74),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g78 ( 
.A(n_74),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_77),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_69),
.B1(n_49),
.B2(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_75),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_37),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_83),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_84),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_41),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_81),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_41),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2x1p5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_93),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_91),
.B(n_39),
.Y(n_99)
);

NAND4xp75_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_37),
.C(n_53),
.D(n_7),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_94),
.B(n_40),
.C(n_42),
.Y(n_101)
);

NAND4xp25_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_94),
.C(n_40),
.D(n_98),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_53),
.B(n_100),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_53),
.B(n_42),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_42),
.B1(n_6),
.B2(n_5),
.Y(n_105)
);


endmodule