module fake_jpeg_2842_n_193 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_193);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_4),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_1),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_63),
.B1(n_62),
.B2(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_49),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_86),
.B1(n_76),
.B2(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_92),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_54),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_66),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_63),
.B1(n_62),
.B2(n_68),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_54),
.B1(n_65),
.B2(n_67),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_76),
.B1(n_74),
.B2(n_72),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_64),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_77),
.B1(n_65),
.B2(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_70),
.B1(n_88),
.B2(n_55),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_106),
.B1(n_88),
.B2(n_84),
.Y(n_118)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_57),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_55),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_74),
.B1(n_72),
.B2(n_66),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_108),
.Y(n_111)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_110),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_58),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_121),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_61),
.C(n_59),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_9),
.C(n_10),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_125),
.B1(n_95),
.B2(n_91),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_58),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_117),
.C(n_112),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_56),
.B1(n_51),
.B2(n_91),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_130),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_70),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_3),
.CI(n_5),
.CON(n_136),
.SN(n_136)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_16),
.A3(n_18),
.B1(n_19),
.B2(n_20),
.C1(n_21),
.C2(n_22),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_105),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_145),
.C(n_151),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_142),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_143),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_147),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_122),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_126),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_150),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_14),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_148),
.B(n_149),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_15),
.Y(n_149)
);

INVxp33_ASAP7_75t_SL g150 ( 
.A(n_122),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_31),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_16),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_25),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_164),
.B(n_151),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_129),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_142),
.C(n_29),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_165),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_23),
.B(n_24),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_131),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_168),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_175),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_134),
.B1(n_144),
.B2(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_172),
.C(n_177),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_27),
.B(n_33),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_34),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_36),
.C(n_37),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_171),
.C(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_183),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_167),
.A3(n_155),
.B1(n_159),
.B2(n_153),
.C1(n_162),
.C2(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_184),
.B(n_185),
.Y(n_189)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_177),
.C(n_167),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_180),
.C(n_164),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_186),
.A3(n_155),
.B1(n_162),
.B2(n_42),
.C1(n_43),
.C2(n_38),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_190),
.A2(n_189),
.B(n_41),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_40),
.B(n_45),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_47),
.Y(n_193)
);


endmodule