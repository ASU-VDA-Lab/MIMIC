module fake_netlist_6_3175_n_1937 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_597, n_280, n_287, n_353, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_581, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_92, n_599, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1937);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_599;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1937;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_917;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1054;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_699;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_1918;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_608;
wire n_630;
wire n_792;
wire n_1328;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1563;
wire n_1912;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_1165;
wire n_702;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_1520;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_937;
wire n_1682;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_776;
wire n_1823;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_879;
wire n_959;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_652;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_1028;
wire n_1922;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_861;
wire n_857;
wire n_967;
wire n_1884;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_1260;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_1423;
wire n_1935;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_506),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_235),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_24),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_582),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_95),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_528),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_34),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_186),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_549),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_400),
.Y(n_616)
);

CKINVDCx16_ASAP7_75t_R g617 ( 
.A(n_233),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_566),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_75),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_320),
.Y(n_620)
);

CKINVDCx6p67_ASAP7_75t_R g621 ( 
.A(n_552),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_600),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_213),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_603),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_30),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_567),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_87),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_202),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_599),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_581),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_384),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_589),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_40),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_46),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_290),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_123),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_372),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_316),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_327),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_592),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_30),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_541),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_64),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_123),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_291),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_319),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_312),
.Y(n_647)
);

BUFx8_ASAP7_75t_SL g648 ( 
.A(n_290),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_76),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_543),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_201),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_93),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_533),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_587),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_524),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_538),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_440),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_51),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_369),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_586),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_243),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_605),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_596),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_526),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_525),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_604),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_575),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_322),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_88),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_406),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_423),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_504),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_218),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_545),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_583),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_444),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_106),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_12),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_88),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_532),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_119),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_13),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_415),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_536),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_247),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_152),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_354),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_426),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_321),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_420),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_505),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_562),
.Y(n_692)
);

BUFx10_ASAP7_75t_L g693 ( 
.A(n_199),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_577),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_547),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_591),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_439),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_544),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_502),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_601),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_61),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_28),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_523),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_595),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_342),
.Y(n_705)
);

BUFx8_ASAP7_75t_SL g706 ( 
.A(n_602),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_274),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_265),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_401),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_302),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_111),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_144),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_76),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_287),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_195),
.Y(n_715)
);

BUFx10_ASAP7_75t_L g716 ( 
.A(n_64),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_246),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_87),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_301),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_590),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_300),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_388),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_7),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_393),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_323),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_5),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_561),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_594),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_108),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_138),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_499),
.Y(n_731)
);

INVx1_ASAP7_75t_SL g732 ( 
.A(n_574),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_399),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_559),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_573),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_430),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_236),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_260),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_209),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_569),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_529),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_344),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_530),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_223),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_578),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_218),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_267),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_404),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_32),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_338),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_564),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_553),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_35),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_531),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_490),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_374),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_141),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_593),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_65),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_56),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_124),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_511),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_570),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_515),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_171),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_118),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_563),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_244),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_413),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_157),
.Y(n_770)
);

CKINVDCx14_ASAP7_75t_R g771 ( 
.A(n_277),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_387),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_606),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_537),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_96),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_555),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_498),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_45),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_468),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_571),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_73),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_548),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_287),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_585),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_535),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_542),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_340),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_363),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_84),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_197),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_330),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_557),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_222),
.Y(n_793)
);

BUFx10_ASAP7_75t_L g794 ( 
.A(n_116),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_358),
.Y(n_795)
);

BUFx10_ASAP7_75t_L g796 ( 
.A(n_325),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_234),
.Y(n_797)
);

BUFx8_ASAP7_75t_SL g798 ( 
.A(n_49),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_576),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_171),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_234),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_554),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_235),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_441),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_117),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_306),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_598),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_135),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_185),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_145),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_588),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_261),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_556),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_568),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_225),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_580),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_383),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_65),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_551),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_437),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_19),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_436),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_558),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_295),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_546),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_539),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_54),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_597),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_54),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_391),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_579),
.Y(n_831)
);

BUFx5_ASAP7_75t_L g832 ( 
.A(n_136),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_560),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_550),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_534),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_364),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_422),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_339),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_274),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_138),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_456),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_288),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_477),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_527),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_101),
.Y(n_845)
);

CKINVDCx16_ASAP7_75t_R g846 ( 
.A(n_455),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_201),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_210),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_42),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_324),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_565),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_572),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_584),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_397),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_285),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_540),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_45),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_832),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_832),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_832),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_656),
.B(n_1),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_832),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_832),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_637),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_830),
.B(n_1),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_706),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_648),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_798),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_701),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_701),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_607),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_655),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_701),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_686),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_616),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_617),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_719),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_615),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_719),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_839),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_624),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_629),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_753),
.Y(n_883)
);

CKINVDCx16_ASAP7_75t_R g884 ( 
.A(n_846),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_719),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_677),
.B(n_0),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_717),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_873),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_871),
.B(n_612),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_875),
.B(n_650),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_881),
.B(n_670),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_873),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_882),
.B(n_687),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_876),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_869),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_870),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_877),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_864),
.B(n_838),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_879),
.Y(n_899)
);

NAND2xp33_ASAP7_75t_SL g900 ( 
.A(n_874),
.B(n_809),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_872),
.B(n_694),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_887),
.B(n_785),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_885),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_868),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_858),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_860),
.B(n_825),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_859),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_862),
.Y(n_908)
);

OA21x2_ASAP7_75t_L g909 ( 
.A1(n_863),
.A2(n_622),
.B(n_610),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_886),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_861),
.B(n_841),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_865),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_884),
.B(n_883),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_880),
.B(n_672),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_866),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_883),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_867),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_894),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_912),
.B(n_642),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_901),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_907),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_888),
.B(n_742),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_895),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_895),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_913),
.Y(n_925)
);

AND2x6_ASAP7_75t_L g926 ( 
.A(n_905),
.B(n_618),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_889),
.B(n_771),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_896),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_890),
.B(n_878),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_902),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_891),
.B(n_817),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_896),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_897),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_901),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_916),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_908),
.Y(n_936)
);

OAI22xp33_ASAP7_75t_SL g937 ( 
.A1(n_911),
.A2(n_723),
.B1(n_638),
.B2(n_643),
.Y(n_937)
);

INVx5_ASAP7_75t_L g938 ( 
.A(n_915),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_892),
.B(n_662),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_917),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_899),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_903),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_910),
.B(n_692),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_906),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_909),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_893),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_898),
.B(n_636),
.Y(n_947)
);

XNOR2xp5_ASAP7_75t_L g948 ( 
.A(n_904),
.B(n_722),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_909),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_914),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_900),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_901),
.B(n_724),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_894),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_912),
.A2(n_812),
.B1(n_818),
.B2(n_809),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_888),
.B(n_732),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_912),
.B(n_735),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_905),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_905),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_915),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_941),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_920),
.B(n_793),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_921),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_942),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_930),
.B(n_636),
.Y(n_964)
);

AO22x2_ASAP7_75t_L g965 ( 
.A1(n_956),
.A2(n_726),
.B1(n_790),
.B2(n_633),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_924),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_957),
.Y(n_967)
);

AO22x2_ASAP7_75t_L g968 ( 
.A1(n_951),
.A2(n_824),
.B1(n_619),
.B2(n_652),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_944),
.B(n_626),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_958),
.Y(n_970)
);

AO22x2_ASAP7_75t_L g971 ( 
.A1(n_943),
.A2(n_689),
.B1(n_708),
.B2(n_682),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_933),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_935),
.Y(n_973)
);

AO22x2_ASAP7_75t_L g974 ( 
.A1(n_952),
.A2(n_797),
.B1(n_669),
.B2(n_681),
.Y(n_974)
);

NAND2x1p5_ASAP7_75t_L g975 ( 
.A(n_938),
.B(n_733),
.Y(n_975)
);

NAND2x1p5_ASAP7_75t_L g976 ( 
.A(n_938),
.B(n_959),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_934),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_923),
.B(n_649),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_950),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_936),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_918),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_936),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_922),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_940),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_928),
.Y(n_985)
);

OAI221xp5_ASAP7_75t_L g986 ( 
.A1(n_931),
.A2(n_730),
.B1(n_747),
.B2(n_715),
.C(n_710),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_925),
.B(n_693),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_932),
.B(n_751),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_932),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_926),
.Y(n_990)
);

OA22x2_ASAP7_75t_L g991 ( 
.A1(n_946),
.A2(n_613),
.B1(n_620),
.B2(n_611),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_945),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_L g993 ( 
.A(n_949),
.B(n_630),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_947),
.B(n_693),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_939),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_953),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_927),
.B(n_776),
.Y(n_997)
);

AO22x2_ASAP7_75t_L g998 ( 
.A1(n_948),
.A2(n_815),
.B1(n_768),
.B2(n_646),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_955),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_929),
.Y(n_1000)
);

OAI221xp5_ASAP7_75t_L g1001 ( 
.A1(n_954),
.A2(n_614),
.B1(n_761),
.B2(n_661),
.C(n_647),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_949),
.Y(n_1002)
);

AO22x2_ASAP7_75t_L g1003 ( 
.A1(n_937),
.A2(n_800),
.B1(n_845),
.B2(n_774),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_926),
.B(n_788),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_926),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_930),
.B(n_791),
.Y(n_1006)
);

BUFx8_ASAP7_75t_L g1007 ( 
.A(n_925),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_931),
.A2(n_731),
.B1(n_764),
.B2(n_728),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_941),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_941),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_930),
.B(n_814),
.Y(n_1011)
);

NAND2x1p5_ASAP7_75t_L g1012 ( 
.A(n_938),
.B(n_632),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_944),
.B(n_639),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_930),
.B(n_712),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_941),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_944),
.B(n_654),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_941),
.Y(n_1017)
);

NOR2xp67_ASAP7_75t_L g1018 ( 
.A(n_959),
.B(n_631),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_941),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_921),
.Y(n_1020)
);

AO22x2_ASAP7_75t_L g1021 ( 
.A1(n_919),
.A2(n_660),
.B1(n_664),
.B2(n_657),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_941),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_944),
.B(n_665),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_931),
.A2(n_640),
.B1(n_659),
.B2(n_653),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_944),
.B(n_674),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_941),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_941),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_930),
.B(n_852),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_944),
.B(n_675),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_944),
.B(n_690),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_930),
.B(n_712),
.Y(n_1031)
);

AO22x2_ASAP7_75t_L g1032 ( 
.A1(n_919),
.A2(n_698),
.B1(n_700),
.B2(n_697),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_941),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_920),
.B(n_705),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_952),
.B(n_809),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_931),
.A2(n_663),
.B1(n_671),
.B2(n_667),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_941),
.Y(n_1037)
);

OAI221xp5_ASAP7_75t_L g1038 ( 
.A1(n_931),
.A2(n_853),
.B1(n_843),
.B2(n_802),
.C(n_762),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_941),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_920),
.B(n_727),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_941),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_921),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_941),
.Y(n_1043)
);

AO22x2_ASAP7_75t_L g1044 ( 
.A1(n_919),
.A2(n_782),
.B1(n_822),
.B2(n_811),
.Y(n_1044)
);

OAI221xp5_ASAP7_75t_L g1045 ( 
.A1(n_931),
.A2(n_833),
.B1(n_834),
.B2(n_813),
.C(n_804),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_920),
.B(n_836),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_941),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_1000),
.B(n_995),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_999),
.B(n_799),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_979),
.B(n_680),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_1011),
.B(n_683),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_SL g1052 ( 
.A(n_994),
.B(n_997),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_983),
.B(n_823),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1002),
.B(n_688),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_992),
.B(n_691),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_964),
.B(n_716),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_1014),
.B(n_695),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_1031),
.B(n_699),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_969),
.B(n_703),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_973),
.B(n_704),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_960),
.B(n_709),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_963),
.B(n_720),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_967),
.B(n_734),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_970),
.B(n_736),
.Y(n_1064)
);

NAND2xp33_ASAP7_75t_SL g1065 ( 
.A(n_990),
.B(n_608),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1013),
.B(n_740),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_1015),
.B(n_741),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_1017),
.B(n_1019),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_1022),
.B(n_743),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_980),
.B(n_326),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_1026),
.B(n_745),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_SL g1073 ( 
.A(n_990),
.B(n_609),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_1027),
.B(n_748),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_1033),
.B(n_750),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_1037),
.B(n_752),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_1039),
.B(n_754),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_1041),
.B(n_755),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_1043),
.B(n_758),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_1047),
.B(n_763),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_1006),
.B(n_767),
.Y(n_1081)
);

NAND2xp33_ASAP7_75t_SL g1082 ( 
.A(n_987),
.B(n_625),
.Y(n_1082)
);

NAND2xp33_ASAP7_75t_SL g1083 ( 
.A(n_1004),
.B(n_673),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_977),
.B(n_769),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_982),
.B(n_772),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_1016),
.B(n_773),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1023),
.B(n_777),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1025),
.B(n_780),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_981),
.B(n_716),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1029),
.B(n_784),
.Y(n_1090)
);

NAND2xp33_ASAP7_75t_SL g1091 ( 
.A(n_1028),
.B(n_725),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1030),
.B(n_786),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_1018),
.B(n_787),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_962),
.B(n_792),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1020),
.B(n_795),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_996),
.B(n_972),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_1034),
.B(n_328),
.Y(n_1097)
);

NAND2xp33_ASAP7_75t_SL g1098 ( 
.A(n_1040),
.B(n_738),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_976),
.B(n_807),
.Y(n_1099)
);

NAND2xp33_ASAP7_75t_SL g1100 ( 
.A(n_1046),
.B(n_789),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1024),
.B(n_816),
.Y(n_1101)
);

NAND2xp33_ASAP7_75t_SL g1102 ( 
.A(n_985),
.B(n_803),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_1036),
.B(n_819),
.Y(n_1103)
);

NAND2xp33_ASAP7_75t_SL g1104 ( 
.A(n_989),
.B(n_827),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_1042),
.B(n_820),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_975),
.B(n_826),
.Y(n_1106)
);

NAND2xp33_ASAP7_75t_SL g1107 ( 
.A(n_966),
.B(n_961),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1044),
.B(n_828),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1008),
.B(n_831),
.Y(n_1109)
);

NAND2xp33_ASAP7_75t_SL g1110 ( 
.A(n_978),
.B(n_842),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_988),
.B(n_835),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1021),
.B(n_837),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_991),
.B(n_844),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_1012),
.B(n_854),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1005),
.B(n_856),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_SL g1116 ( 
.A(n_1032),
.B(n_857),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1007),
.B(n_618),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_984),
.B(n_618),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_965),
.B(n_684),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_1003),
.B(n_684),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_993),
.B(n_666),
.Y(n_1121)
);

NAND2xp33_ASAP7_75t_SL g1122 ( 
.A(n_971),
.B(n_623),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_1038),
.B(n_696),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1045),
.B(n_696),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_974),
.B(n_696),
.Y(n_1125)
);

NAND2xp33_ASAP7_75t_SL g1126 ( 
.A(n_986),
.B(n_627),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_1035),
.B(n_756),
.Y(n_1127)
);

NAND2xp33_ASAP7_75t_SL g1128 ( 
.A(n_1035),
.B(n_628),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1001),
.B(n_634),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_968),
.B(n_676),
.Y(n_1130)
);

NAND2xp33_ASAP7_75t_SL g1131 ( 
.A(n_998),
.B(n_635),
.Y(n_1131)
);

NAND2xp33_ASAP7_75t_SL g1132 ( 
.A(n_1000),
.B(n_641),
.Y(n_1132)
);

NAND2xp33_ASAP7_75t_SL g1133 ( 
.A(n_1000),
.B(n_644),
.Y(n_1133)
);

NAND2xp33_ASAP7_75t_SL g1134 ( 
.A(n_1000),
.B(n_645),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_SL g1135 ( 
.A(n_1000),
.B(n_651),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1000),
.B(n_756),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1000),
.B(n_779),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1000),
.B(n_851),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1000),
.B(n_851),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1000),
.B(n_812),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1000),
.B(n_818),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1000),
.B(n_818),
.Y(n_1142)
);

NAND2xp33_ASAP7_75t_SL g1143 ( 
.A(n_1000),
.B(n_658),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1000),
.B(n_829),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1000),
.B(n_829),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_995),
.B(n_621),
.Y(n_1146)
);

NAND2xp33_ASAP7_75t_SL g1147 ( 
.A(n_1000),
.B(n_668),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1000),
.B(n_678),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_995),
.B(n_679),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1000),
.B(n_685),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_995),
.B(n_702),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1000),
.B(n_707),
.Y(n_1152)
);

NAND2xp33_ASAP7_75t_SL g1153 ( 
.A(n_1000),
.B(n_711),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1000),
.B(n_713),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_995),
.B(n_714),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_995),
.B(n_718),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1000),
.B(n_721),
.Y(n_1157)
);

NAND2xp33_ASAP7_75t_SL g1158 ( 
.A(n_1000),
.B(n_729),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1000),
.B(n_737),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_SL g1160 ( 
.A(n_1000),
.B(n_739),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1000),
.B(n_744),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1000),
.B(n_746),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1000),
.B(n_749),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1000),
.B(n_757),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1000),
.B(n_759),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1000),
.B(n_760),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1000),
.B(n_765),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1000),
.B(n_766),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_995),
.B(n_770),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_995),
.B(n_775),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1000),
.B(n_778),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1053),
.B(n_781),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_SL g1173 ( 
.A(n_1056),
.B(n_794),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1049),
.B(n_783),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1048),
.B(n_801),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1149),
.B(n_805),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1151),
.B(n_806),
.Y(n_1177)
);

INVx3_ASAP7_75t_SL g1178 ( 
.A(n_1117),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_1089),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1066),
.A2(n_331),
.B(n_329),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1121),
.A2(n_333),
.B(n_332),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1069),
.A2(n_335),
.B(n_334),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_SL g1183 ( 
.A1(n_1054),
.A2(n_337),
.B(n_336),
.Y(n_1183)
);

NAND3x1_ASAP7_75t_L g1184 ( 
.A(n_1146),
.B(n_796),
.C(n_794),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1155),
.B(n_1169),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1156),
.B(n_808),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1096),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1071),
.Y(n_1188)
);

INVxp67_ASAP7_75t_L g1189 ( 
.A(n_1113),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1071),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1170),
.B(n_810),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1055),
.A2(n_840),
.B(n_821),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1120),
.A2(n_848),
.B(n_847),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1059),
.A2(n_343),
.B(n_341),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1052),
.A2(n_849),
.B1(n_855),
.B2(n_850),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1067),
.B(n_2),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1082),
.B(n_1051),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1084),
.A2(n_346),
.B(n_345),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1097),
.B(n_796),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_1102),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1105),
.A2(n_1095),
.B(n_1094),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1087),
.A2(n_348),
.B(n_347),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1090),
.A2(n_350),
.B(n_349),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1061),
.A2(n_352),
.B(n_351),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1057),
.B(n_1058),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1129),
.A2(n_1103),
.B(n_1101),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1091),
.B(n_3),
.Y(n_1207)
);

AO21x1_ASAP7_75t_L g1208 ( 
.A1(n_1119),
.A2(n_3),
.B(n_4),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1112),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1130),
.B(n_4),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1081),
.B(n_5),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1099),
.A2(n_1115),
.B(n_1106),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1085),
.A2(n_355),
.B(n_353),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1140),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1141),
.Y(n_1215)
);

BUFx2_ASAP7_75t_R g1216 ( 
.A(n_1125),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1111),
.B(n_356),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1086),
.B(n_1088),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1092),
.A2(n_359),
.B(n_357),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1116),
.A2(n_361),
.B1(n_362),
.B2(n_360),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1062),
.B(n_6),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1142),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1144),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1108),
.A2(n_8),
.A3(n_6),
.B(n_7),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1145),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1107),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1098),
.B(n_365),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1065),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1063),
.A2(n_367),
.B1(n_368),
.B2(n_366),
.Y(n_1229)
);

AND2x2_ASAP7_75t_SL g1230 ( 
.A(n_1083),
.B(n_8),
.Y(n_1230)
);

AOI221x1_ASAP7_75t_L g1231 ( 
.A1(n_1122),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.C(n_12),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1064),
.A2(n_371),
.B(n_370),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1068),
.A2(n_1070),
.B1(n_1074),
.B2(n_1072),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1060),
.B(n_1050),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1075),
.B(n_9),
.Y(n_1235)
);

AO21x2_ASAP7_75t_L g1236 ( 
.A1(n_1093),
.A2(n_375),
.B(n_373),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1148),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1073),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1076),
.B(n_10),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1126),
.A2(n_14),
.A3(n_11),
.B(n_13),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1136),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1077),
.A2(n_377),
.B(n_376),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_SL g1243 ( 
.A1(n_1150),
.A2(n_14),
.B(n_15),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1078),
.A2(n_379),
.B1(n_380),
.B2(n_378),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1079),
.A2(n_382),
.B(n_381),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1080),
.B(n_16),
.Y(n_1246)
);

AOI21xp33_ASAP7_75t_L g1247 ( 
.A1(n_1152),
.A2(n_16),
.B(n_17),
.Y(n_1247)
);

O2A1O1Ixp5_ASAP7_75t_L g1248 ( 
.A1(n_1137),
.A2(n_1138),
.B(n_1139),
.C(n_1109),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_SL g1249 ( 
.A1(n_1118),
.A2(n_386),
.B(n_385),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1132),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1154),
.A2(n_390),
.B1(n_392),
.B2(n_389),
.Y(n_1251)
);

INVx3_ASAP7_75t_SL g1252 ( 
.A(n_1157),
.Y(n_1252)
);

CKINVDCx11_ASAP7_75t_R g1253 ( 
.A(n_1100),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1133),
.A2(n_22),
.B(n_18),
.C(n_21),
.Y(n_1254)
);

AOI21x1_ASAP7_75t_SL g1255 ( 
.A1(n_1131),
.A2(n_21),
.B(n_22),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1159),
.A2(n_395),
.B(n_394),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1114),
.A2(n_398),
.B(n_396),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1161),
.B(n_23),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1162),
.B(n_24),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1110),
.B(n_402),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1163),
.A2(n_405),
.B(n_403),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1207),
.A2(n_1104),
.B1(n_1165),
.B2(n_1164),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1201),
.A2(n_1124),
.B(n_1123),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1188),
.B(n_1166),
.Y(n_1264)
);

CKINVDCx11_ASAP7_75t_R g1265 ( 
.A(n_1253),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1190),
.B(n_1167),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_SL g1267 ( 
.A1(n_1206),
.A2(n_1168),
.B(n_1171),
.C(n_1127),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1185),
.A2(n_1135),
.B(n_1134),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1242),
.A2(n_1158),
.B(n_1153),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1198),
.A2(n_1160),
.B(n_1147),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1226),
.Y(n_1271)
);

OR2x6_ASAP7_75t_L g1272 ( 
.A(n_1212),
.B(n_1128),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1176),
.B(n_1143),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1213),
.A2(n_1257),
.B(n_1181),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1230),
.B(n_25),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1187),
.B(n_407),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1248),
.A2(n_409),
.B(n_408),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1197),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1278)
);

AOI21xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1252),
.A2(n_26),
.B(n_27),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1177),
.B(n_28),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1260),
.B(n_411),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1218),
.A2(n_412),
.B(n_410),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1209),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1189),
.Y(n_1284)
);

AO21x2_ASAP7_75t_L g1285 ( 
.A1(n_1183),
.A2(n_416),
.B(n_414),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1208),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1178),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1231),
.A2(n_418),
.A3(n_419),
.B(n_417),
.Y(n_1288)
);

AO21x2_ASAP7_75t_L g1289 ( 
.A1(n_1196),
.A2(n_424),
.B(n_421),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1194),
.A2(n_427),
.B(n_425),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1219),
.A2(n_429),
.B(n_428),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1186),
.B(n_1191),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1261),
.A2(n_432),
.B(n_431),
.Y(n_1293)
);

NAND2x1p5_ASAP7_75t_L g1294 ( 
.A(n_1237),
.B(n_1227),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1228),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_SL g1296 ( 
.A1(n_1256),
.A2(n_434),
.B(n_435),
.C(n_433),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1233),
.A2(n_442),
.A3(n_443),
.B(n_438),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1202),
.A2(n_446),
.B(n_445),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1238),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1234),
.Y(n_1300)
);

INVx3_ASAP7_75t_L g1301 ( 
.A(n_1234),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1223),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1203),
.A2(n_448),
.B(n_447),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1255),
.A2(n_450),
.B(n_449),
.Y(n_1304)
);

INVxp33_ASAP7_75t_L g1305 ( 
.A(n_1175),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1200),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1172),
.A2(n_452),
.B(n_451),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1214),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1249),
.A2(n_454),
.B(n_453),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1215),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1174),
.B(n_37),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1250),
.A2(n_458),
.A3(n_459),
.B(n_457),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1225),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1217),
.Y(n_1314)
);

AOI22x1_ASAP7_75t_L g1315 ( 
.A1(n_1241),
.A2(n_461),
.B1(n_462),
.B2(n_460),
.Y(n_1315)
);

OR2x6_ASAP7_75t_L g1316 ( 
.A(n_1199),
.B(n_463),
.Y(n_1316)
);

NAND2x1p5_ASAP7_75t_L g1317 ( 
.A(n_1205),
.B(n_464),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1180),
.A2(n_466),
.B(n_465),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1222),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1254),
.A2(n_469),
.A3(n_470),
.B(n_467),
.Y(n_1320)
);

OR2x6_ASAP7_75t_L g1321 ( 
.A(n_1243),
.B(n_471),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1192),
.B(n_38),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1210),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1229),
.A2(n_1244),
.A3(n_1251),
.B(n_1182),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1204),
.A2(n_473),
.B(n_472),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1232),
.A2(n_475),
.B(n_474),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1245),
.A2(n_478),
.B(n_476),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1211),
.Y(n_1328)
);

INVxp67_ASAP7_75t_SL g1329 ( 
.A(n_1258),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1193),
.B(n_1259),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1221),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1216),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1195),
.B(n_39),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1235),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1247),
.A2(n_1239),
.B1(n_1246),
.B2(n_1220),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1240),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1236),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1184),
.A2(n_480),
.B(n_479),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_SL g1339 ( 
.A1(n_1240),
.A2(n_482),
.B(n_481),
.Y(n_1339)
);

NAND2x1p5_ASAP7_75t_L g1340 ( 
.A(n_1240),
.B(n_488),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1224),
.A2(n_484),
.B(n_483),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1224),
.A2(n_486),
.B(n_485),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1188),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1201),
.A2(n_489),
.B(n_487),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1179),
.Y(n_1345)
);

NAND2x1p5_ASAP7_75t_L g1346 ( 
.A(n_1226),
.B(n_493),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_SL g1347 ( 
.A1(n_1206),
.A2(n_492),
.B(n_494),
.C(n_491),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1201),
.A2(n_496),
.B(n_495),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1179),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1201),
.A2(n_500),
.B(n_497),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1179),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1206),
.A2(n_503),
.B(n_501),
.Y(n_1352)
);

OAI221xp5_ASAP7_75t_L g1353 ( 
.A1(n_1173),
.A2(n_44),
.B1(n_41),
.B2(n_43),
.C(n_47),
.Y(n_1353)
);

OAI211xp5_ASAP7_75t_L g1354 ( 
.A1(n_1207),
.A2(n_48),
.B(n_44),
.C(n_47),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1201),
.A2(n_508),
.B(n_507),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1302),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1345),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1308),
.Y(n_1358)
);

BUFx12f_ASAP7_75t_L g1359 ( 
.A(n_1265),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1349),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_SL g1361 ( 
.A(n_1295),
.B(n_509),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1287),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1313),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1351),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1301),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1287),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1322),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1274),
.A2(n_512),
.B(n_510),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1292),
.B(n_51),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1310),
.Y(n_1370)
);

AO21x2_ASAP7_75t_L g1371 ( 
.A1(n_1277),
.A2(n_514),
.B(n_513),
.Y(n_1371)
);

OR2x6_ASAP7_75t_L g1372 ( 
.A(n_1300),
.B(n_516),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1305),
.A2(n_55),
.B1(n_52),
.B2(n_53),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1335),
.A2(n_1280),
.B(n_1329),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1275),
.B(n_1331),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1333),
.B(n_1328),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1314),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1319),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1344),
.A2(n_1350),
.B(n_1348),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1334),
.B(n_52),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1264),
.B(n_517),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1343),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1284),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1266),
.Y(n_1384)
);

AOI211xp5_ASAP7_75t_L g1385 ( 
.A1(n_1353),
.A2(n_56),
.B(n_53),
.C(n_55),
.Y(n_1385)
);

AND2x6_ASAP7_75t_L g1386 ( 
.A(n_1286),
.B(n_1323),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1271),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1336),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1294),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1340),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1311),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1276),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1332),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1321),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1316),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1330),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1297),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1268),
.A2(n_57),
.B(n_58),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1355),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1312),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1263),
.A2(n_519),
.B(n_518),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1272),
.B(n_520),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1341),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1288),
.Y(n_1404)
);

INVx5_ASAP7_75t_L g1405 ( 
.A(n_1272),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1283),
.B(n_1321),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1317),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1299),
.B(n_59),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1262),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1346),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1278),
.B(n_60),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1312),
.Y(n_1412)
);

INVx8_ASAP7_75t_L g1413 ( 
.A(n_1359),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1375),
.B(n_1338),
.Y(n_1414)
);

NAND2xp33_ASAP7_75t_R g1415 ( 
.A(n_1395),
.B(n_1273),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1362),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1376),
.B(n_1297),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1360),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1407),
.B(n_1320),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_R g1420 ( 
.A(n_1361),
.B(n_1337),
.Y(n_1420)
);

BUFx10_ASAP7_75t_L g1421 ( 
.A(n_1393),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1391),
.B(n_1267),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1383),
.B(n_1320),
.Y(n_1423)
);

XNOR2xp5_ASAP7_75t_L g1424 ( 
.A(n_1384),
.B(n_1354),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1374),
.B(n_1307),
.Y(n_1425)
);

BUFx10_ASAP7_75t_L g1426 ( 
.A(n_1381),
.Y(n_1426)
);

XOR2xp5_ASAP7_75t_L g1427 ( 
.A(n_1364),
.B(n_1281),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1366),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1388),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1396),
.B(n_1306),
.Y(n_1430)
);

XNOR2xp5_ASAP7_75t_L g1431 ( 
.A(n_1392),
.B(n_1315),
.Y(n_1431)
);

XNOR2xp5_ASAP7_75t_L g1432 ( 
.A(n_1357),
.B(n_1269),
.Y(n_1432)
);

NAND2xp33_ASAP7_75t_R g1433 ( 
.A(n_1402),
.B(n_1291),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1366),
.B(n_1270),
.Y(n_1434)
);

BUFx10_ASAP7_75t_L g1435 ( 
.A(n_1381),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1405),
.B(n_1352),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1369),
.B(n_1279),
.Y(n_1437)
);

NAND2xp33_ASAP7_75t_SL g1438 ( 
.A(n_1394),
.B(n_1293),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_R g1439 ( 
.A(n_1410),
.B(n_521),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1365),
.B(n_1285),
.Y(n_1440)
);

NAND2xp33_ASAP7_75t_R g1441 ( 
.A(n_1365),
.B(n_1342),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1405),
.B(n_1377),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1387),
.Y(n_1443)
);

OR2x6_ASAP7_75t_L g1444 ( 
.A(n_1372),
.B(n_1282),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1405),
.B(n_1309),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1370),
.Y(n_1446)
);

NAND2xp33_ASAP7_75t_R g1447 ( 
.A(n_1411),
.B(n_1304),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1406),
.B(n_1289),
.Y(n_1448)
);

NAND2xp33_ASAP7_75t_R g1449 ( 
.A(n_1380),
.B(n_1290),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1414),
.B(n_1358),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1429),
.Y(n_1451)
);

NOR2xp67_ASAP7_75t_L g1452 ( 
.A(n_1422),
.B(n_1389),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1417),
.B(n_1378),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1446),
.Y(n_1454)
);

AND2x4_ASAP7_75t_SL g1455 ( 
.A(n_1421),
.B(n_1377),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1443),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1423),
.B(n_1390),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1448),
.B(n_1382),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1442),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1432),
.B(n_1404),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1440),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1425),
.A2(n_1398),
.B1(n_1408),
.B2(n_1367),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1416),
.Y(n_1463)
);

INVxp33_ASAP7_75t_L g1464 ( 
.A(n_1427),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1434),
.Y(n_1465)
);

NOR2xp67_ASAP7_75t_L g1466 ( 
.A(n_1431),
.B(n_1390),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1438),
.A2(n_1409),
.B1(n_1373),
.B2(n_1386),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1418),
.B(n_1400),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1419),
.B(n_1400),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1441),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1437),
.B(n_1397),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1428),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1445),
.B(n_1412),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1415),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1430),
.B(n_1356),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1424),
.B(n_1363),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1436),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1426),
.B(n_1403),
.Y(n_1478)
);

AOI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1420),
.A2(n_1385),
.B1(n_1339),
.B2(n_1347),
.C(n_1296),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1435),
.B(n_1372),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1444),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1439),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1447),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1449),
.B(n_1403),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1463),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1458),
.B(n_1371),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1456),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1471),
.Y(n_1488)
);

AND3x2_ASAP7_75t_L g1489 ( 
.A(n_1474),
.B(n_1413),
.C(n_1399),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1464),
.B(n_1482),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1456),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1460),
.B(n_1401),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1461),
.B(n_1379),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1483),
.B(n_1450),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1454),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1477),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1453),
.B(n_1473),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1465),
.B(n_1368),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1457),
.B(n_1298),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1454),
.B(n_1303),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1470),
.B(n_1325),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1459),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1484),
.B(n_1324),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1469),
.B(n_1326),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1476),
.B(n_1324),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1478),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1466),
.B(n_1327),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1475),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1452),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1459),
.Y(n_1510)
);

OAI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1479),
.A2(n_1433),
.B1(n_1318),
.B2(n_66),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1455),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1472),
.Y(n_1513)
);

OAI221xp5_ASAP7_75t_L g1514 ( 
.A1(n_1467),
.A2(n_68),
.B1(n_63),
.B2(n_67),
.C(n_69),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1480),
.Y(n_1515)
);

NAND2x1_ASAP7_75t_L g1516 ( 
.A(n_1477),
.B(n_63),
.Y(n_1516)
);

INVx5_ASAP7_75t_L g1517 ( 
.A(n_1472),
.Y(n_1517)
);

OAI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1462),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.C(n_70),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1468),
.B(n_70),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1451),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1462),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.C(n_74),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1451),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1468),
.B(n_71),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1454),
.Y(n_1524)
);

INVx4_ASAP7_75t_L g1525 ( 
.A(n_1472),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1468),
.B(n_72),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_L g1527 ( 
.A(n_1479),
.B(n_74),
.C(n_75),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1451),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1451),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1481),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1517),
.B(n_77),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1496),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1530),
.B(n_77),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1530),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1508),
.B(n_78),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1488),
.B(n_78),
.Y(n_1536)
);

OR3x2_ASAP7_75t_L g1537 ( 
.A(n_1505),
.B(n_79),
.C(n_80),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1509),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1497),
.B(n_81),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1494),
.B(n_81),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1506),
.B(n_82),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1493),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1520),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1522),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1503),
.B(n_83),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1487),
.B(n_83),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1486),
.B(n_85),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1528),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1529),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1491),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1495),
.B(n_86),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1510),
.B(n_89),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1517),
.B(n_1525),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1524),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1515),
.Y(n_1555)
);

NAND2x1_ASAP7_75t_L g1556 ( 
.A(n_1502),
.B(n_90),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1501),
.B(n_91),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1492),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1500),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1513),
.B(n_91),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1490),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1512),
.B(n_92),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1485),
.B(n_93),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1517),
.B(n_94),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1504),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1519),
.B(n_1523),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1499),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1498),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1526),
.B(n_1507),
.Y(n_1569)
);

AND2x4_ASAP7_75t_SL g1570 ( 
.A(n_1489),
.B(n_522),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1516),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1511),
.B(n_94),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1527),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1518),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1514),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1521),
.B(n_97),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1530),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1488),
.B(n_97),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1530),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1496),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1508),
.B(n_98),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1496),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1508),
.B(n_98),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1530),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1508),
.B(n_99),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1488),
.B(n_99),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1488),
.B(n_100),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1530),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1497),
.B(n_100),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1496),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1530),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1497),
.B(n_102),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1538),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1547),
.B(n_103),
.Y(n_1594)
);

NAND2xp33_ASAP7_75t_R g1595 ( 
.A(n_1564),
.B(n_104),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1552),
.Y(n_1596)
);

NAND2xp33_ASAP7_75t_R g1597 ( 
.A(n_1564),
.B(n_1533),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1571),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1574),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1573),
.A2(n_108),
.B1(n_105),
.B2(n_107),
.C(n_109),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1572),
.A2(n_1575),
.B1(n_1576),
.B2(n_1545),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1569),
.Y(n_1602)
);

AO221x2_ASAP7_75t_L g1603 ( 
.A1(n_1537),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.C(n_112),
.Y(n_1603)
);

NOR2x1_ASAP7_75t_L g1604 ( 
.A(n_1553),
.B(n_1533),
.Y(n_1604)
);

XNOR2xp5_ASAP7_75t_L g1605 ( 
.A(n_1566),
.B(n_1539),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1565),
.B(n_112),
.Y(n_1606)
);

AO221x2_ASAP7_75t_L g1607 ( 
.A1(n_1557),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.C(n_116),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1532),
.B(n_114),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1552),
.Y(n_1609)
);

NOR2x1_ASAP7_75t_L g1610 ( 
.A(n_1531),
.B(n_1535),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1580),
.B(n_1582),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1590),
.B(n_117),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1534),
.Y(n_1613)
);

NOR2x1_ASAP7_75t_L g1614 ( 
.A(n_1581),
.B(n_1583),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1548),
.B(n_118),
.Y(n_1615)
);

OAI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1567),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1542),
.B(n_121),
.Y(n_1617)
);

AO221x2_ASAP7_75t_L g1618 ( 
.A1(n_1551),
.A2(n_125),
.B1(n_122),
.B2(n_124),
.C(n_126),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1570),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1549),
.B(n_127),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1554),
.B(n_128),
.Y(n_1621)
);

AO221x2_ASAP7_75t_L g1622 ( 
.A1(n_1540),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.C(n_131),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1585),
.B(n_129),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1536),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1568),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_1625)
);

NOR2x1_ASAP7_75t_L g1626 ( 
.A(n_1578),
.B(n_1586),
.Y(n_1626)
);

OAI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1587),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1543),
.B(n_134),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1577),
.B(n_136),
.Y(n_1629)
);

AO221x2_ASAP7_75t_L g1630 ( 
.A1(n_1579),
.A2(n_140),
.B1(n_137),
.B2(n_139),
.C(n_142),
.Y(n_1630)
);

CKINVDCx20_ASAP7_75t_R g1631 ( 
.A(n_1589),
.Y(n_1631)
);

OAI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1584),
.A2(n_1588),
.B1(n_1591),
.B2(n_1559),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1544),
.B(n_143),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1550),
.B(n_1541),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1546),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1546),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1560),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1592),
.B(n_149),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1563),
.B(n_150),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_R g1640 ( 
.A(n_1562),
.B(n_150),
.Y(n_1640)
);

NOR4xp25_ASAP7_75t_SL g1641 ( 
.A(n_1553),
.B(n_153),
.C(n_151),
.D(n_152),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1561),
.B(n_154),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1561),
.B(n_155),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1555),
.B(n_156),
.Y(n_1644)
);

AND2x4_ASAP7_75t_SL g1645 ( 
.A(n_1552),
.B(n_158),
.Y(n_1645)
);

NAND2xp33_ASAP7_75t_SL g1646 ( 
.A(n_1556),
.B(n_159),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1555),
.B(n_160),
.Y(n_1647)
);

CKINVDCx16_ASAP7_75t_R g1648 ( 
.A(n_1552),
.Y(n_1648)
);

NAND2xp33_ASAP7_75t_SL g1649 ( 
.A(n_1556),
.B(n_160),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1561),
.B(n_161),
.Y(n_1650)
);

NAND2xp33_ASAP7_75t_SL g1651 ( 
.A(n_1556),
.B(n_161),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1574),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_1652)
);

OAI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1573),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.C(n_165),
.Y(n_1653)
);

NOR2x1_ASAP7_75t_L g1654 ( 
.A(n_1553),
.B(n_166),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1555),
.B(n_167),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1563),
.Y(n_1656)
);

NOR2x1_ASAP7_75t_L g1657 ( 
.A(n_1553),
.B(n_168),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1558),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1555),
.B(n_169),
.Y(n_1659)
);

OAI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1573),
.A2(n_173),
.B1(n_170),
.B2(n_172),
.Y(n_1660)
);

NAND2xp33_ASAP7_75t_SL g1661 ( 
.A(n_1556),
.B(n_173),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1555),
.B(n_174),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1598),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1614),
.B(n_175),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1603),
.A2(n_176),
.B(n_177),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1640),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1595),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1593),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1602),
.B(n_178),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1611),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1624),
.B(n_179),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1626),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1628),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1633),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1620),
.Y(n_1675)
);

OR2x6_ASAP7_75t_L g1676 ( 
.A(n_1654),
.B(n_180),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1596),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1609),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1613),
.Y(n_1679)
);

OR2x6_ASAP7_75t_L g1680 ( 
.A(n_1657),
.B(n_181),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1635),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1656),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1617),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1634),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1608),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1629),
.B(n_182),
.Y(n_1686)
);

OAI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1599),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.C(n_185),
.Y(n_1687)
);

CKINVDCx16_ASAP7_75t_R g1688 ( 
.A(n_1597),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1605),
.B(n_187),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1610),
.B(n_188),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1631),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1655),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1644),
.B(n_1647),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1612),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1645),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1659),
.B(n_189),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1662),
.B(n_189),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1621),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1601),
.B(n_190),
.Y(n_1699)
);

AO21x2_ASAP7_75t_L g1700 ( 
.A1(n_1615),
.A2(n_190),
.B(n_191),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1594),
.B(n_1623),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1632),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1630),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1639),
.B(n_192),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1638),
.B(n_193),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1642),
.B(n_194),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1643),
.B(n_196),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1650),
.B(n_198),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1606),
.B(n_200),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1600),
.B(n_203),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1618),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1607),
.B(n_203),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1652),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1607),
.B(n_207),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1646),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1622),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1649),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1636),
.B(n_207),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1625),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1637),
.B(n_208),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1651),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1627),
.Y(n_1722)
);

NAND3x1_ASAP7_75t_L g1723 ( 
.A(n_1619),
.B(n_1661),
.C(n_1641),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1616),
.B(n_211),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1660),
.B(n_212),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1653),
.B(n_212),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1604),
.B(n_213),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1595),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1640),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1640),
.Y(n_1730)
);

AOI222xp33_ASAP7_75t_L g1731 ( 
.A1(n_1600),
.A2(n_216),
.B1(n_219),
.B2(n_214),
.C1(n_215),
.C2(n_217),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1598),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1604),
.B(n_215),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1611),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1658),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1602),
.B(n_216),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1611),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1604),
.B(n_220),
.Y(n_1738)
);

AND3x1_ASAP7_75t_L g1739 ( 
.A(n_1604),
.B(n_220),
.C(n_221),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1611),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1602),
.B(n_221),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1640),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1624),
.B(n_222),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1598),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1598),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1648),
.A2(n_227),
.B1(n_224),
.B2(n_226),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1658),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1602),
.B(n_228),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1648),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1640),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1604),
.B(n_228),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1604),
.B(n_229),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1598),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1595),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1598),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1640),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1598),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1604),
.B(n_230),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1604),
.B(n_230),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1598),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1602),
.B(n_231),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1611),
.Y(n_1762)
);

NAND2x1_ASAP7_75t_SL g1763 ( 
.A(n_1604),
.B(n_232),
.Y(n_1763)
);

BUFx3_ASAP7_75t_L g1764 ( 
.A(n_1596),
.Y(n_1764)
);

O2A1O1Ixp5_ASAP7_75t_L g1765 ( 
.A1(n_1703),
.A2(n_239),
.B(n_237),
.C(n_238),
.Y(n_1765)
);

AOI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1665),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1688),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_1767)
);

NOR2x1_ASAP7_75t_L g1768 ( 
.A(n_1738),
.B(n_245),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1735),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1747),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1672),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.C(n_251),
.Y(n_1771)
);

O2A1O1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1667),
.A2(n_252),
.B(n_250),
.C(n_251),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1728),
.B(n_252),
.Y(n_1773)
);

INVx1_ASAP7_75t_SL g1774 ( 
.A(n_1763),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1749),
.Y(n_1775)
);

OAI32xp33_ASAP7_75t_L g1776 ( 
.A1(n_1716),
.A2(n_255),
.A3(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1738),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1739),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1677),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1723),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1759),
.B(n_258),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1666),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1683),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1681),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1682),
.B(n_1679),
.Y(n_1785)
);

AOI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1699),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.C(n_263),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1711),
.B(n_262),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1691),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_SL g1789 ( 
.A(n_1754),
.B(n_263),
.Y(n_1789)
);

O2A1O1Ixp33_ASAP7_75t_L g1790 ( 
.A1(n_1712),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_1790)
);

AO211x2_ASAP7_75t_L g1791 ( 
.A1(n_1702),
.A2(n_267),
.B(n_264),
.C(n_266),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1670),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1692),
.B(n_268),
.Y(n_1793)
);

AOI322xp5_ASAP7_75t_L g1794 ( 
.A1(n_1714),
.A2(n_268),
.A3(n_269),
.B1(n_270),
.B2(n_271),
.C1(n_272),
.C2(n_273),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1684),
.B(n_269),
.Y(n_1795)
);

OAI31xp33_ASAP7_75t_L g1796 ( 
.A1(n_1715),
.A2(n_277),
.A3(n_275),
.B(n_276),
.Y(n_1796)
);

AOI21xp33_ASAP7_75t_L g1797 ( 
.A1(n_1710),
.A2(n_275),
.B(n_276),
.Y(n_1797)
);

OAI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1717),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1719),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_1799)
);

AND2x4_ASAP7_75t_SL g1800 ( 
.A(n_1676),
.B(n_1680),
.Y(n_1800)
);

NOR3xp33_ASAP7_75t_L g1801 ( 
.A(n_1687),
.B(n_281),
.C(n_282),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1734),
.Y(n_1802)
);

INVxp67_ASAP7_75t_L g1803 ( 
.A(n_1721),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1737),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1740),
.Y(n_1805)
);

INVxp67_ASAP7_75t_L g1806 ( 
.A(n_1727),
.Y(n_1806)
);

O2A1O1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1676),
.A2(n_285),
.B(n_283),
.C(n_284),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1725),
.A2(n_286),
.B(n_289),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1663),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1722),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1732),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1685),
.B(n_294),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1733),
.B(n_296),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1744),
.Y(n_1814)
);

AOI31xp33_ASAP7_75t_L g1815 ( 
.A1(n_1729),
.A2(n_299),
.A3(n_297),
.B(n_298),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1713),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1730),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1745),
.B(n_305),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1753),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1742),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1755),
.Y(n_1821)
);

INVxp67_ASAP7_75t_L g1822 ( 
.A(n_1751),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1752),
.B(n_1758),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1757),
.B(n_307),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1762),
.Y(n_1825)
);

OAI32xp33_ASAP7_75t_L g1826 ( 
.A1(n_1726),
.A2(n_309),
.A3(n_307),
.B1(n_308),
.B2(n_310),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1731),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1694),
.B(n_311),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1680),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1675),
.B(n_313),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1673),
.B(n_314),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1674),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1760),
.B(n_314),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1668),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1690),
.B(n_315),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1750),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1669),
.Y(n_1837)
);

NOR2xp67_ASAP7_75t_L g1838 ( 
.A(n_1664),
.B(n_317),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1698),
.B(n_1678),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1764),
.B(n_318),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1780),
.B(n_1700),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1777),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1788),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1782),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1783),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1769),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1774),
.B(n_1779),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1770),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1800),
.A2(n_1718),
.B1(n_1689),
.B2(n_1709),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1784),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1803),
.B(n_1701),
.Y(n_1851)
);

CKINVDCx16_ASAP7_75t_R g1852 ( 
.A(n_1789),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1837),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1766),
.A2(n_1718),
.B1(n_1724),
.B2(n_1756),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1834),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1775),
.B(n_1695),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1839),
.B(n_1696),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1817),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1785),
.B(n_1697),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1820),
.B(n_1693),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1836),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1823),
.B(n_1736),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1768),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1832),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1806),
.B(n_1671),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_1793),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1792),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1822),
.B(n_1686),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_SL g1869 ( 
.A1(n_1808),
.A2(n_1720),
.B1(n_1746),
.B2(n_1743),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1802),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1804),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1831),
.B(n_1704),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1805),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1809),
.B(n_1706),
.Y(n_1874)
);

NOR2x1_ASAP7_75t_L g1875 ( 
.A(n_1838),
.B(n_1741),
.Y(n_1875)
);

NOR3xp33_ASAP7_75t_L g1876 ( 
.A(n_1790),
.B(n_1708),
.C(n_1707),
.Y(n_1876)
);

NOR2x1_ASAP7_75t_L g1877 ( 
.A(n_1815),
.B(n_1748),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1819),
.B(n_1811),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1787),
.B(n_1705),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1824),
.B(n_1814),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1821),
.B(n_1761),
.Y(n_1881)
);

INVx2_ASAP7_75t_SL g1882 ( 
.A(n_1840),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1842),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1863),
.Y(n_1884)
);

INVx1_ASAP7_75t_SL g1885 ( 
.A(n_1844),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1852),
.B(n_1773),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1858),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1856),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1845),
.Y(n_1889)
);

INVx8_ASAP7_75t_L g1890 ( 
.A(n_1857),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1846),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1848),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1868),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1850),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1855),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1861),
.Y(n_1896)
);

BUFx4_ASAP7_75t_SL g1897 ( 
.A(n_1853),
.Y(n_1897)
);

INVx1_ASAP7_75t_SL g1898 ( 
.A(n_1875),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1864),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1867),
.Y(n_1900)
);

INVx2_ASAP7_75t_SL g1901 ( 
.A(n_1878),
.Y(n_1901)
);

INVx1_ASAP7_75t_SL g1902 ( 
.A(n_1866),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1870),
.Y(n_1903)
);

O2A1O1Ixp5_ASAP7_75t_SL g1904 ( 
.A1(n_1884),
.A2(n_1847),
.B(n_1873),
.C(n_1871),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1890),
.Y(n_1905)
);

NAND4xp25_ASAP7_75t_SL g1906 ( 
.A(n_1898),
.B(n_1877),
.C(n_1841),
.D(n_1794),
.Y(n_1906)
);

AOI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1896),
.A2(n_1801),
.B1(n_1885),
.B2(n_1886),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1883),
.A2(n_1854),
.B1(n_1767),
.B2(n_1772),
.C(n_1798),
.Y(n_1908)
);

AOI211xp5_ASAP7_75t_L g1909 ( 
.A1(n_1902),
.A2(n_1826),
.B(n_1797),
.C(n_1807),
.Y(n_1909)
);

NOR3xp33_ASAP7_75t_L g1910 ( 
.A(n_1887),
.B(n_1851),
.C(n_1843),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1888),
.B(n_1849),
.Y(n_1911)
);

NOR4xp25_ASAP7_75t_L g1912 ( 
.A(n_1889),
.B(n_1786),
.C(n_1829),
.D(n_1771),
.Y(n_1912)
);

OAI211xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1893),
.A2(n_1869),
.B(n_1796),
.C(n_1876),
.Y(n_1913)
);

NOR3xp33_ASAP7_75t_L g1914 ( 
.A(n_1901),
.B(n_1860),
.C(n_1865),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1890),
.B(n_1859),
.Y(n_1915)
);

OAI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1891),
.A2(n_1765),
.B(n_1778),
.Y(n_1916)
);

OA22x2_ASAP7_75t_L g1917 ( 
.A1(n_1907),
.A2(n_1882),
.B1(n_1880),
.B2(n_1827),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1915),
.B(n_1874),
.Y(n_1918)
);

AOI322xp5_ASAP7_75t_L g1919 ( 
.A1(n_1908),
.A2(n_1879),
.A3(n_1892),
.B1(n_1862),
.B2(n_1872),
.C1(n_1900),
.C2(n_1899),
.Y(n_1919)
);

XNOR2x1_ASAP7_75t_L g1920 ( 
.A(n_1905),
.B(n_1791),
.Y(n_1920)
);

NOR3xp33_ASAP7_75t_L g1921 ( 
.A(n_1906),
.B(n_1895),
.C(n_1894),
.Y(n_1921)
);

XOR2xp5_ASAP7_75t_L g1922 ( 
.A(n_1920),
.B(n_1911),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1918),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1917),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1921),
.Y(n_1925)
);

NAND3xp33_ASAP7_75t_L g1926 ( 
.A(n_1925),
.B(n_1904),
.C(n_1919),
.Y(n_1926)
);

NOR3xp33_ASAP7_75t_SL g1927 ( 
.A(n_1923),
.B(n_1913),
.C(n_1916),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1924),
.B(n_1914),
.Y(n_1928)
);

NAND5xp2_ASAP7_75t_L g1929 ( 
.A(n_1927),
.B(n_1910),
.C(n_1909),
.D(n_1922),
.E(n_1903),
.Y(n_1929)
);

OR3x1_ASAP7_75t_L g1930 ( 
.A(n_1929),
.B(n_1897),
.C(n_1776),
.Y(n_1930)
);

AO21x2_ASAP7_75t_L g1931 ( 
.A1(n_1930),
.A2(n_1926),
.B(n_1928),
.Y(n_1931)
);

AOI31xp33_ASAP7_75t_L g1932 ( 
.A1(n_1931),
.A2(n_1781),
.A3(n_1835),
.B(n_1813),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1932),
.A2(n_1912),
.B1(n_1818),
.B2(n_1833),
.Y(n_1933)
);

AOI21xp33_ASAP7_75t_L g1934 ( 
.A1(n_1933),
.A2(n_1881),
.B(n_1828),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_1934),
.Y(n_1935)
);

OAI221xp5_ASAP7_75t_R g1936 ( 
.A1(n_1935),
.A2(n_1810),
.B1(n_1799),
.B2(n_1816),
.C(n_1812),
.Y(n_1936)
);

OAI31xp33_ASAP7_75t_L g1937 ( 
.A1(n_1936),
.A2(n_1830),
.A3(n_1795),
.B(n_1825),
.Y(n_1937)
);


endmodule