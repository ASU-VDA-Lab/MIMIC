module fake_jpeg_31601_n_491 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_491);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_491;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_53),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_15),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_54),
.B(n_64),
.Y(n_134)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_55),
.Y(n_143)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g118 ( 
.A(n_56),
.Y(n_118)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_61),
.B(n_67),
.Y(n_125)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_49),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_33),
.B(n_17),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_25),
.A2(n_17),
.B1(n_14),
.B2(n_2),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_41),
.B1(n_32),
.B2(n_48),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_31),
.Y(n_73)
);

CKINVDCx6p67_ASAP7_75t_R g148 ( 
.A(n_73),
.Y(n_148)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx2_ASAP7_75t_SL g151 ( 
.A(n_75),
.Y(n_151)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_28),
.B(n_14),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_78),
.B(n_87),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_0),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_0),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_92),
.B(n_96),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

CKINVDCx9p33_ASAP7_75t_R g153 ( 
.A(n_93),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_97),
.Y(n_113)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_23),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_104),
.A2(n_105),
.B1(n_116),
.B2(n_42),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_33),
.B1(n_26),
.B2(n_22),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_30),
.B1(n_20),
.B2(n_46),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_107),
.A2(n_108),
.B1(n_131),
.B2(n_149),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_30),
.B1(n_20),
.B2(n_46),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_30),
.B1(n_47),
.B2(n_21),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_110),
.A2(n_146),
.B1(n_39),
.B2(n_47),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_48),
.B1(n_26),
.B2(n_42),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_46),
.B1(n_32),
.B2(n_41),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_92),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_147),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_64),
.B(n_18),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_142),
.B(n_1),
.C(n_2),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_80),
.A2(n_21),
.B1(n_39),
.B2(n_34),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_75),
.B(n_18),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_94),
.A2(n_32),
.B1(n_41),
.B2(n_21),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_93),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_73),
.B(n_22),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_122),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_157),
.B(n_169),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_100),
.B1(n_84),
.B2(n_43),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_118),
.A2(n_44),
.B1(n_35),
.B2(n_43),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_159),
.A2(n_170),
.B1(n_176),
.B2(n_209),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_44),
.B(n_35),
.C(n_96),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_160),
.B(n_165),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_161),
.A2(n_168),
.B1(n_174),
.B2(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_39),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_162),
.B(n_197),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_164),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_148),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_167),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_141),
.B1(n_110),
.B2(n_146),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_180),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_70),
.B1(n_59),
.B2(n_60),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_134),
.A2(n_24),
.B(n_47),
.C(n_34),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_175),
.B(n_177),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_79),
.B1(n_82),
.B2(n_51),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_34),
.B(n_24),
.C(n_23),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_131),
.A2(n_149),
.B1(n_107),
.B2(n_108),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_179),
.B(n_185),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_114),
.B(n_81),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_113),
.Y(n_185)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_118),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_192),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g212 ( 
.A(n_188),
.B(n_203),
.CI(n_204),
.CON(n_212),
.SN(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_128),
.A2(n_24),
.B(n_23),
.C(n_3),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_189),
.A2(n_123),
.B(n_111),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_117),
.A2(n_69),
.B1(n_65),
.B2(n_90),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_190),
.A2(n_191),
.B1(n_201),
.B2(n_174),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_121),
.A2(n_83),
.B1(n_23),
.B2(n_3),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_124),
.B(n_135),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_194),
.Y(n_235)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_129),
.A2(n_23),
.B(n_4),
.Y(n_196)
);

OR2x6_ASAP7_75t_L g245 ( 
.A(n_196),
.B(n_6),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_119),
.B(n_3),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_136),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_109),
.Y(n_202)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_123),
.B(n_4),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_119),
.B(n_137),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_122),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_103),
.Y(n_206)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_138),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_137),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_210),
.A2(n_213),
.B(n_236),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_163),
.A2(n_126),
.B1(n_103),
.B2(n_136),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_184),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_229),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_160),
.A2(n_120),
.B1(n_130),
.B2(n_126),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_223),
.A2(n_238),
.B1(n_248),
.B2(n_187),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_228),
.A2(n_191),
.B1(n_183),
.B2(n_182),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_181),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_162),
.A2(n_122),
.B(n_101),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_170),
.A2(n_144),
.B1(n_132),
.B2(n_127),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_164),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_165),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_168),
.A2(n_144),
.B1(n_132),
.B2(n_127),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_241),
.A2(n_207),
.B1(n_167),
.B2(n_202),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_178),
.A2(n_138),
.B1(n_115),
.B2(n_9),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_201),
.C(n_197),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_166),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_248)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_185),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_254),
.A2(n_189),
.B(n_177),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_255),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_231),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_278),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_257),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_258),
.A2(n_269),
.B(n_290),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_188),
.C(n_204),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_280),
.C(n_287),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_215),
.A2(n_203),
.B1(n_188),
.B2(n_161),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

OAI21xp33_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_201),
.B(n_191),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_262),
.A2(n_295),
.B(n_255),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_264),
.A2(n_279),
.B1(n_283),
.B2(n_293),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_203),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_267),
.Y(n_329)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_175),
.B(n_171),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_216),
.B(n_191),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_272),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_179),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_212),
.B(n_205),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_275),
.B(n_285),
.Y(n_313)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_210),
.A2(n_190),
.B(n_193),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_276),
.A2(n_286),
.B(n_246),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_231),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_224),
.A2(n_198),
.B1(n_207),
.B2(n_202),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_212),
.B(n_199),
.C(n_157),
.Y(n_280)
);

INVx13_ASAP7_75t_L g281 ( 
.A(n_225),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_281),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_224),
.A2(n_167),
.B1(n_208),
.B2(n_186),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_211),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_289),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_212),
.B(n_11),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_245),
.A2(n_200),
.B(n_195),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_245),
.B(n_236),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_287),
.B(n_288),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_220),
.B(n_11),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_227),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_245),
.A2(n_11),
.B(n_12),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_228),
.B(n_235),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_291),
.Y(n_319)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_225),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_249),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_213),
.A2(n_241),
.B1(n_233),
.B2(n_218),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_219),
.Y(n_294)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_233),
.A2(n_218),
.B(n_222),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_274),
.A2(n_222),
.B(n_221),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_304),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_275),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_306),
.C(n_320),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_221),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_312),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_310),
.A2(n_311),
.B(n_327),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_240),
.B(n_246),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_256),
.B(n_234),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_314),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_249),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_316),
.B(n_322),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_278),
.B(n_261),
.Y(n_317)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_253),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_325),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_285),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_272),
.B(n_234),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_243),
.C(n_239),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_330),
.C(n_289),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_243),
.C(n_239),
.Y(n_330)
);

AND2x2_ASAP7_75t_SL g332 ( 
.A(n_271),
.B(n_214),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_332),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_321),
.A2(n_264),
.B1(n_291),
.B2(n_277),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_335),
.A2(n_340),
.B1(n_351),
.B2(n_355),
.Y(n_367)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_269),
.C(n_260),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_302),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_321),
.A2(n_279),
.B1(n_307),
.B2(n_299),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_341),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_299),
.A2(n_270),
.B1(n_276),
.B2(n_262),
.Y(n_342)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_343),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_286),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_347),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_296),
.A2(n_293),
.B1(n_283),
.B2(n_276),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_346),
.A2(n_350),
.B(n_297),
.Y(n_374)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_306),
.B(n_288),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_359),
.C(n_361),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_276),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_SL g351 ( 
.A(n_301),
.B(n_273),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_301),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_358),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_307),
.A2(n_290),
.B1(n_258),
.B2(n_286),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_294),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_313),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_304),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_318),
.B(n_268),
.C(n_263),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_323),
.Y(n_360)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_360),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_300),
.B(n_263),
.C(n_252),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_331),
.A2(n_282),
.B1(n_227),
.B2(n_251),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_362),
.A2(n_330),
.B1(n_319),
.B2(n_326),
.Y(n_369)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_363),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_339),
.B(n_319),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_368),
.A2(n_328),
.B1(n_313),
.B2(n_332),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_369),
.A2(n_337),
.B1(n_357),
.B2(n_345),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_392),
.Y(n_403)
);

NOR2x1_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_298),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_387),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_374),
.A2(n_376),
.B(n_384),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_353),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_375),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_364),
.A2(n_327),
.B(n_310),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_352),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_377),
.B(n_388),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_341),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_379),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_333),
.A2(n_303),
.B1(n_309),
.B2(n_324),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_381),
.A2(n_389),
.B1(n_334),
.B2(n_332),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_298),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_382),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_364),
.A2(n_311),
.B(n_302),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_336),
.A2(n_327),
.B(n_317),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

INVxp33_ASAP7_75t_SL g387 ( 
.A(n_356),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_322),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_350),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_391),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_366),
.A2(n_346),
.B1(n_336),
.B2(n_362),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_394),
.A2(n_378),
.B1(n_324),
.B2(n_309),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_395),
.B(n_409),
.Y(n_425)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_390),
.Y(n_397)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

XNOR2x1_ASAP7_75t_L g435 ( 
.A(n_399),
.B(n_292),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_344),
.C(n_347),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_408),
.C(n_412),
.Y(n_417)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_390),
.Y(n_404)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_404),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_366),
.A2(n_342),
.B1(n_331),
.B2(n_332),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_405),
.A2(n_373),
.B1(n_380),
.B2(n_385),
.Y(n_428)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_406),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_344),
.C(n_337),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_371),
.B(n_348),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_411),
.Y(n_432)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_365),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_349),
.C(n_359),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_375),
.B(n_360),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_413),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_361),
.C(n_328),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_368),
.C(n_370),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_415),
.B(n_392),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_421),
.Y(n_440)
);

A2O1A1Ixp33_ASAP7_75t_SL g419 ( 
.A1(n_398),
.A2(n_376),
.B(n_386),
.C(n_374),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_419),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_367),
.C(n_369),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_403),
.C(n_414),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_367),
.C(n_384),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_427),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_402),
.B(n_391),
.C(n_385),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_428),
.A2(n_394),
.B1(n_400),
.B2(n_415),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_398),
.B(n_380),
.Y(n_429)
);

A2O1A1O1Ixp25_ASAP7_75t_L g446 ( 
.A1(n_429),
.A2(n_409),
.B(n_411),
.C(n_404),
.D(n_406),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_431),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_401),
.A2(n_378),
.B(n_329),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_433),
.A2(n_401),
.B(n_410),
.Y(n_439)
);

FAx1_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_309),
.CI(n_292),
.CON(n_434),
.SN(n_434)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_434),
.B(n_413),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_435),
.B(n_405),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_439),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_443),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_438),
.B(n_448),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_432),
.B(n_407),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_447),
.Y(n_456)
);

NOR2x1_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_429),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_395),
.C(n_403),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_420),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_423),
.A2(n_393),
.B1(n_396),
.B2(n_397),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_419),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_424),
.A2(n_396),
.B(n_416),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_450),
.A2(n_422),
.B(n_434),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_442),
.A2(n_430),
.B1(n_422),
.B2(n_435),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_281),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_440),
.B(n_417),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_455),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_444),
.B(n_434),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_459),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_462),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_419),
.Y(n_461)
);

AOI31xp67_ASAP7_75t_SL g468 ( 
.A1(n_461),
.A2(n_419),
.A3(n_446),
.B(n_443),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_425),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_441),
.A2(n_447),
.B(n_442),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_463),
.A2(n_425),
.B(n_250),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_456),
.B(n_436),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_466),
.B(n_468),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_453),
.B(n_329),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_472),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_470),
.B(n_471),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_460),
.B(n_453),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_257),
.Y(n_472)
);

AOI322xp5_ASAP7_75t_L g473 ( 
.A1(n_459),
.A2(n_281),
.A3(n_242),
.B1(n_250),
.B2(n_267),
.C1(n_257),
.C2(n_252),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_473),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_474),
.B(n_454),
.C(n_451),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_477),
.B(n_478),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_464),
.C(n_462),
.Y(n_478)
);

A2O1A1O1Ixp25_ASAP7_75t_L g481 ( 
.A1(n_467),
.A2(n_232),
.B(n_454),
.C(n_457),
.D(n_470),
.Y(n_481)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_481),
.Y(n_485)
);

AO21x1_ASAP7_75t_L g482 ( 
.A1(n_476),
.A2(n_474),
.B(n_232),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_482),
.Y(n_487)
);

BUFx24_ASAP7_75t_SL g484 ( 
.A(n_480),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_484),
.A2(n_483),
.B(n_485),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_486),
.B(n_487),
.Y(n_488)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_488),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_486),
.A2(n_475),
.B(n_479),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_489),
.Y(n_491)
);


endmodule