module real_jpeg_29125_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_297, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_297;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_292;
wire n_286;
wire n_288;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_290;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_285;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_55;
wire n_240;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_202;
wire n_295;
wire n_128;
wire n_213;
wire n_179;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_0),
.A2(n_73),
.B1(n_74),
.B2(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_0),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_0),
.A2(n_32),
.B1(n_35),
.B2(n_122),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_122),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_122),
.Y(n_235)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_1),
.Y(n_85)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_2),
.A2(n_46),
.B1(n_73),
.B2(n_74),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_46),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_2),
.A2(n_32),
.B1(n_35),
.B2(n_46),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_3),
.B(n_26),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_25),
.B(n_26),
.C(n_135),
.D(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_3),
.B(n_48),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_3),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_3),
.A2(n_84),
.B(n_152),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_3),
.A2(n_44),
.B(n_47),
.C(n_183),
.D(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_3),
.B(n_44),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_3),
.A2(n_45),
.B(n_71),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_3),
.A2(n_73),
.B1(n_74),
.B2(n_167),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_4),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_4),
.A2(n_32),
.B1(n_35),
.B2(n_147),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_147),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_4),
.A2(n_73),
.B1(n_74),
.B2(n_147),
.Y(n_252)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_7),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_7),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_76),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_7),
.A2(n_32),
.B1(n_35),
.B2(n_76),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_76),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_73),
.B1(n_74),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_8),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_99),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_8),
.A2(n_32),
.B1(n_35),
.B2(n_99),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_99),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_32),
.B1(n_35),
.B2(n_40),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_11),
.A2(n_26),
.B(n_28),
.C(n_31),
.Y(n_25)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_12),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_12),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_111)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_15),
.A2(n_32),
.B1(n_35),
.B2(n_54),
.Y(n_222)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_100),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_20),
.B(n_100),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_81),
.B2(n_82),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_55),
.B1(n_56),
.B2(n_80),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_23),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_23),
.A2(n_24),
.B(n_41),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_36),
.B2(n_38),
.Y(n_24)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_25),
.A2(n_31),
.B1(n_36),
.B2(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_25),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_25),
.A2(n_31),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_26),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_26),
.A2(n_45),
.A3(n_183),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g134 ( 
.A1(n_27),
.A2(n_30),
.A3(n_35),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_27),
.B(n_50),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_29),
.B(n_32),
.Y(n_136)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2x1_ASAP7_75t_SL g84 ( 
.A(n_32),
.B(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_35),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_62),
.B(n_63),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_43),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_45),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_48),
.B1(n_53),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_47),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_47),
.A2(n_48),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_50),
.Y(n_194)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_66),
.B2(n_79),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_63),
.B1(n_94),
.B2(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_62),
.A2(n_211),
.B(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_62),
.A2(n_63),
.B1(n_114),
.B2(n_238),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_63),
.B(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_63),
.A2(n_146),
.B(n_148),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_63),
.B(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_63),
.A2(n_148),
.B(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_67),
.A2(n_120),
.B(n_123),
.Y(n_119)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_68),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_68),
.A2(n_69),
.B1(n_121),
.B2(n_252),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_69),
.B(n_98),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_70),
.A2(n_73),
.B(n_167),
.C(n_225),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_73),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_77),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_77),
.B(n_167),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_77),
.A2(n_97),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_90),
.B(n_95),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_95),
.B1(n_96),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_83),
.A2(n_91),
.B1(n_92),
.B2(n_104),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B(n_89),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_89),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_84),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_84),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_84),
.B(n_154),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_84),
.A2(n_86),
.B1(n_192),
.B2(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_84),
.A2(n_88),
.B1(n_111),
.B2(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_86),
.A2(n_159),
.B(n_169),
.Y(n_168)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_87),
.B(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_87),
.A2(n_170),
.B(n_191),
.Y(n_190)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_88),
.B(n_167),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_103),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.C(n_107),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_284)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_107),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_115),
.C(n_119),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_108),
.A2(n_109),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_110),
.B(n_113),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_115),
.B(n_119),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_116),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_117),
.A2(n_118),
.B(n_202),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_118),
.B(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_118),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_123),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI321xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_276),
.A3(n_285),
.B1(n_290),
.B2(n_295),
.C(n_297),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_240),
.C(n_272),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_214),
.B(n_239),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_197),
.B(n_213),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_178),
.B(n_196),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_155),
.B(n_177),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_133),
.B(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_137),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_138),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_145),
.C(n_150),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_164),
.B(n_176),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_163),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_160),
.A2(n_162),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_171),
.B(n_175),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_168),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_181),
.B(n_198),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_186),
.CI(n_189),
.CON(n_181),
.SN(n_181)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_193),
.Y(n_209)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_208),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_209),
.C(n_210),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_205),
.C(n_206),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_201),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_207),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_215),
.B(n_216),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_227),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_219),
.C(n_227),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_219)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_226),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_233),
.C(n_236),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_235),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_241),
.A2(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_259),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_242),
.B(n_259),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_254),
.C(n_258),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_246),
.C(n_253),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_253),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_250),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_258),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_257),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_259)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_268),
.C(n_271),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_265),
.C(n_266),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_283),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_283),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.C(n_282),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_286),
.A2(n_291),
.B(n_294),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);


endmodule