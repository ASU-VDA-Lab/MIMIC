module real_jpeg_31351_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_0),
.Y(n_136)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_1),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_1),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_1),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_1),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_1),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_1),
.B(n_321),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_2),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_3),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_3),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_3),
.B(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_3),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_3),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_4),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_4),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_4),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_4),
.B(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_6),
.Y(n_143)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_6),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_6),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_7),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_7),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_7),
.B(n_93),
.Y(n_92)
);

NAND2x1_ASAP7_75t_L g122 ( 
.A(n_7),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_7),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_8),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_8),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_8),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_8),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_8),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_8),
.B(n_244),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_8),
.B(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_9),
.Y(n_94)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_10),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_10),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_10),
.B(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_11),
.Y(n_129)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_12),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_13),
.Y(n_151)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_13),
.Y(n_211)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_14),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_14),
.B(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_14),
.B(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_14),
.B(n_87),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_15),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_15),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_15),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_15),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_15),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_15),
.B(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_193),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_192),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_169),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_20),
.B(n_169),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_103),
.Y(n_20)
);

MAJx2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.C(n_89),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_23),
.B(n_90),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_25),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.C(n_34),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_26),
.A2(n_27),
.B1(n_34),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_29),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_30),
.B(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_34),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_43),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_38),
.B(n_43),
.C(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_42),
.Y(n_161)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_47),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_49),
.B(n_171),
.Y(n_170)
);

OAI21x1_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_68),
.B(n_88),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_50),
.A2(n_51),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_52),
.Y(n_154)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_54),
.B(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_56),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_56),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_58),
.B(n_64),
.C(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_61),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_62),
.Y(n_238)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_65),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_65),
.B(n_316),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_67),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_77),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_77),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_69),
.A2(n_77),
.B1(n_78),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_69),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_70),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_70),
.B(n_108),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_114),
.Y(n_212)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_76),
.Y(n_322)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.C(n_85),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_79),
.A2(n_85),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_79),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_80),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_81),
.B(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_84),
.Y(n_205)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_84),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_85),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_96),
.C(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_130),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_108),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_108),
.A2(n_243),
.B1(n_247),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_120),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_155),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_144),
.C(n_152),
.Y(n_131)
);

XOR2x2_ASAP7_75t_L g190 ( 
.A(n_132),
.B(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_138),
.C(n_141),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_133),
.B(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_135),
.Y(n_279)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_146),
.B(n_148),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_153),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_159)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_190),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_170),
.B(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_190),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_185),
.C(n_186),
.Y(n_172)
);

XOR2x2_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_223),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.C(n_183),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_249)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_183),
.A2(n_184),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_187),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_226),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_224),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_224),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_217),
.C(n_222),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_212),
.C(n_213),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_212),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.C(n_206),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_L g287 ( 
.A(n_200),
.B(n_207),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_202),
.B(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_R g340 ( 
.A(n_202),
.B(n_287),
.Y(n_340)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_222),
.Y(n_252)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

OAI21x1_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_253),
.B(n_344),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_251),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_232),
.B(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.C(n_248),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_233),
.B(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_235),
.B(n_248),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.C(n_242),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_236),
.A2(n_239),
.B1(n_240),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_242),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_251),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_337),
.B(n_343),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_293),
.B(n_336),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_283),
.Y(n_255)
);

NAND2xp33_ASAP7_75t_L g336 ( 
.A(n_256),
.B(n_283),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_275),
.C(n_280),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_257),
.A2(n_258),
.B1(n_304),
.B2(n_306),
.Y(n_303)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_269),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_268),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_268),
.C(n_269),
.Y(n_285)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_280),
.B1(n_281),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_278),
.Y(n_296)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_290),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_289),
.B(n_339),
.C(n_340),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_290),
.Y(n_339)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_307),
.B(n_335),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_303),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_295),
.B(n_303),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.C(n_298),
.Y(n_295)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_332),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_297),
.Y(n_332)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_328),
.B(n_334),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_323),
.B(n_327),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_314),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_314),
.Y(n_327)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_315),
.B(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_320),
.Y(n_329)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_330),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_341),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_341),
.Y(n_343)
);


endmodule