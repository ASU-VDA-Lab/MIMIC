module fake_jpeg_18154_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_44),
.B(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_46),
.B(n_64),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_23),
.B1(n_25),
.B2(n_18),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_53),
.B1(n_67),
.B2(n_30),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_70),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_23),
.B1(n_25),
.B2(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_19),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_58),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_25),
.B1(n_27),
.B2(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_55),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_19),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_1),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_65),
.B(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_16),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_34),
.A2(n_24),
.B1(n_29),
.B2(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_72),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_33),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_1),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_73),
.B1(n_71),
.B2(n_63),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_40),
.B1(n_32),
.B2(n_30),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_89),
.B(n_58),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_46),
.A2(n_62),
.B1(n_26),
.B2(n_28),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_32),
.CI(n_29),
.CON(n_83),
.SN(n_83)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_83),
.B(n_94),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_60),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_86),
.C(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_101),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_28),
.C(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_95),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_51),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_SL g126 ( 
.A(n_96),
.B(n_5),
.C(n_7),
.Y(n_126)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_98),
.Y(n_111)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_14),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_3),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_3),
.C(n_4),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_123),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_110),
.B1(n_117),
.B2(n_130),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_73),
.B1(n_64),
.B2(n_59),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_68),
.B1(n_56),
.B2(n_59),
.Y(n_113)
);

AO22x1_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_80),
.B1(n_95),
.B2(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_124),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_68),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_121),
.B(n_10),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_48),
.B1(n_68),
.B2(n_52),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_52),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_48),
.B1(n_6),
.B2(n_7),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_98),
.B1(n_90),
.B2(n_13),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_14),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_126),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_7),
.C(n_9),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_102),
.C(n_101),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_78),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_10),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_147),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_104),
.B1(n_83),
.B2(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_139),
.Y(n_157)
);

AO21x2_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_91),
.B(n_94),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_143),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_89),
.B1(n_87),
.B2(n_86),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_144),
.A2(n_154),
.B(n_127),
.Y(n_160)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_11),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_11),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_149),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_122),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_152),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_111),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_150),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_109),
.B1(n_110),
.B2(n_105),
.Y(n_154)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_109),
.A3(n_123),
.B1(n_106),
.B2(n_118),
.C1(n_126),
.C2(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_148),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_107),
.B(n_113),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_160),
.B(n_163),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_118),
.C(n_113),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_164),
.C(n_165),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_124),
.B(n_127),
.C(n_144),
.D(n_154),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_137),
.C(n_132),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_133),
.C(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_135),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_161),
.C(n_139),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_136),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_180),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_143),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_140),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_181),
.B(n_140),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_140),
.B1(n_133),
.B2(n_134),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_184),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_186),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_157),
.B(n_162),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_187),
.A2(n_181),
.B(n_192),
.Y(n_200)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_194),
.B1(n_185),
.B2(n_140),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_155),
.B1(n_163),
.B2(n_140),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_155),
.B(n_164),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_184),
.B(n_173),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_176),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_200),
.A2(n_187),
.B(n_196),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

NAND4xp25_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_139),
.C(n_183),
.D(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_206),
.B1(n_196),
.B2(n_188),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_176),
.C(n_178),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_173),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_193),
.B(n_191),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_SL g207 ( 
.A(n_204),
.B(n_189),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_210),
.B(n_206),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_212),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_201),
.C(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_214),
.B(n_215),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_198),
.B(n_205),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_216),
.A2(n_210),
.B(n_198),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_217),
.A2(n_200),
.B(n_145),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_199),
.B(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_218),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_146),
.Y(n_223)
);


endmodule