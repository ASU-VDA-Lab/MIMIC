module fake_ibex_256_n_1150 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_195, n_163, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1150);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1150;

wire n_1084;
wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1011;
wire n_992;
wire n_1148;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_1143;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_418;
wire n_510;
wire n_845;
wire n_972;
wire n_947;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_1106;
wire n_1129;
wire n_449;
wire n_1131;
wire n_547;
wire n_1134;
wire n_727;
wire n_1138;
wire n_1077;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_1147;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_1140;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_1144;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_470;
wire n_276;
wire n_339;
wire n_259;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_1109;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_1112;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1068;
wire n_325;
wire n_301;
wire n_617;
wire n_496;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_1141;
wire n_694;
wire n_523;
wire n_787;
wire n_977;
wire n_1075;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_1081;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1101;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_1082;
wire n_1137;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_607;
wire n_427;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1028;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_1135;
wire n_973;
wire n_1146;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1142;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_433;
wire n_439;
wire n_299;
wire n_704;
wire n_949;
wire n_1007;
wire n_1126;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_1115;
wire n_935;
wire n_869;
wire n_998;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1100;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_567;
wire n_516;
wire n_548;
wire n_943;
wire n_1057;
wire n_1049;
wire n_763;
wire n_1086;
wire n_745;
wire n_329;
wire n_1149;
wire n_447;
wire n_940;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_706;
wire n_624;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_615;
wire n_512;
wire n_950;
wire n_685;
wire n_1026;
wire n_397;
wire n_366;
wire n_283;
wire n_894;
wire n_803;
wire n_1033;
wire n_1118;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_223;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_285;
wire n_379;
wire n_1128;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_1145;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_1139;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_1119;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_1095;
wire n_361;
wire n_1085;
wire n_455;
wire n_1136;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1005;
wire n_1102;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_874;
wire n_890;
wire n_816;
wire n_912;
wire n_921;
wire n_1105;
wire n_1058;
wire n_677;
wire n_489;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_1038;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_74),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_100),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_37),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_128),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_126),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_96),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_76),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_173),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_21),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_29),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_53),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_88),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_182),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_45),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_109),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_180),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_166),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_60),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_147),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_71),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_155),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_16),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_95),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_107),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_130),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_44),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_98),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_42),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_144),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_91),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_106),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_13),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_133),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_13),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_4),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_18),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_62),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_36),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_55),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_176),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_5),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_2),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_189),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_44),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_11),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_9),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_138),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_52),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_50),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_39),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_200),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_25),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_119),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_82),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_115),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_151),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_114),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_158),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_175),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_79),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_94),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_116),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_18),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_5),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_137),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_97),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_156),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_64),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_104),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_143),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_54),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_46),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_65),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_43),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_86),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_183),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_45),
.B(n_61),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_108),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_24),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_167),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_127),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_131),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_101),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_1),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_113),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_188),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_136),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_125),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_153),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_26),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_84),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_140),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_4),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_66),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_197),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_80),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_171),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_87),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_191),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_132),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_72),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_142),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_105),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_85),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_37),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_68),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_38),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_9),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_199),
.B(n_51),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_134),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_201),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_16),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_0),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_33),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_168),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_157),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_139),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_92),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_48),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_38),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_89),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_149),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_29),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_6),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_67),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_20),
.B(n_195),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_11),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_10),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_178),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_121),
.B(n_146),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_78),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_41),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_42),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_43),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_22),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_14),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_148),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_198),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_186),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_19),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_19),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_48),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_32),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_15),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_40),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_57),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_32),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_117),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_2),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_L g358 ( 
.A(n_0),
.B(n_124),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_10),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_202),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_276),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_343),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g363 ( 
.A(n_236),
.B(n_56),
.Y(n_363)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_236),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_354),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_280),
.B(n_3),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_202),
.Y(n_367)
);

OAI22x1_ASAP7_75t_R g368 ( 
.A1(n_336),
.A2(n_344),
.B1(n_342),
.B2(n_212),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g369 ( 
.A(n_236),
.B(n_58),
.Y(n_369)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_339),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_202),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_203),
.Y(n_372)
);

OAI22x1_ASAP7_75t_R g373 ( 
.A1(n_336),
.A2(n_344),
.B1(n_342),
.B2(n_212),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_252),
.Y(n_374)
);

OA21x2_ASAP7_75t_L g375 ( 
.A1(n_203),
.A2(n_103),
.B(n_196),
.Y(n_375)
);

CKINVDCx6p67_ASAP7_75t_R g376 ( 
.A(n_339),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_322),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_215),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_252),
.Y(n_379)
);

BUFx12f_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_202),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_247),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_210),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_269),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_215),
.Y(n_386)
);

INVx6_ASAP7_75t_L g387 ( 
.A(n_347),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_210),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_3),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_274),
.B(n_6),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_258),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_269),
.Y(n_392)
);

AOI22x1_ASAP7_75t_SL g393 ( 
.A1(n_224),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_306),
.B(n_12),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_220),
.A2(n_111),
.B(n_192),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_262),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_397)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_216),
.Y(n_398)
);

BUFx8_ASAP7_75t_SL g399 ( 
.A(n_224),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_258),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_17),
.Y(n_402)
);

OA21x2_ASAP7_75t_L g403 ( 
.A1(n_220),
.A2(n_118),
.B(n_190),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_269),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_226),
.B(n_244),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_343),
.B(n_20),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_214),
.B(n_23),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_240),
.B(n_24),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_225),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_244),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_206),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_225),
.B(n_27),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_219),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_304),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_219),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_209),
.B(n_28),
.Y(n_416)
);

OA21x2_ASAP7_75t_L g417 ( 
.A1(n_228),
.A2(n_123),
.B(n_187),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

BUFx12f_ASAP7_75t_L g419 ( 
.A(n_216),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_269),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_295),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_305),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_422)
);

BUFx12f_ASAP7_75t_L g423 ( 
.A(n_218),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_250),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_251),
.A2(n_135),
.B(n_185),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_251),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_271),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_286),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_288),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_288),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_242),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_296),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_245),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_204),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_272),
.B(n_34),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_326),
.B(n_35),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_282),
.B(n_35),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_227),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_292),
.B(n_36),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_271),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_286),
.Y(n_441)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_286),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_320),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_286),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_293),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_321),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_271),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_293),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_327),
.Y(n_449)
);

AOI22x1_ASAP7_75t_SL g450 ( 
.A1(n_257),
.A2(n_290),
.B1(n_323),
.B2(n_352),
.Y(n_450)
);

BUFx12f_ASAP7_75t_L g451 ( 
.A(n_218),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_340),
.Y(n_452)
);

BUFx8_ASAP7_75t_SL g453 ( 
.A(n_257),
.Y(n_453)
);

AND2x2_ASAP7_75t_SL g454 ( 
.A(n_317),
.B(n_141),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_348),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_205),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_349),
.B(n_40),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_312),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_271),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_350),
.B(n_47),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_312),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_353),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_314),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_359),
.B(n_49),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_231),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_207),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_234),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_217),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_238),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_229),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_232),
.B(n_49),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_466),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_398),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_360),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_363),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_378),
.B(n_296),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_385),
.B(n_221),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_461),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_461),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_370),
.B(n_394),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_360),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_411),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_364),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_385),
.B(n_221),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_364),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_398),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_364),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_387),
.B(n_233),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_360),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_370),
.B(n_345),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_377),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_364),
.Y(n_492)
);

BUFx4f_ASAP7_75t_L g493 ( 
.A(n_363),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_387),
.Y(n_494)
);

AND2x2_ASAP7_75t_SL g495 ( 
.A(n_454),
.B(n_235),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_466),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_367),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_432),
.B(n_346),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_367),
.Y(n_499)
);

AND2x2_ASAP7_75t_SL g500 ( 
.A(n_454),
.B(n_237),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_419),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_434),
.B(n_346),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_363),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_367),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_434),
.B(n_241),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_470),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_371),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_363),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_363),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_371),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_419),
.B(n_323),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_381),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_378),
.B(n_253),
.Y(n_513)
);

NOR2x1p5_ASAP7_75t_L g514 ( 
.A(n_376),
.B(n_254),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_381),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_377),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_456),
.B(n_260),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_423),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_456),
.B(n_287),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_362),
.B(n_208),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_384),
.Y(n_521)
);

BUFx4f_ASAP7_75t_L g522 ( 
.A(n_369),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_387),
.B(n_298),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_384),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_386),
.B(n_301),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_386),
.B(n_313),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_470),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_362),
.B(n_211),
.Y(n_528)
);

OAI22xp33_ASAP7_75t_L g529 ( 
.A1(n_366),
.A2(n_316),
.B1(n_315),
.B2(n_328),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_401),
.B(n_331),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_369),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_372),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_455),
.B(n_332),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_372),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_392),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_380),
.B(n_285),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_455),
.B(n_335),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_404),
.Y(n_538)
);

CKINVDCx8_ASAP7_75t_R g539 ( 
.A(n_368),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_438),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_436),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_382),
.B(n_255),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_361),
.B(n_256),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_436),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_404),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_383),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_365),
.B(n_213),
.Y(n_547)
);

AO21x2_ASAP7_75t_L g548 ( 
.A1(n_412),
.A2(n_396),
.B(n_407),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_438),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_L g550 ( 
.A1(n_397),
.A2(n_355),
.B1(n_249),
.B2(n_341),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_423),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_420),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_383),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_380),
.B(n_222),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_451),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_467),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_374),
.B(n_261),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_388),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_388),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_379),
.B(n_465),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_413),
.B(n_351),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_428),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_428),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_428),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_436),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_409),
.Y(n_566)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_467),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_399),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_441),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_441),
.Y(n_570)
);

INVx8_ASAP7_75t_L g571 ( 
.A(n_369),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_441),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_441),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_444),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_413),
.B(n_223),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_444),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_444),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_426),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_444),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_447),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_426),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_414),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_468),
.B(n_230),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_465),
.B(n_239),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_429),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_447),
.Y(n_586)
);

AOI21x1_ASAP7_75t_L g587 ( 
.A1(n_412),
.A2(n_311),
.B(n_268),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_429),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_430),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_430),
.Y(n_590)
);

BUFx6f_ASAP7_75t_SL g591 ( 
.A(n_369),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_447),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_469),
.B(n_263),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_448),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_447),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_459),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_459),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_459),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_448),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_459),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_442),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_442),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_442),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_442),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_458),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_431),
.B(n_270),
.Y(n_606)
);

AOI21x1_ASAP7_75t_L g607 ( 
.A1(n_390),
.A2(n_324),
.B(n_356),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_414),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_476),
.B(n_389),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_482),
.B(n_451),
.Y(n_610)
);

AOI22x1_ASAP7_75t_SL g611 ( 
.A1(n_473),
.A2(n_399),
.B1(n_453),
.B2(n_405),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_571),
.B(n_369),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_476),
.B(n_406),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_575),
.B(n_471),
.Y(n_614)
);

OAI221xp5_ASAP7_75t_L g615 ( 
.A1(n_549),
.A2(n_435),
.B1(n_408),
.B2(n_457),
.C(n_460),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_575),
.B(n_418),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_533),
.B(n_418),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_508),
.B(n_437),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_L g619 ( 
.A(n_501),
.B(n_445),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_495),
.A2(n_464),
.B1(n_437),
.B2(n_439),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_495),
.A2(n_402),
.B1(n_464),
.B2(n_439),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g622 ( 
.A(n_550),
.B(n_410),
.C(n_421),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_483),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_533),
.B(n_416),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_483),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_485),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_556),
.B(n_402),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_537),
.B(n_477),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_537),
.B(n_416),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_485),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_532),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_561),
.B(n_433),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_532),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_561),
.B(n_443),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_484),
.B(n_446),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_518),
.B(n_422),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_490),
.B(n_449),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_505),
.B(n_452),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_534),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_546),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_500),
.A2(n_462),
.B1(n_395),
.B2(n_391),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_513),
.B(n_400),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_540),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_546),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_571),
.B(n_243),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_473),
.Y(n_646)
);

NOR2x1p5_ASAP7_75t_L g647 ( 
.A(n_501),
.B(n_373),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_486),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_513),
.B(n_415),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_L g650 ( 
.A(n_529),
.B(n_424),
.C(n_277),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_553),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_493),
.B(n_246),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_517),
.B(n_519),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_553),
.Y(n_654)
);

AND2x2_ASAP7_75t_SL g655 ( 
.A(n_500),
.B(n_375),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_525),
.B(n_248),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_502),
.B(n_424),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_487),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_526),
.B(n_259),
.Y(n_659)
);

BUFx5_ASAP7_75t_L g660 ( 
.A(n_503),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_526),
.B(n_583),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_571),
.B(n_264),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_584),
.B(n_265),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_522),
.B(n_266),
.Y(n_664)
);

INVxp33_ASAP7_75t_SL g665 ( 
.A(n_486),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_584),
.B(n_560),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_530),
.B(n_458),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_593),
.B(n_267),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_522),
.B(n_273),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_558),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_488),
.B(n_275),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_559),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_492),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_475),
.B(n_278),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_608),
.B(n_279),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_567),
.B(n_281),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_518),
.B(n_453),
.Y(n_677)
);

BUFx6f_ASAP7_75t_SL g678 ( 
.A(n_536),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_531),
.B(n_283),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_539),
.A2(n_393),
.B1(n_445),
.B2(n_463),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_523),
.B(n_284),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_531),
.B(n_294),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_514),
.B(n_450),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_543),
.B(n_299),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_480),
.B(n_289),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_566),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_491),
.B(n_445),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_542),
.B(n_300),
.Y(n_688)
);

OR2x6_ASAP7_75t_L g689 ( 
.A(n_514),
.B(n_334),
.Y(n_689)
);

NOR2xp67_ASAP7_75t_L g690 ( 
.A(n_551),
.B(n_445),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_520),
.B(n_291),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_539),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_L g693 ( 
.A1(n_511),
.A2(n_463),
.B1(n_358),
.B2(n_325),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_544),
.A2(n_463),
.B1(n_375),
.B2(n_403),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_544),
.B(n_302),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_472),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_528),
.B(n_307),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_491),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_565),
.B(n_303),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_565),
.B(n_308),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_606),
.B(n_309),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_L g702 ( 
.A(n_551),
.B(n_463),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_547),
.B(n_310),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_503),
.B(n_318),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_472),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_516),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_582),
.B(n_319),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_494),
.B(n_329),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_494),
.B(n_330),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_472),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_557),
.B(n_333),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_555),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_655),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_643),
.B(n_509),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_R g715 ( 
.A(n_712),
.B(n_555),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_643),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_623),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_706),
.B(n_498),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_706),
.B(n_554),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_655),
.A2(n_548),
.B(n_509),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_628),
.B(n_541),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_694),
.A2(n_548),
.B(n_403),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_694),
.A2(n_607),
.B(n_587),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_638),
.A2(n_578),
.B(n_605),
.C(n_581),
.Y(n_724)
);

NAND2x1p5_ASAP7_75t_L g725 ( 
.A(n_698),
.B(n_578),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_631),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_L g727 ( 
.A(n_653),
.B(n_568),
.C(n_536),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_621),
.A2(n_591),
.B1(n_607),
.B2(n_599),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_632),
.B(n_581),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_634),
.B(n_585),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_618),
.A2(n_425),
.B(n_417),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_620),
.A2(n_661),
.B1(n_641),
.B2(n_615),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_638),
.B(n_585),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_637),
.A2(n_635),
.B(n_666),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_609),
.B(n_588),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_613),
.B(n_588),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_617),
.A2(n_590),
.B(n_589),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_614),
.A2(n_591),
.B1(n_590),
.B2(n_589),
.Y(n_738)
);

BUFx4f_ASAP7_75t_L g739 ( 
.A(n_683),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_667),
.B(n_594),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_624),
.B(n_594),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_629),
.A2(n_605),
.B(n_599),
.C(n_337),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_616),
.B(n_536),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_649),
.B(n_536),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_627),
.B(n_604),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_642),
.B(n_663),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_650),
.A2(n_496),
.B1(n_506),
.B2(n_527),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_657),
.A2(n_506),
.B(n_527),
.C(n_440),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_610),
.B(n_601),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_633),
.A2(n_506),
.B(n_527),
.C(n_440),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_656),
.B(n_427),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_646),
.B(n_427),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_648),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_639),
.A2(n_644),
.B(n_640),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_650),
.B(n_604),
.C(n_603),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_659),
.B(n_602),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_677),
.B(n_603),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_703),
.B(n_478),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_651),
.A2(n_479),
.B1(n_478),
.B2(n_338),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_703),
.B(n_59),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_654),
.A2(n_600),
.B(n_598),
.C(n_597),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_695),
.A2(n_538),
.B(n_489),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_670),
.A2(n_600),
.B(n_598),
.C(n_597),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_625),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_687),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_622),
.A2(n_596),
.B(n_595),
.C(n_592),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_676),
.B(n_691),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_626),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_699),
.A2(n_545),
.B(n_497),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_630),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_672),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_636),
.B(n_63),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_691),
.B(n_697),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_697),
.B(n_69),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_636),
.B(n_70),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_700),
.A2(n_552),
.B(n_507),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_SL g777 ( 
.A1(n_678),
.A2(n_596),
.B1(n_595),
.B2(n_592),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_658),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_686),
.A2(n_535),
.B(n_499),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_685),
.B(n_73),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_622),
.A2(n_586),
.B1(n_580),
.B2(n_579),
.Y(n_781)
);

OAI21xp33_ASAP7_75t_L g782 ( 
.A1(n_684),
.A2(n_586),
.B(n_580),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_685),
.B(n_75),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_636),
.A2(n_577),
.B1(n_576),
.B2(n_574),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_673),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_708),
.A2(n_573),
.B1(n_572),
.B2(n_570),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_701),
.B(n_77),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_688),
.B(n_83),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_660),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_689),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_696),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_709),
.A2(n_524),
.B(n_564),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_647),
.B(n_90),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_668),
.A2(n_524),
.B1(n_564),
.B2(n_563),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_674),
.A2(n_682),
.B(n_679),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_705),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_709),
.A2(n_521),
.B(n_563),
.C(n_562),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_689),
.B(n_93),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_711),
.B(n_99),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_716),
.B(n_683),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_734),
.B(n_681),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_753),
.B(n_683),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_729),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_725),
.Y(n_804)
);

AO21x2_ASAP7_75t_L g805 ( 
.A1(n_722),
.A2(n_693),
.B(n_652),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_731),
.A2(n_662),
.B(n_645),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_734),
.B(n_680),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_732),
.B(n_680),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_746),
.B(n_619),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_720),
.A2(n_664),
.B(n_669),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_730),
.B(n_690),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_725),
.B(n_689),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_720),
.A2(n_704),
.B(n_675),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_723),
.A2(n_671),
.B(n_707),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_718),
.B(n_702),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_772),
.B(n_692),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_721),
.B(n_693),
.Y(n_817)
);

AOI21xp33_ASAP7_75t_L g818 ( 
.A1(n_766),
.A2(n_710),
.B(n_521),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_757),
.B(n_611),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_726),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_740),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_715),
.Y(n_822)
);

BUFx4_ASAP7_75t_SL g823 ( 
.A(n_727),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_771),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_767),
.A2(n_515),
.B(n_504),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_735),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_775),
.B(n_660),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_744),
.B(n_102),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_717),
.Y(n_829)
);

NAND2x1p5_ASAP7_75t_L g830 ( 
.A(n_764),
.B(n_569),
.Y(n_830)
);

OAI21x1_ASAP7_75t_SL g831 ( 
.A1(n_754),
.A2(n_110),
.B(n_112),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_773),
.B(n_120),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_736),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_724),
.A2(n_512),
.B(n_510),
.Y(n_834)
);

BUFx12f_ASAP7_75t_L g835 ( 
.A(n_790),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_SL g836 ( 
.A1(n_798),
.A2(n_719),
.B(n_745),
.C(n_749),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_733),
.B(n_122),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_751),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_764),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_743),
.B(n_145),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_739),
.Y(n_841)
);

AO31x2_ASAP7_75t_L g842 ( 
.A1(n_742),
.A2(n_481),
.A3(n_474),
.B(n_154),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_741),
.B(n_150),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_752),
.B(n_152),
.Y(n_844)
);

AO31x2_ASAP7_75t_L g845 ( 
.A1(n_738),
.A2(n_797),
.A3(n_728),
.B(n_748),
.Y(n_845)
);

AO22x1_ASAP7_75t_L g846 ( 
.A1(n_793),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_737),
.A2(n_713),
.B1(n_755),
.B2(n_760),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_765),
.B(n_163),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_756),
.B(n_164),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_781),
.A2(n_165),
.B(n_169),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_778),
.B(n_170),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_761),
.A2(n_172),
.B(n_174),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_763),
.A2(n_177),
.B(n_179),
.Y(n_853)
);

NAND2x1p5_ASAP7_75t_L g854 ( 
.A(n_778),
.B(n_789),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_768),
.B(n_770),
.Y(n_855)
);

BUFx12f_ASAP7_75t_L g856 ( 
.A(n_739),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_785),
.B(n_713),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_713),
.B(n_747),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_758),
.Y(n_859)
);

AOI21xp33_ASAP7_75t_L g860 ( 
.A1(n_784),
.A2(n_774),
.B(n_780),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_779),
.A2(n_769),
.B(n_776),
.Y(n_861)
);

AOI21x1_ASAP7_75t_L g862 ( 
.A1(n_787),
.A2(n_788),
.B(n_799),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_714),
.B(n_796),
.Y(n_863)
);

AO31x2_ASAP7_75t_L g864 ( 
.A1(n_759),
.A2(n_750),
.A3(n_794),
.B(n_783),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_791),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_777),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_786),
.B(n_792),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_795),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_782),
.A2(n_762),
.B(n_795),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_716),
.B(n_706),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_720),
.A2(n_722),
.B(n_723),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_726),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_720),
.A2(n_722),
.B(n_723),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_716),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_734),
.B(n_732),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_734),
.B(n_732),
.Y(n_876)
);

INVx4_ASAP7_75t_SL g877 ( 
.A(n_726),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_753),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_725),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_729),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_729),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_720),
.A2(n_722),
.B(n_723),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_720),
.A2(n_722),
.B(n_723),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_716),
.B(n_405),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_716),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_726),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_722),
.A2(n_612),
.B(n_522),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_720),
.A2(n_722),
.B(n_723),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_734),
.A2(n_495),
.B1(n_500),
.B2(n_733),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_722),
.A2(n_612),
.B(n_522),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_734),
.B(n_732),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_734),
.B(n_732),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_726),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_720),
.A2(n_722),
.B(n_723),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_716),
.B(n_746),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_725),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_889),
.A2(n_821),
.B1(n_808),
.B2(n_875),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_896),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_826),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_895),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_824),
.Y(n_901)
);

AOI21xp33_ASAP7_75t_L g902 ( 
.A1(n_836),
.A2(n_891),
.B(n_876),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_895),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_829),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_878),
.Y(n_905)
);

AO21x2_ASAP7_75t_L g906 ( 
.A1(n_871),
.A2(n_894),
.B(n_883),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_803),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_889),
.A2(n_807),
.B1(n_817),
.B2(n_833),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_856),
.Y(n_909)
);

OA21x2_ASAP7_75t_L g910 ( 
.A1(n_871),
.A2(n_894),
.B(n_873),
.Y(n_910)
);

INVx4_ASAP7_75t_L g911 ( 
.A(n_877),
.Y(n_911)
);

AOI221xp5_ASAP7_75t_L g912 ( 
.A1(n_880),
.A2(n_881),
.B1(n_892),
.B2(n_821),
.C(n_859),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_855),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_886),
.Y(n_914)
);

CKINVDCx16_ASAP7_75t_R g915 ( 
.A(n_835),
.Y(n_915)
);

AOI21xp33_ASAP7_75t_L g916 ( 
.A1(n_847),
.A2(n_801),
.B(n_814),
.Y(n_916)
);

NOR2x1_ASAP7_75t_L g917 ( 
.A(n_870),
.B(n_879),
.Y(n_917)
);

OAI21x1_ASAP7_75t_SL g918 ( 
.A1(n_850),
.A2(n_831),
.B(n_853),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_804),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_838),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_879),
.B(n_841),
.Y(n_921)
);

OR2x6_ASAP7_75t_L g922 ( 
.A(n_827),
.B(n_874),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_885),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_822),
.Y(n_924)
);

AO31x2_ASAP7_75t_L g925 ( 
.A1(n_847),
.A2(n_869),
.A3(n_890),
.B(n_887),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_809),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_815),
.B(n_828),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_811),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_884),
.B(n_812),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_857),
.B(n_858),
.Y(n_930)
);

OAI221xp5_ASAP7_75t_L g931 ( 
.A1(n_802),
.A2(n_888),
.B1(n_883),
.B2(n_882),
.C(n_873),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_827),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_877),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_844),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_893),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_877),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_893),
.Y(n_937)
);

NAND3xp33_ASAP7_75t_L g938 ( 
.A(n_868),
.B(n_813),
.C(n_846),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_848),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_L g940 ( 
.A(n_868),
.B(n_810),
.C(n_852),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_863),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_865),
.B(n_839),
.Y(n_942)
);

NAND3xp33_ASAP7_75t_SL g943 ( 
.A(n_850),
.B(n_814),
.C(n_853),
.Y(n_943)
);

BUFx12f_ASAP7_75t_L g944 ( 
.A(n_816),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_865),
.B(n_839),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_819),
.A2(n_816),
.B1(n_858),
.B2(n_867),
.Y(n_946)
);

AO21x2_ASAP7_75t_L g947 ( 
.A1(n_861),
.A2(n_860),
.B(n_862),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_823),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_800),
.B(n_854),
.Y(n_949)
);

OAI21x1_ASAP7_75t_SL g950 ( 
.A1(n_852),
.A2(n_810),
.B(n_806),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_832),
.A2(n_837),
.B(n_843),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_854),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_866),
.A2(n_840),
.B1(n_805),
.B2(n_849),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_851),
.Y(n_954)
);

AO21x2_ASAP7_75t_L g955 ( 
.A1(n_805),
.A2(n_818),
.B(n_834),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_820),
.B(n_872),
.Y(n_956)
);

BUFx8_ASAP7_75t_L g957 ( 
.A(n_866),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_845),
.B(n_830),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_845),
.B(n_830),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_845),
.B(n_864),
.Y(n_960)
);

AOI22x1_ASAP7_75t_L g961 ( 
.A1(n_825),
.A2(n_834),
.B1(n_864),
.B2(n_842),
.Y(n_961)
);

BUFx2_ASAP7_75t_R g962 ( 
.A(n_842),
.Y(n_962)
);

AO31x2_ASAP7_75t_L g963 ( 
.A1(n_864),
.A2(n_847),
.A3(n_876),
.B(n_875),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_875),
.A2(n_892),
.B(n_891),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_895),
.A2(n_405),
.B1(n_665),
.B2(n_706),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_826),
.Y(n_966)
);

AO21x2_ASAP7_75t_L g967 ( 
.A1(n_871),
.A2(n_882),
.B(n_873),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_822),
.Y(n_968)
);

BUFx4f_ASAP7_75t_L g969 ( 
.A(n_856),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_833),
.B(n_734),
.Y(n_970)
);

NAND3xp33_ASAP7_75t_L g971 ( 
.A(n_868),
.B(n_727),
.C(n_650),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_826),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_850),
.A2(n_892),
.B(n_876),
.Y(n_973)
);

NAND2x1p5_ASAP7_75t_L g974 ( 
.A(n_879),
.B(n_821),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_826),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_911),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_898),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_970),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_930),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_911),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_899),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_931),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_915),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_910),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_931),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_912),
.A2(n_908),
.B1(n_899),
.B2(n_897),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_922),
.Y(n_987)
);

INVx4_ASAP7_75t_L g988 ( 
.A(n_922),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_941),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_913),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_974),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_923),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_964),
.A2(n_908),
.B(n_897),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_912),
.A2(n_946),
.B1(n_934),
.B2(n_932),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_901),
.Y(n_995)
);

OAI222xp33_ASAP7_75t_L g996 ( 
.A1(n_922),
.A2(n_946),
.B1(n_965),
.B2(n_905),
.C1(n_917),
.C2(n_932),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_907),
.Y(n_997)
);

AO21x2_ASAP7_75t_L g998 ( 
.A1(n_943),
.A2(n_950),
.B(n_902),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_958),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_920),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_929),
.A2(n_944),
.B1(n_926),
.B2(n_928),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_904),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_919),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_960),
.B(n_906),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_SL g1005 ( 
.A1(n_957),
.A2(n_918),
.B1(n_921),
.B2(n_972),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_963),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_906),
.B(n_967),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_963),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_967),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_914),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_959),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_921),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_964),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_929),
.A2(n_927),
.B1(n_971),
.B2(n_903),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_956),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_966),
.B(n_975),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_914),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_978),
.Y(n_1018)
);

INVx6_ASAP7_75t_L g1019 ( 
.A(n_980),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_978),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1004),
.B(n_947),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_981),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_977),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_983),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_1011),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1004),
.B(n_982),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_985),
.A2(n_948),
.B1(n_927),
.B2(n_957),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_L g1028 ( 
.A(n_1001),
.B(n_902),
.C(n_961),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_1014),
.A2(n_962),
.B(n_953),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_980),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_990),
.B(n_900),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_992),
.B(n_909),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_1003),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_999),
.B(n_955),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1006),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_990),
.B(n_949),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_977),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_977),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1006),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_995),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_976),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_976),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_1007),
.B(n_925),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_994),
.A2(n_939),
.B1(n_954),
.B2(n_943),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_999),
.B(n_955),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1007),
.B(n_925),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1025),
.B(n_1011),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1026),
.B(n_1008),
.Y(n_1048)
);

OR2x6_ASAP7_75t_SL g1049 ( 
.A(n_1034),
.B(n_986),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_1022),
.Y(n_1050)
);

AND2x4_ASAP7_75t_SL g1051 ( 
.A(n_1030),
.B(n_987),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_1019),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1026),
.B(n_1008),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1035),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1035),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1046),
.B(n_1009),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1046),
.B(n_1009),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1039),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_1025),
.B(n_986),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_1021),
.B(n_993),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1021),
.B(n_993),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1043),
.B(n_984),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_1023),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1018),
.B(n_979),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1018),
.B(n_979),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1054),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1061),
.B(n_1043),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1061),
.B(n_1043),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1050),
.B(n_1040),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1054),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1056),
.B(n_1043),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1050),
.B(n_1033),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1056),
.B(n_1045),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_1063),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_1052),
.B(n_1024),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1057),
.B(n_1045),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_1060),
.B(n_1034),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_1063),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1048),
.B(n_1020),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1055),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_1079),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1074),
.B(n_1060),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1069),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1066),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1066),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_1079),
.B(n_1052),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_1078),
.B(n_1057),
.Y(n_1088)
);

OR2x2_ASAP7_75t_L g1089 ( 
.A(n_1078),
.B(n_1047),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1070),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1070),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1081),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1073),
.B(n_1077),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1081),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1072),
.Y(n_1095)
);

INVxp67_ASAP7_75t_SL g1096 ( 
.A(n_1087),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1089),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_SL g1098 ( 
.A1(n_1087),
.A2(n_1075),
.B(n_1076),
.C(n_996),
.Y(n_1098)
);

AOI32xp33_ASAP7_75t_L g1099 ( 
.A1(n_1082),
.A2(n_1075),
.A3(n_1071),
.B1(n_1067),
.B2(n_1068),
.Y(n_1099)
);

NAND5xp2_ASAP7_75t_L g1100 ( 
.A(n_1095),
.B(n_1005),
.C(n_1027),
.D(n_1044),
.E(n_1029),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_1088),
.B(n_1073),
.Y(n_1101)
);

INVxp67_ASAP7_75t_SL g1102 ( 
.A(n_1091),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1093),
.A2(n_1049),
.B1(n_1019),
.B2(n_1030),
.Y(n_1103)
);

NAND4xp75_ASAP7_75t_L g1104 ( 
.A(n_1084),
.B(n_1068),
.C(n_1067),
.D(n_1071),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1085),
.B(n_1077),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1093),
.A2(n_1049),
.B1(n_1047),
.B2(n_1059),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1083),
.B(n_1080),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1091),
.Y(n_1108)
);

AOI321xp33_ASAP7_75t_L g1109 ( 
.A1(n_1106),
.A2(n_994),
.A3(n_1059),
.B1(n_1053),
.B2(n_1090),
.C(n_1086),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1104),
.A2(n_1019),
.B1(n_1030),
.B2(n_1051),
.Y(n_1110)
);

AOI321xp33_ASAP7_75t_L g1111 ( 
.A1(n_1106),
.A2(n_1103),
.A3(n_1096),
.B1(n_1097),
.B2(n_1105),
.C(n_1100),
.Y(n_1111)
);

OAI322xp33_ASAP7_75t_L g1112 ( 
.A1(n_1101),
.A2(n_1092),
.A3(n_1094),
.B1(n_1032),
.B2(n_1065),
.C1(n_1064),
.C2(n_1058),
.Y(n_1112)
);

OAI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1102),
.A2(n_1019),
.B1(n_1037),
.B2(n_1038),
.Y(n_1113)
);

AOI21xp33_ASAP7_75t_SL g1114 ( 
.A1(n_1099),
.A2(n_1042),
.B(n_1041),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1105),
.A2(n_1051),
.B(n_969),
.C(n_976),
.Y(n_1115)
);

NAND4xp25_ASAP7_75t_SL g1116 ( 
.A(n_1107),
.B(n_968),
.C(n_1028),
.D(n_1012),
.Y(n_1116)
);

AOI22x1_ASAP7_75t_L g1117 ( 
.A1(n_1111),
.A2(n_1098),
.B1(n_980),
.B2(n_988),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1114),
.B(n_1108),
.Y(n_1118)
);

NOR5xp2_ASAP7_75t_L g1119 ( 
.A(n_1112),
.B(n_938),
.C(n_940),
.D(n_916),
.E(n_1013),
.Y(n_1119)
);

OAI22x1_ASAP7_75t_L g1120 ( 
.A1(n_1116),
.A2(n_987),
.B1(n_988),
.B2(n_1042),
.Y(n_1120)
);

OAI21xp33_ASAP7_75t_L g1121 ( 
.A1(n_1115),
.A2(n_1094),
.B(n_1062),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1113),
.B(n_1055),
.Y(n_1122)
);

NOR4xp25_ASAP7_75t_L g1123 ( 
.A(n_1109),
.B(n_1016),
.C(n_997),
.D(n_1000),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_L g1124 ( 
.A(n_1118),
.B(n_1122),
.C(n_1121),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1117),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1123),
.B(n_1110),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1120),
.B(n_1058),
.Y(n_1127)
);

NAND2x1_ASAP7_75t_SL g1128 ( 
.A(n_1119),
.B(n_980),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1127),
.Y(n_1129)
);

NOR4xp25_ASAP7_75t_L g1130 ( 
.A(n_1125),
.B(n_997),
.C(n_1000),
.D(n_995),
.Y(n_1130)
);

NAND3xp33_ASAP7_75t_SL g1131 ( 
.A(n_1126),
.B(n_968),
.C(n_924),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_SL g1132 ( 
.A1(n_1128),
.A2(n_987),
.B(n_988),
.Y(n_1132)
);

AO22x2_ASAP7_75t_L g1133 ( 
.A1(n_1124),
.A2(n_987),
.B1(n_988),
.B2(n_989),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1131),
.B(n_969),
.Y(n_1134)
);

NOR4xp75_ASAP7_75t_L g1135 ( 
.A(n_1132),
.B(n_976),
.C(n_973),
.D(n_1041),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1129),
.B(n_1130),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1134),
.A2(n_1133),
.B(n_989),
.Y(n_1137)
);

OAI322xp33_ASAP7_75t_L g1138 ( 
.A1(n_1136),
.A2(n_1133),
.A3(n_1012),
.B1(n_1031),
.B2(n_1015),
.C1(n_1036),
.C2(n_991),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1135),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1138),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1137),
.B(n_1139),
.Y(n_1141)
);

XOR2x1_ASAP7_75t_L g1142 ( 
.A(n_1139),
.B(n_933),
.Y(n_1142)
);

OA22x2_ASAP7_75t_L g1143 ( 
.A1(n_1140),
.A2(n_1141),
.B1(n_1142),
.B2(n_1051),
.Y(n_1143)
);

OA22x2_ASAP7_75t_L g1144 ( 
.A1(n_1143),
.A2(n_936),
.B1(n_933),
.B2(n_1010),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1144),
.A2(n_951),
.B(n_942),
.Y(n_1145)
);

AOI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1145),
.A2(n_945),
.B1(n_942),
.B2(n_952),
.C(n_937),
.Y(n_1146)
);

OAI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1146),
.A2(n_1017),
.B1(n_1010),
.B2(n_952),
.Y(n_1147)
);

OA21x2_ASAP7_75t_L g1148 ( 
.A1(n_1147),
.A2(n_945),
.B(n_951),
.Y(n_1148)
);

AOI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_1148),
.A2(n_937),
.B1(n_935),
.B2(n_1010),
.C(n_1002),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1149),
.A2(n_1010),
.B1(n_1017),
.B2(n_998),
.Y(n_1150)
);


endmodule