module real_aes_8355_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_519;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g163 ( .A(n_0), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_0), .A2(n_498), .B1(n_511), .B2(n_519), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_1), .A2(n_49), .B1(n_482), .B2(n_484), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_2), .A2(n_30), .B1(n_90), .B2(n_99), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_3), .B(n_110), .Y(n_174) );
AND2x6_ASAP7_75t_L g108 ( .A(n_4), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g494 ( .A(n_4), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_4), .B(n_524), .Y(n_523) );
AO22x2_ASAP7_75t_L g401 ( .A1(n_5), .A2(n_25), .B1(n_402), .B2(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g106 ( .A(n_6), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_7), .B(n_97), .Y(n_117) );
INVx1_ASAP7_75t_L g155 ( .A(n_8), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_9), .B(n_111), .Y(n_179) );
AO32x2_ASAP7_75t_L g142 ( .A1(n_10), .A2(n_107), .A3(n_110), .B1(n_143), .B2(n_147), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g121 ( .A(n_11), .B(n_99), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_12), .B(n_111), .Y(n_165) );
AO22x2_ASAP7_75t_L g405 ( .A1(n_13), .A2(n_28), .B1(n_402), .B2(n_406), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_14), .A2(n_40), .B1(n_90), .B2(n_99), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_15), .A2(n_42), .B1(n_506), .B2(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_15), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g96 ( .A1(n_16), .A2(n_62), .B1(n_97), .B2(n_99), .Y(n_96) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_17), .B(n_99), .Y(n_136) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_18), .A2(n_32), .B1(n_464), .B2(n_469), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_19), .A2(n_58), .B1(n_474), .B2(n_478), .Y(n_473) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_20), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_21), .B(n_102), .Y(n_199) );
AOI22xp5_ASAP7_75t_SL g390 ( .A1(n_22), .A2(n_391), .B1(n_392), .B2(n_487), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_22), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_23), .B(n_102), .Y(n_140) );
INVx2_ASAP7_75t_L g92 ( .A(n_24), .Y(n_92) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_26), .B(n_99), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_27), .B(n_102), .Y(n_124) );
OAI221xp5_ASAP7_75t_L g514 ( .A1(n_28), .A2(n_45), .B1(n_56), .B2(n_515), .C(n_516), .Y(n_514) );
INVxp67_ASAP7_75t_L g517 ( .A(n_28), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g453 ( .A1(n_29), .A2(n_57), .B1(n_454), .B2(n_459), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_31), .Y(n_424) );
OAI22xp5_ASAP7_75t_SL g500 ( .A1(n_33), .A2(n_41), .B1(n_501), .B2(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_33), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_34), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_35), .B(n_99), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g89 ( .A1(n_36), .A2(n_69), .B1(n_90), .B2(n_93), .Y(n_89) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_37), .B(n_99), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_38), .B(n_99), .Y(n_157) );
INVx1_ASAP7_75t_L g529 ( .A(n_38), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_39), .B(n_161), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_41), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g183 ( .A1(n_42), .A2(n_47), .B1(n_97), .B2(n_99), .Y(n_183) );
INVx1_ASAP7_75t_L g506 ( .A(n_42), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_43), .B(n_99), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_44), .B(n_99), .Y(n_198) );
AO22x2_ASAP7_75t_L g411 ( .A1(n_45), .A2(n_65), .B1(n_402), .B2(n_406), .Y(n_411) );
INVxp67_ASAP7_75t_L g518 ( .A(n_45), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_46), .Y(n_412) );
INVx1_ASAP7_75t_L g109 ( .A(n_48), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_50), .B(n_99), .Y(n_164) );
INVx1_ASAP7_75t_L g105 ( .A(n_51), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_52), .Y(n_515) );
AO32x2_ASAP7_75t_L g87 ( .A1(n_53), .A2(n_88), .A3(n_101), .B1(n_107), .B2(n_110), .Y(n_87) );
INVx1_ASAP7_75t_L g197 ( .A(n_54), .Y(n_197) );
INVx1_ASAP7_75t_L g132 ( .A(n_55), .Y(n_132) );
AO22x2_ASAP7_75t_L g409 ( .A1(n_56), .A2(n_71), .B1(n_402), .B2(n_403), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_59), .B(n_97), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_60), .A2(n_504), .B1(n_505), .B2(n_508), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_60), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_61), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_63), .B(n_90), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_64), .B(n_97), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_66), .Y(n_395) );
INVx2_ASAP7_75t_L g103 ( .A(n_67), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_68), .B(n_97), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_70), .A2(n_76), .B1(n_97), .B2(n_98), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_72), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_73), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g402 ( .A(n_74), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_74), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_75), .B(n_97), .Y(n_195) );
AOI221xp5_ASAP7_75t_SL g77 ( .A1(n_78), .A2(n_384), .B1(n_389), .B2(n_488), .C(n_495), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
AND3x1_ASAP7_75t_L g81 ( .A(n_82), .B(n_304), .C(n_352), .Y(n_81) );
NOR4xp25_ASAP7_75t_L g82 ( .A(n_83), .B(n_232), .C(n_277), .D(n_291), .Y(n_82) );
OAI311xp33_ASAP7_75t_L g83 ( .A1(n_84), .A2(n_148), .A3(n_175), .B1(n_185), .C1(n_200), .Y(n_83) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_85), .B(n_112), .Y(n_84) );
OAI21xp33_ASAP7_75t_L g185 ( .A1(n_85), .A2(n_186), .B(n_188), .Y(n_185) );
AND2x2_ASAP7_75t_L g293 ( .A(n_85), .B(n_220), .Y(n_293) );
AND2x2_ASAP7_75t_L g350 ( .A(n_85), .B(n_236), .Y(n_350) );
BUFx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g243 ( .A(n_86), .B(n_141), .Y(n_243) );
AND2x2_ASAP7_75t_L g300 ( .A(n_86), .B(n_248), .Y(n_300) );
INVx1_ASAP7_75t_L g341 ( .A(n_86), .Y(n_341) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_87), .Y(n_209) );
AND2x2_ASAP7_75t_L g250 ( .A(n_87), .B(n_141), .Y(n_250) );
AND2x2_ASAP7_75t_L g254 ( .A(n_87), .B(n_142), .Y(n_254) );
INVx1_ASAP7_75t_L g266 ( .A(n_87), .Y(n_266) );
OAI22xp5_ASAP7_75t_SL g88 ( .A1(n_89), .A2(n_94), .B1(n_96), .B2(n_100), .Y(n_88) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
BUFx3_ASAP7_75t_L g93 ( .A(n_91), .Y(n_93) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_91), .Y(n_99) );
AND2x6_ASAP7_75t_L g387 ( .A(n_91), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g98 ( .A(n_92), .Y(n_98) );
INVx1_ASAP7_75t_L g162 ( .A(n_92), .Y(n_162) );
INVx2_ASAP7_75t_L g123 ( .A(n_94), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_94), .A2(n_144), .B1(n_145), .B2(n_146), .Y(n_143) );
OAI22xp5_ASAP7_75t_L g181 ( .A1(n_94), .A2(n_145), .B1(n_182), .B2(n_183), .Y(n_181) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx3_ASAP7_75t_L g100 ( .A(n_95), .Y(n_100) );
INVx1_ASAP7_75t_L g119 ( .A(n_95), .Y(n_119) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_95), .Y(n_139) );
INVx1_ASAP7_75t_L g388 ( .A(n_95), .Y(n_388) );
INVx2_ASAP7_75t_L g156 ( .A(n_97), .Y(n_156) );
INVx3_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx3_ASAP7_75t_L g131 ( .A(n_99), .Y(n_131) );
INVx5_ASAP7_75t_L g134 ( .A(n_100), .Y(n_134) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_102), .A2(n_114), .B(n_124), .Y(n_113) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_102), .A2(n_129), .B(n_140), .Y(n_128) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_104), .Y(n_102) );
AND2x2_ASAP7_75t_L g111 ( .A(n_103), .B(n_104), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
NAND3xp33_ASAP7_75t_L g180 ( .A(n_107), .B(n_181), .C(n_184), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_107), .A2(n_193), .B(n_196), .Y(n_192) );
AND2x2_ASAP7_75t_L g386 ( .A(n_107), .B(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI21xp5_ASAP7_75t_L g114 ( .A1(n_108), .A2(n_115), .B(n_120), .Y(n_114) );
OAI21xp5_ASAP7_75t_L g129 ( .A1(n_108), .A2(n_130), .B(n_135), .Y(n_129) );
OAI21xp5_ASAP7_75t_L g153 ( .A1(n_108), .A2(n_154), .B(n_159), .Y(n_153) );
OAI21xp5_ASAP7_75t_L g167 ( .A1(n_108), .A2(n_168), .B(n_171), .Y(n_167) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_109), .Y(n_492) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_110), .A2(n_167), .B(n_174), .Y(n_166) );
INVx4_ASAP7_75t_L g184 ( .A(n_110), .Y(n_184) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_125), .Y(n_112) );
AND2x2_ASAP7_75t_L g187 ( .A(n_113), .B(n_141), .Y(n_187) );
INVx2_ASAP7_75t_L g221 ( .A(n_113), .Y(n_221) );
AND2x2_ASAP7_75t_L g236 ( .A(n_113), .B(n_142), .Y(n_236) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_113), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_113), .B(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g256 ( .A(n_113), .B(n_219), .Y(n_256) );
INVx1_ASAP7_75t_L g268 ( .A(n_113), .Y(n_268) );
INVx1_ASAP7_75t_L g309 ( .A(n_113), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_113), .B(n_209), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_117), .B(n_118), .Y(n_115) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B(n_123), .Y(n_120) );
O2A1O1Ixp5_ASAP7_75t_L g196 ( .A1(n_123), .A2(n_160), .B(n_197), .C(n_198), .Y(n_196) );
NOR2xp67_ASAP7_75t_L g125 ( .A(n_126), .B(n_141), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g186 ( .A(n_127), .B(n_187), .Y(n_186) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_127), .Y(n_214) );
AND2x2_ASAP7_75t_SL g267 ( .A(n_127), .B(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g271 ( .A(n_127), .B(n_141), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_127), .B(n_266), .Y(n_329) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g219 ( .A(n_128), .Y(n_219) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_128), .Y(n_235) );
OR2x2_ASAP7_75t_L g308 ( .A(n_128), .B(n_309), .Y(n_308) );
O2A1O1Ixp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_132), .B(n_133), .C(n_134), .Y(n_130) );
INVx2_ASAP7_75t_L g145 ( .A(n_134), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_134), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_134), .A2(n_194), .B(n_195), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g158 ( .A(n_138), .Y(n_158) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx2_ASAP7_75t_L g215 ( .A(n_142), .Y(n_215) );
AND2x2_ASAP7_75t_L g220 ( .A(n_142), .B(n_221), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g159 ( .A1(n_145), .A2(n_160), .B(n_163), .C(n_164), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_145), .A2(n_172), .B(n_173), .Y(n_171) );
INVx2_ASAP7_75t_L g152 ( .A(n_147), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_148), .B(n_203), .Y(n_366) );
INVx1_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g336 ( .A(n_149), .B(n_177), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_166), .Y(n_149) );
AND2x2_ASAP7_75t_L g212 ( .A(n_150), .B(n_203), .Y(n_212) );
INVx2_ASAP7_75t_L g224 ( .A(n_150), .Y(n_224) );
AND2x2_ASAP7_75t_L g258 ( .A(n_150), .B(n_206), .Y(n_258) );
AND2x2_ASAP7_75t_L g325 ( .A(n_150), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_151), .B(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g205 ( .A(n_151), .B(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g245 ( .A(n_151), .B(n_166), .Y(n_245) );
AND2x2_ASAP7_75t_L g262 ( .A(n_151), .B(n_263), .Y(n_262) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_165), .Y(n_151) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_152), .A2(n_192), .B(n_199), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_157), .C(n_158), .Y(n_154) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_163), .A2(n_499), .B1(n_513), .B2(n_521), .Y(n_530) );
AND2x2_ASAP7_75t_L g188 ( .A(n_166), .B(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g206 ( .A(n_166), .Y(n_206) );
AND2x2_ASAP7_75t_L g211 ( .A(n_166), .B(n_191), .Y(n_211) );
AND2x2_ASAP7_75t_L g284 ( .A(n_166), .B(n_263), .Y(n_284) );
AND2x2_ASAP7_75t_L g349 ( .A(n_166), .B(n_339), .Y(n_349) );
OAI311xp33_ASAP7_75t_L g232 ( .A1(n_175), .A2(n_233), .A3(n_237), .B1(n_239), .C1(n_259), .Y(n_232) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g244 ( .A(n_176), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g303 ( .A(n_176), .B(n_211), .Y(n_303) );
AND2x2_ASAP7_75t_L g377 ( .A(n_176), .B(n_258), .Y(n_377) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_177), .B(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g312 ( .A(n_177), .Y(n_312) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx3_ASAP7_75t_L g203 ( .A(n_178), .Y(n_203) );
NOR2x1_ASAP7_75t_L g275 ( .A(n_178), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g332 ( .A(n_178), .B(n_206), .Y(n_332) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx1_ASAP7_75t_L g229 ( .A(n_179), .Y(n_229) );
AO21x1_ASAP7_75t_L g228 ( .A1(n_181), .A2(n_184), .B(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g207 ( .A(n_187), .B(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g260 ( .A(n_187), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g340 ( .A(n_187), .B(n_341), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g239 ( .A1(n_188), .A2(n_220), .B1(n_240), .B2(n_244), .C(n_246), .Y(n_239) );
INVx1_ASAP7_75t_L g364 ( .A(n_189), .Y(n_364) );
OR2x2_ASAP7_75t_L g330 ( .A(n_190), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g225 ( .A(n_191), .B(n_206), .Y(n_225) );
OR2x2_ASAP7_75t_L g227 ( .A(n_191), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g252 ( .A(n_191), .Y(n_252) );
INVx2_ASAP7_75t_L g263 ( .A(n_191), .Y(n_263) );
AND2x2_ASAP7_75t_L g290 ( .A(n_191), .B(n_228), .Y(n_290) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_191), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_207), .B1(n_210), .B2(n_213), .C(n_216), .Y(n_200) );
INVx1_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
AND2x2_ASAP7_75t_L g301 ( .A(n_203), .B(n_211), .Y(n_301) );
AND2x2_ASAP7_75t_L g351 ( .A(n_203), .B(n_205), .Y(n_351) );
INVx2_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g238 ( .A(n_205), .B(n_209), .Y(n_238) );
AND2x2_ASAP7_75t_L g317 ( .A(n_205), .B(n_290), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_206), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g276 ( .A(n_206), .Y(n_276) );
OAI21xp33_ASAP7_75t_L g286 ( .A1(n_207), .A2(n_287), .B(n_289), .Y(n_286) );
OR2x2_ASAP7_75t_L g230 ( .A(n_208), .B(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g296 ( .A(n_208), .B(n_256), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_208), .B(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g273 ( .A(n_209), .B(n_242), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_209), .B(n_356), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_210), .B(n_236), .Y(n_346) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
AND2x2_ASAP7_75t_L g269 ( .A(n_211), .B(n_224), .Y(n_269) );
INVx1_ASAP7_75t_L g285 ( .A(n_212), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_222), .B1(n_226), .B2(n_230), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g248 ( .A(n_219), .Y(n_248) );
INVx1_ASAP7_75t_L g261 ( .A(n_219), .Y(n_261) );
INVx1_ASAP7_75t_L g231 ( .A(n_220), .Y(n_231) );
AND2x2_ASAP7_75t_L g302 ( .A(n_220), .B(n_248), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_220), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_225), .Y(n_222) );
OR2x2_ASAP7_75t_L g226 ( .A(n_223), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_223), .B(n_339), .Y(n_338) );
NOR2xp67_ASAP7_75t_L g370 ( .A(n_223), .B(n_371), .Y(n_370) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g373 ( .A(n_225), .B(n_325), .Y(n_373) );
INVx1_ASAP7_75t_SL g339 ( .A(n_227), .Y(n_339) );
AND2x2_ASAP7_75t_L g279 ( .A(n_228), .B(n_263), .Y(n_279) );
INVx1_ASAP7_75t_L g326 ( .A(n_228), .Y(n_326) );
OAI222xp33_ASAP7_75t_L g367 ( .A1(n_233), .A2(n_323), .B1(n_368), .B2(n_369), .C1(n_372), .C2(n_374), .Y(n_367) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
INVx1_ASAP7_75t_L g288 ( .A(n_235), .Y(n_288) );
AND2x2_ASAP7_75t_L g299 ( .A(n_236), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_236), .B(n_341), .Y(n_368) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_238), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g343 ( .A(n_240), .Y(n_343) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_SL g281 ( .A(n_243), .Y(n_281) );
AND2x2_ASAP7_75t_L g360 ( .A(n_243), .B(n_321), .Y(n_360) );
AND2x2_ASAP7_75t_L g383 ( .A(n_243), .B(n_267), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_245), .B(n_279), .Y(n_278) );
OAI32xp33_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .A3(n_251), .B1(n_253), .B2(n_257), .Y(n_246) );
BUFx2_ASAP7_75t_L g321 ( .A(n_248), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_249), .B(n_267), .Y(n_348) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g287 ( .A(n_250), .B(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g355 ( .A(n_250), .B(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g344 ( .A(n_251), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g315 ( .A(n_254), .B(n_288), .Y(n_315) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OAI221xp5_ASAP7_75t_SL g277 ( .A1(n_256), .A2(n_278), .B1(n_280), .B2(n_282), .C(n_286), .Y(n_277) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g289 ( .A(n_258), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g295 ( .A(n_258), .B(n_279), .Y(n_295) );
AOI221xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_262), .B1(n_264), .B2(n_269), .C(n_270), .Y(n_259) );
INVx1_ASAP7_75t_L g378 ( .A(n_260), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_261), .B(n_355), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g274 ( .A(n_262), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_267), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g333 ( .A(n_267), .Y(n_333) );
BUFx3_ASAP7_75t_L g356 ( .A(n_268), .Y(n_356) );
INVx1_ASAP7_75t_SL g297 ( .A(n_269), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_269), .B(n_311), .Y(n_310) );
AOI21xp33_ASAP7_75t_SL g270 ( .A1(n_271), .A2(n_272), .B(n_274), .Y(n_270) );
OAI221xp5_ASAP7_75t_L g375 ( .A1(n_271), .A2(n_372), .B1(n_376), .B2(n_378), .C(n_379), .Y(n_375) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g318 ( .A(n_276), .B(n_279), .Y(n_318) );
INVx1_ASAP7_75t_L g382 ( .A(n_276), .Y(n_382) );
INVx2_ASAP7_75t_L g371 ( .A(n_279), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_279), .B(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g324 ( .A(n_284), .B(n_325), .Y(n_324) );
OAI221xp5_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_294), .B1(n_296), .B2(n_297), .C(n_298), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_301), .B1(n_302), .B2(n_303), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_300), .A2(n_362), .B1(n_363), .B2(n_365), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_303), .A2(n_380), .B(n_383), .Y(n_379) );
NOR4xp25_ASAP7_75t_SL g304 ( .A(n_305), .B(n_313), .C(n_322), .D(n_342), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_310), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B1(n_319), .B2(n_320), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g358 ( .A(n_318), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_327), .B1(n_330), .B2(n_333), .C(n_334), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g345 ( .A(n_325), .Y(n_345) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI21xp5_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_337), .B(n_340), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI211xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B(n_346), .C(n_347), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_350), .B2(n_351), .Y(n_347) );
CKINVDCx14_ASAP7_75t_R g357 ( .A(n_351), .Y(n_357) );
NOR3xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_367), .C(n_375), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .B1(n_358), .B2(n_359), .C(n_361), .Y(n_353) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
CKINVDCx16_ASAP7_75t_R g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_385), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_386), .Y(n_385) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_387), .A2(n_491), .B(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_390), .Y(n_389) );
OAI322xp33_ASAP7_75t_L g495 ( .A1(n_391), .A2(n_496), .A3(n_497), .B1(n_525), .B2(n_526), .C1(n_529), .C2(n_530), .Y(n_495) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_451), .Y(n_392) );
INVxp67_ASAP7_75t_L g525 ( .A(n_393), .Y(n_525) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_418), .C(n_438), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_412), .B2(n_413), .Y(n_394) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_407), .Y(n_398) );
INVx2_ASAP7_75t_L g477 ( .A(n_399), .Y(n_477) );
OR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_405), .Y(n_399) );
AND2x2_ASAP7_75t_L g417 ( .A(n_400), .B(n_405), .Y(n_417) );
AND2x2_ASAP7_75t_L g458 ( .A(n_400), .B(n_437), .Y(n_458) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g421 ( .A(n_401), .B(n_405), .Y(n_421) );
AND2x2_ASAP7_75t_L g431 ( .A(n_401), .B(n_411), .Y(n_431) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_404), .Y(n_406) );
INVx2_ASAP7_75t_L g437 ( .A(n_405), .Y(n_437) );
INVx1_ASAP7_75t_L g471 ( .A(n_405), .Y(n_471) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_408), .B(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g480 ( .A(n_408), .B(n_458), .Y(n_480) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g423 ( .A(n_409), .Y(n_423) );
INVx1_ASAP7_75t_L g430 ( .A(n_409), .Y(n_430) );
INVx1_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_409), .B(n_411), .Y(n_462) );
AND2x2_ASAP7_75t_L g422 ( .A(n_410), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g468 ( .A(n_411), .B(n_450), .Y(n_468) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g467 ( .A(n_417), .B(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g483 ( .A(n_417), .B(n_422), .Y(n_483) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_424), .B1(n_425), .B2(n_432), .C(n_433), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x6_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g447 ( .A(n_421), .Y(n_447) );
AND2x2_ASAP7_75t_L g457 ( .A(n_422), .B(n_458), .Y(n_457) );
AND2x6_ASAP7_75t_L g476 ( .A(n_422), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g436 ( .A(n_430), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g435 ( .A(n_431), .B(n_436), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g441 ( .A(n_431), .B(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g442 ( .A(n_437), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B1(n_443), .B2(n_444), .Y(n_438) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
CKINVDCx16_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
OR2x6_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVxp67_ASAP7_75t_L g496 ( .A(n_451), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_472), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_463), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g460 ( .A(n_458), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g486 ( .A(n_458), .B(n_468), .Y(n_486) );
BUFx2_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x6_ASAP7_75t_L g470 ( .A(n_462), .B(n_471), .Y(n_470) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx4_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx8_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_481), .Y(n_472) );
INVx2_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
INVx11_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx4f_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_SL g489 ( .A(n_490), .B(n_493), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND3x1_ASAP7_75t_SL g513 ( .A(n_491), .B(n_493), .C(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g521 ( .A(n_491), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_492), .B(n_494), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_503), .B1(n_509), .B2(n_510), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_500), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_503), .Y(n_510) );
INVx1_ASAP7_75t_L g508 ( .A(n_505), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
INVxp67_ASAP7_75t_L g524 ( .A(n_514), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
endmodule