module fake_jpeg_26146_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_42),
.Y(n_49)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_29),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_53),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_19),
.B1(n_32),
.B2(n_20),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_41),
.B1(n_36),
.B2(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_20),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_19),
.B1(n_32),
.B2(n_20),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_38),
.B1(n_28),
.B2(n_43),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_19),
.B1(n_32),
.B2(n_25),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_40),
.B1(n_36),
.B2(n_41),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_59),
.Y(n_89)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_64),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_65),
.B(n_91),
.Y(n_127)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_69),
.A2(n_71),
.B1(n_92),
.B2(n_57),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_36),
.B1(n_41),
.B2(n_40),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_77),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_74),
.A2(n_94),
.B1(n_21),
.B2(n_50),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_78),
.B1(n_86),
.B2(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_28),
.B1(n_38),
.B2(n_43),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_24),
.B1(n_16),
.B2(n_26),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_84),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_81),
.B(n_95),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_35),
.C(n_29),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_33),
.C(n_30),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_30),
.B1(n_17),
.B2(n_33),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_21),
.B1(n_26),
.B2(n_59),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_16),
.B1(n_24),
.B2(n_30),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_50),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_50),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_28),
.B1(n_37),
.B2(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_37),
.B1(n_31),
.B2(n_27),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_93),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_16),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_98),
.Y(n_119)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_58),
.B(n_37),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_31),
.B(n_27),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_101),
.A2(n_115),
.B(n_117),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_27),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_126),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_108),
.B1(n_114),
.B2(n_123),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_12),
.C(n_11),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_15),
.B(n_12),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_68),
.A2(n_37),
.B1(n_57),
.B2(n_48),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_21),
.B(n_26),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_64),
.A2(n_22),
.B(n_34),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_35),
.B(n_59),
.C(n_50),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_122),
.B(n_90),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_33),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_67),
.A2(n_59),
.B1(n_30),
.B2(n_33),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_63),
.B1(n_69),
.B2(n_71),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_134),
.B1(n_147),
.B2(n_109),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_65),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_141),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_65),
.B1(n_75),
.B2(n_78),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_89),
.B(n_91),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_142),
.B(n_156),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_84),
.B1(n_97),
.B2(n_81),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_136),
.A2(n_143),
.B(n_150),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_96),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_138),
.B(n_139),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_87),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_140),
.B(n_151),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_98),
.Y(n_141)
);

OAI22x1_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_35),
.B1(n_22),
.B2(n_34),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_144),
.A2(n_156),
.B1(n_149),
.B2(n_66),
.Y(n_166)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_148),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_111),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_77),
.B1(n_66),
.B2(n_76),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_112),
.A2(n_92),
.B(n_1),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_111),
.B(n_72),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_155),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_72),
.Y(n_155)
);

OR2x4_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_22),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_110),
.B(n_17),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_106),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_158),
.Y(n_178)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_169),
.B1(n_131),
.B2(n_154),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_167),
.B(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_182),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_121),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_170),
.B(n_188),
.Y(n_221)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_172),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_122),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_122),
.C(n_126),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_190),
.C(n_0),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_149),
.B(n_135),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_180),
.A2(n_143),
.B(n_127),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_158),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_181),
.Y(n_194)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_102),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_192),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_186),
.B(n_187),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_125),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_127),
.C(n_117),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_153),
.B(n_101),
.Y(n_192)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_208),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_199),
.B1(n_205),
.B2(n_218),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_132),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_222),
.C(n_217),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_133),
.B1(n_134),
.B2(n_150),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_162),
.B(n_178),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_115),
.Y(n_204)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_174),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_133),
.B1(n_128),
.B2(n_107),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_125),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_108),
.B1(n_123),
.B2(n_114),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_218),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_172),
.B1(n_185),
.B2(n_164),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_120),
.B1(n_124),
.B2(n_152),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_124),
.Y(n_214)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

OAI221xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_15),
.B1(n_9),
.B2(n_7),
.C(n_10),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_120),
.B1(n_17),
.B2(n_23),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_180),
.A2(n_23),
.B1(n_34),
.B2(n_2),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_203),
.B1(n_221),
.B2(n_193),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_SL g220 ( 
.A1(n_165),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_220)
);

AO22x2_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_223),
.B(n_231),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_238),
.B1(n_210),
.B2(n_212),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_197),
.A2(n_190),
.B1(n_174),
.B2(n_163),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_228),
.A2(n_215),
.B1(n_219),
.B2(n_195),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_201),
.Y(n_249)
);

AOI221x1_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_189),
.B1(n_162),
.B2(n_183),
.C(n_165),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_236),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_181),
.C(n_178),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_240),
.C(n_222),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_200),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_206),
.A2(n_173),
.B(n_161),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_244),
.B(n_243),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_202),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_10),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_173),
.C(n_171),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_7),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_220),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_220),
.B1(n_4),
.B2(n_5),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_194),
.B(n_2),
.Y(n_244)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_245),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_240),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_247),
.A2(n_264),
.B1(n_257),
.B2(n_261),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_248),
.A2(n_263),
.B1(n_224),
.B2(n_243),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_258),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_244),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_252),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_202),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_257),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_209),
.C(n_206),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_261),
.C(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_244),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_259),
.B(n_265),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_193),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_196),
.C(n_220),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_254),
.B(n_225),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_267),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_270),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_223),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_249),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_276),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_238),
.B1(n_234),
.B2(n_227),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_13),
.B1(n_14),
.B2(n_5),
.Y(n_294)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_228),
.Y(n_276)
);

XOR2x2_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_224),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_243),
.B(n_13),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_232),
.C(n_241),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_279),
.A2(n_264),
.B(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_269),
.B(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_270),
.C(n_276),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_278),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_266),
.B(n_263),
.Y(n_290)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_3),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_13),
.C(n_14),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_272),
.C(n_268),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_294),
.A2(n_4),
.B1(n_5),
.B2(n_285),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_302),
.C(n_284),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_298),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_299),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_277),
.B1(n_272),
.B2(n_271),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_4),
.B1(n_5),
.B2(n_288),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_4),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_289),
.B(n_293),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_309),
.B(n_299),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_287),
.B(n_284),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_307),
.A2(n_298),
.B(n_303),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_306),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_282),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_295),
.C(n_282),
.Y(n_312)
);

INVx11_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_317),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_314),
.A2(n_316),
.B(n_309),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_315),
.B(n_316),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_318),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_312),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);


endmodule