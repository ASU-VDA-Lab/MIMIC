module fake_netlist_5_1419_n_777 (n_137, n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_777);

input n_137;
input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_777;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_139;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_443;
wire n_372;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_568;
wire n_509;
wire n_147;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_138;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_681;
wire n_584;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_142;
wire n_743;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_144;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_679;
wire n_707;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_728;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_34),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_0),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_37),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_1),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_60),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_59),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_92),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_109),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_15),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_35),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_105),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_75),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_128),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_57),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_113),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_110),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_68),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_63),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_49),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_125),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_78),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_38),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_16),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_71),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_58),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_65),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_72),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_30),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_39),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_66),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_24),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_13),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_L g189 ( 
.A(n_52),
.B(n_94),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_41),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_69),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_74),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_129),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_81),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_0),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_1),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_139),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_142),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_144),
.A2(n_2),
.B(n_3),
.Y(n_208)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_148),
.B(n_21),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_163),
.Y(n_214)
);

BUFx8_ASAP7_75t_SL g215 ( 
.A(n_194),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_188),
.Y(n_218)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_165),
.A2(n_4),
.B(n_5),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_147),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_144),
.Y(n_225)
);

BUFx8_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_153),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_155),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_156),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_183),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_215),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_224),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_202),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_235),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g245 ( 
.A(n_235),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_202),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_237),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_195),
.B(n_157),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_R g255 ( 
.A(n_218),
.B(n_143),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_234),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_203),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_198),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_218),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_R g265 ( 
.A(n_214),
.B(n_149),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_205),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_210),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_235),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_210),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_235),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_197),
.B(n_158),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_205),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_205),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_211),
.B(n_159),
.Y(n_275)
);

AO22x2_ASAP7_75t_L g276 ( 
.A1(n_232),
.A2(n_189),
.B1(n_6),
.B2(n_7),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_211),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_216),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_L g279 ( 
.A(n_211),
.B(n_160),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_229),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_226),
.Y(n_281)
);

OR2x2_ASAP7_75t_SL g282 ( 
.A(n_208),
.B(n_200),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_198),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_226),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_225),
.B(n_199),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_201),
.B(n_162),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

NOR3xp33_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_219),
.C(n_169),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_254),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_259),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_164),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_255),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_243),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_239),
.B(n_198),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_206),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_209),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_265),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_274),
.B(n_180),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_206),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_263),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_225),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_244),
.B(n_206),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_206),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_206),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_207),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_285),
.A2(n_209),
.B1(n_171),
.B2(n_185),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_250),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_207),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_207),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_SL g316 ( 
.A(n_284),
.B(n_208),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_275),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_268),
.B(n_207),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_253),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_225),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_268),
.B(n_207),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_261),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_277),
.B(n_166),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_256),
.B(n_174),
.Y(n_325)
);

NAND2xp33_ASAP7_75t_L g326 ( 
.A(n_257),
.B(n_209),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_241),
.B(n_175),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_213),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_261),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_246),
.B(n_249),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_261),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_251),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_266),
.A2(n_219),
.B(n_220),
.C(n_196),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_276),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_267),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_281),
.A2(n_230),
.B(n_212),
.C(n_196),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_269),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_264),
.B(n_213),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_238),
.B(n_177),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_240),
.B(n_178),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_242),
.B(n_213),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_248),
.B(n_213),
.Y(n_344)
);

NAND3xp33_ASAP7_75t_L g345 ( 
.A(n_260),
.B(n_213),
.C(n_228),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_244),
.B(n_221),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_244),
.B(n_221),
.Y(n_348)
);

AND3x1_ASAP7_75t_L g349 ( 
.A(n_272),
.B(n_230),
.C(n_220),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_L g350 ( 
.A(n_270),
.B(n_209),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_244),
.B(n_221),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_255),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_289),
.A2(n_209),
.B1(n_208),
.B2(n_226),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_290),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_287),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_309),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_304),
.B(n_209),
.Y(n_358)
);

NOR3xp33_ASAP7_75t_SL g359 ( 
.A(n_343),
.B(n_181),
.C(n_186),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

AND2x6_ASAP7_75t_L g361 ( 
.A(n_290),
.B(n_204),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_228),
.B1(n_223),
.B2(n_222),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_187),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_304),
.B(n_221),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_346),
.B(n_221),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_R g366 ( 
.A(n_299),
.B(n_192),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_318),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_294),
.Y(n_368)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_312),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_303),
.Y(n_371)
);

BUFx6f_ASAP7_75t_SL g372 ( 
.A(n_337),
.Y(n_372)
);

BUFx6f_ASAP7_75t_SL g373 ( 
.A(n_333),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_193),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_320),
.Y(n_375)
);

NAND2x1p5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_222),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_320),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_22),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_340),
.B(n_344),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_352),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_313),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_222),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_340),
.B(n_222),
.Y(n_383)
);

HB1xp67_ASAP7_75t_SL g384 ( 
.A(n_330),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_222),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_307),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_334),
.A2(n_217),
.B(n_212),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_L g388 ( 
.A(n_317),
.B(n_223),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_348),
.B(n_223),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_321),
.B(n_293),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_349),
.A2(n_228),
.B1(n_223),
.B2(n_217),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_295),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_339),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_310),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_292),
.A2(n_228),
.B1(n_223),
.B2(n_204),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_295),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_302),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_324),
.B(n_228),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_302),
.Y(n_400)
);

O2A1O1Ixp33_ASAP7_75t_L g401 ( 
.A1(n_332),
.A2(n_338),
.B(n_335),
.C(n_336),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g402 ( 
.A(n_332),
.B(n_23),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_312),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_345),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_348),
.B(n_25),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_300),
.B(n_5),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_351),
.B(n_26),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_351),
.B(n_27),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_308),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_311),
.B(n_6),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_288),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_331),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_297),
.B(n_28),
.Y(n_417)
);

OAI221xp5_ASAP7_75t_L g418 ( 
.A1(n_301),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_306),
.B(n_29),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_326),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_325),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_331),
.Y(n_422)
);

OAI21xp33_ASAP7_75t_L g423 ( 
.A1(n_408),
.A2(n_327),
.B(n_341),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_360),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_379),
.B(n_342),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_386),
.A2(n_350),
.B(n_298),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_378),
.B(n_421),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_395),
.A2(n_296),
.B(n_314),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_387),
.A2(n_323),
.B(n_322),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_316),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_378),
.B(n_319),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_388),
.A2(n_328),
.B(n_93),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_371),
.B(n_12),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_407),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_367),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_415),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_392),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_397),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_380),
.B(n_31),
.Y(n_439)
);

NAND2x1p5_ASAP7_75t_L g440 ( 
.A(n_354),
.B(n_32),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_369),
.A2(n_96),
.B(n_136),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_369),
.A2(n_95),
.B(n_135),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_357),
.Y(n_443)
);

O2A1O1Ixp33_ASAP7_75t_L g444 ( 
.A1(n_401),
.A2(n_14),
.B(n_16),
.C(n_17),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_354),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_353),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_446)
);

O2A1O1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_414),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_394),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_420),
.A2(n_20),
.B1(n_33),
.B2(n_36),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_369),
.A2(n_40),
.B(n_42),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_418),
.A2(n_362),
.B1(n_384),
.B2(n_405),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_370),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_361),
.B(n_385),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_363),
.B(n_43),
.C(n_44),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_355),
.B(n_45),
.Y(n_455)
);

O2A1O1Ixp5_ASAP7_75t_SL g456 ( 
.A1(n_383),
.A2(n_375),
.B(n_377),
.C(n_413),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_407),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_361),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_361),
.B(n_50),
.Y(n_459)
);

A2O1A1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_399),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_361),
.B(n_55),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_393),
.A2(n_56),
.B(n_62),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_356),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_412),
.Y(n_464)
);

BUFx12f_ASAP7_75t_L g465 ( 
.A(n_390),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_398),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_374),
.B(n_64),
.Y(n_467)
);

A2O1A1Ixp33_ASAP7_75t_L g468 ( 
.A1(n_381),
.A2(n_67),
.B(n_73),
.C(n_76),
.Y(n_468)
);

O2A1O1Ixp33_ASAP7_75t_SL g469 ( 
.A1(n_417),
.A2(n_77),
.B(n_80),
.C(n_82),
.Y(n_469)
);

BUFx12f_ASAP7_75t_L g470 ( 
.A(n_390),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_412),
.Y(n_472)
);

NAND2x1p5_ASAP7_75t_L g473 ( 
.A(n_393),
.B(n_83),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_393),
.A2(n_84),
.B(n_85),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_368),
.B(n_86),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_359),
.B(n_88),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_373),
.B(n_89),
.Y(n_477)
);

NAND3xp33_ASAP7_75t_SL g478 ( 
.A(n_366),
.B(n_90),
.C(n_91),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_358),
.A2(n_97),
.B(n_98),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_419),
.A2(n_99),
.B(n_101),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_403),
.B(n_103),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_434),
.Y(n_482)
);

OAI21x1_ASAP7_75t_SL g483 ( 
.A1(n_444),
.A2(n_410),
.B(n_409),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_429),
.A2(n_406),
.B(n_365),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_465),
.Y(n_486)
);

OAI21x1_ASAP7_75t_SL g487 ( 
.A1(n_459),
.A2(n_364),
.B(n_382),
.Y(n_487)
);

AO21x2_ASAP7_75t_L g488 ( 
.A1(n_453),
.A2(n_389),
.B(n_396),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_466),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_434),
.Y(n_491)
);

INVx5_ASAP7_75t_L g492 ( 
.A(n_464),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_426),
.A2(n_422),
.B(n_416),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_448),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_473),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_471),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_424),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_475),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_456),
.A2(n_428),
.B(n_453),
.Y(n_499)
);

AOI22x1_ASAP7_75t_L g500 ( 
.A1(n_479),
.A2(n_443),
.B1(n_452),
.B2(n_435),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_464),
.Y(n_501)
);

BUFx2_ASAP7_75t_SL g502 ( 
.A(n_457),
.Y(n_502)
);

BUFx2_ASAP7_75t_SL g503 ( 
.A(n_472),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_437),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_445),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_473),
.Y(n_506)
);

NAND2x1p5_ASAP7_75t_L g507 ( 
.A(n_431),
.B(n_404),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_433),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_432),
.A2(n_376),
.B(n_391),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_476),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_438),
.Y(n_511)
);

CKINVDCx6p67_ASAP7_75t_R g512 ( 
.A(n_439),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_430),
.Y(n_513)
);

AOI22x1_ASAP7_75t_L g514 ( 
.A1(n_440),
.A2(n_404),
.B1(n_403),
.B2(n_402),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_440),
.Y(n_515)
);

INVx8_ASAP7_75t_L g516 ( 
.A(n_476),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_427),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_459),
.A2(n_461),
.B(n_455),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_461),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_477),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_447),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_467),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_425),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_449),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_480),
.A2(n_402),
.B(n_404),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_451),
.A2(n_402),
.B(n_403),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_441),
.A2(n_402),
.B(n_106),
.Y(n_527)
);

CKINVDCx6p67_ASAP7_75t_R g528 ( 
.A(n_481),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_446),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_469),
.Y(n_530)
);

CKINVDCx14_ASAP7_75t_R g531 ( 
.A(n_478),
.Y(n_531)
);

OAI21x1_ASAP7_75t_SL g532 ( 
.A1(n_526),
.A2(n_446),
.B(n_449),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_495),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_517),
.B(n_511),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_485),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_524),
.A2(n_436),
.B1(n_423),
.B2(n_451),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_511),
.Y(n_537)
);

AO21x1_ASAP7_75t_L g538 ( 
.A1(n_519),
.A2(n_436),
.B(n_474),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_524),
.A2(n_373),
.B1(n_458),
.B2(n_372),
.Y(n_539)
);

INVx3_ASAP7_75t_SL g540 ( 
.A(n_516),
.Y(n_540)
);

BUFx2_ASAP7_75t_R g541 ( 
.A(n_486),
.Y(n_541)
);

AO21x1_ASAP7_75t_L g542 ( 
.A1(n_519),
.A2(n_462),
.B(n_450),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_501),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_494),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_529),
.B(n_460),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_494),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_505),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_531),
.A2(n_372),
.B1(n_454),
.B2(n_442),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_501),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_482),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_498),
.Y(n_551)
);

AO21x2_ASAP7_75t_L g552 ( 
.A1(n_487),
.A2(n_483),
.B(n_499),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_523),
.A2(n_468),
.B1(n_107),
.B2(n_108),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_486),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_489),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_496),
.Y(n_556)
);

CKINVDCx11_ASAP7_75t_R g557 ( 
.A(n_490),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_497),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_504),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_491),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_490),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_492),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_491),
.Y(n_563)
);

NAND2x1p5_ASAP7_75t_L g564 ( 
.A(n_495),
.B(n_104),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_482),
.Y(n_565)
);

OAI21x1_ASAP7_75t_L g566 ( 
.A1(n_493),
.A2(n_111),
.B(n_114),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_495),
.Y(n_567)
);

CKINVDCx11_ASAP7_75t_R g568 ( 
.A(n_520),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g569 ( 
.A1(n_493),
.A2(n_115),
.B(n_118),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_521),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_482),
.Y(n_571)
);

A2O1A1Ixp33_ASAP7_75t_L g572 ( 
.A1(n_536),
.A2(n_523),
.B(n_513),
.C(n_516),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_554),
.B(n_516),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_539),
.A2(n_508),
.B(n_520),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_R g575 ( 
.A(n_545),
.B(n_530),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_R g576 ( 
.A(n_545),
.B(n_530),
.Y(n_576)
);

OAI22xp33_ASAP7_75t_L g577 ( 
.A1(n_544),
.A2(n_510),
.B1(n_512),
.B2(n_517),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_R g578 ( 
.A(n_568),
.B(n_557),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_R g579 ( 
.A(n_554),
.B(n_561),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_546),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_547),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_551),
.B(n_505),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_534),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_R g584 ( 
.A(n_534),
.B(n_562),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_561),
.B(n_517),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_534),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_534),
.B(n_515),
.Y(n_587)
);

AND2x2_ASAP7_75t_SL g588 ( 
.A(n_553),
.B(n_495),
.Y(n_588)
);

NOR2x1p5_ASAP7_75t_L g589 ( 
.A(n_535),
.B(n_512),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_R g590 ( 
.A(n_540),
.B(n_516),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_R g591 ( 
.A(n_562),
.B(n_530),
.Y(n_591)
);

AND2x4_ASAP7_75t_SL g592 ( 
.A(n_533),
.B(n_506),
.Y(n_592)
);

A2O1A1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_548),
.A2(n_522),
.B(n_527),
.C(n_518),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_564),
.B(n_503),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_535),
.B(n_515),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_SL g596 ( 
.A1(n_555),
.A2(n_528),
.B(n_483),
.C(n_514),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_541),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_R g598 ( 
.A(n_540),
.B(n_528),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_559),
.B(n_503),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_555),
.A2(n_514),
.B1(n_502),
.B2(n_507),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_564),
.B(n_502),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_532),
.A2(n_522),
.B1(n_495),
.B2(n_506),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_556),
.B(n_506),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_564),
.B(n_506),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_559),
.B(n_506),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_540),
.B(n_556),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_533),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_533),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_532),
.A2(n_500),
.B1(n_487),
.B2(n_507),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_558),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_558),
.B(n_507),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_538),
.A2(n_500),
.B1(n_488),
.B2(n_518),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_537),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_537),
.Y(n_614)
);

AND2x4_ASAP7_75t_SL g615 ( 
.A(n_533),
.B(n_492),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_560),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_560),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_533),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_543),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_R g620 ( 
.A(n_562),
.B(n_525),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_611),
.B(n_552),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_610),
.Y(n_622)
);

OA21x2_ASAP7_75t_L g623 ( 
.A1(n_612),
.A2(n_499),
.B(n_484),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_583),
.B(n_552),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_616),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_617),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_588),
.A2(n_570),
.B1(n_538),
.B2(n_542),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_582),
.B(n_543),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_595),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g630 ( 
.A(n_575),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_613),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_586),
.B(n_552),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_614),
.B(n_549),
.Y(n_633)
);

INVx5_ASAP7_75t_L g634 ( 
.A(n_594),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_603),
.B(n_563),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_572),
.B(n_563),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_608),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_599),
.B(n_549),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_577),
.A2(n_570),
.B1(n_542),
.B2(n_550),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_585),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_574),
.B(n_565),
.Y(n_641)
);

NAND2x1p5_ASAP7_75t_L g642 ( 
.A(n_589),
.B(n_567),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_585),
.Y(n_643)
);

OA21x2_ASAP7_75t_L g644 ( 
.A1(n_593),
.A2(n_484),
.B(n_569),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_619),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_607),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_605),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_587),
.B(n_565),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_618),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_595),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_607),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_594),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_601),
.B(n_580),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_L g654 ( 
.A(n_581),
.B(n_571),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_601),
.B(n_488),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_609),
.B(n_488),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_604),
.B(n_569),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_600),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_621),
.B(n_587),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_625),
.Y(n_660)
);

OAI221xp5_ASAP7_75t_SL g661 ( 
.A1(n_627),
.A2(n_602),
.B1(n_573),
.B2(n_604),
.C(n_576),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_625),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_624),
.B(n_606),
.Y(n_663)
);

AND2x6_ASAP7_75t_SL g664 ( 
.A(n_641),
.B(n_578),
.Y(n_664)
);

NAND2x1_ASAP7_75t_SL g665 ( 
.A(n_658),
.B(n_591),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_621),
.B(n_566),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_634),
.B(n_573),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_626),
.B(n_592),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_634),
.B(n_598),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_634),
.B(n_567),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_637),
.B(n_597),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_631),
.B(n_567),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_631),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_628),
.B(n_579),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_645),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_622),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_638),
.B(n_596),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_655),
.B(n_567),
.Y(n_678)
);

NAND2x1_ASAP7_75t_L g679 ( 
.A(n_652),
.B(n_567),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_655),
.B(n_615),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_647),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_624),
.B(n_509),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_634),
.B(n_590),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_659),
.B(n_678),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_681),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_660),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_659),
.B(n_678),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_666),
.B(n_632),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_667),
.B(n_634),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_660),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_667),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_676),
.B(n_652),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_662),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_666),
.B(n_632),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_682),
.B(n_656),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_663),
.B(n_656),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_682),
.B(n_623),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_675),
.B(n_653),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_662),
.Y(n_699)
);

OAI33xp33_ASAP7_75t_L g700 ( 
.A1(n_698),
.A2(n_677),
.A3(n_653),
.B1(n_674),
.B2(n_673),
.B3(n_636),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_684),
.B(n_680),
.Y(n_701)
);

INVx3_ASAP7_75t_SL g702 ( 
.A(n_689),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_685),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_690),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_692),
.A2(n_630),
.B1(n_639),
.B2(n_584),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_685),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_694),
.B(n_663),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_694),
.B(n_673),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_R g709 ( 
.A1(n_697),
.A2(n_669),
.B(n_664),
.C(n_671),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_696),
.B(n_675),
.Y(n_710)
);

NAND2x1_ASAP7_75t_L g711 ( 
.A(n_689),
.B(n_667),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_711),
.B(n_689),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_703),
.B(n_665),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_706),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_710),
.Y(n_715)
);

INVxp67_ASAP7_75t_SL g716 ( 
.A(n_704),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_712),
.B(n_702),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_712),
.B(n_701),
.Y(n_718)
);

NOR2x1_ASAP7_75t_L g719 ( 
.A(n_713),
.B(n_709),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_713),
.A2(n_700),
.B1(n_705),
.B2(n_691),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_SL g721 ( 
.A1(n_719),
.A2(n_705),
.B(n_642),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_717),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_SL g723 ( 
.A1(n_720),
.A2(n_642),
.B(n_683),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_SL g724 ( 
.A(n_721),
.B(n_661),
.C(n_716),
.Y(n_724)
);

NOR3x1_ASAP7_75t_L g725 ( 
.A(n_723),
.B(n_679),
.C(n_707),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_724),
.B(n_722),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_725),
.A2(n_713),
.B1(n_718),
.B2(n_714),
.Y(n_727)
);

AOI221xp5_ASAP7_75t_L g728 ( 
.A1(n_724),
.A2(n_715),
.B1(n_704),
.B2(n_693),
.C(n_699),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_726),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_728),
.A2(n_668),
.B1(n_629),
.B2(n_679),
.Y(n_730)
);

NOR2x1_ASAP7_75t_L g731 ( 
.A(n_727),
.B(n_649),
.Y(n_731)
);

AO22x2_ASAP7_75t_L g732 ( 
.A1(n_726),
.A2(n_708),
.B1(n_686),
.B2(n_649),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_726),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_726),
.Y(n_734)
);

NOR3xp33_ASAP7_75t_SL g735 ( 
.A(n_733),
.B(n_734),
.C(n_729),
.Y(n_735)
);

NAND4xp75_ASAP7_75t_L g736 ( 
.A(n_731),
.B(n_654),
.C(n_668),
.D(n_651),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_732),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_730),
.B(n_687),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_734),
.A2(n_665),
.B(n_636),
.C(n_696),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_R g740 ( 
.A(n_733),
.B(n_123),
.Y(n_740)
);

AND3x2_ASAP7_75t_L g741 ( 
.A(n_734),
.B(n_670),
.C(n_687),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_740),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_737),
.Y(n_743)
);

NAND4xp25_ASAP7_75t_L g744 ( 
.A(n_739),
.B(n_650),
.C(n_640),
.D(n_680),
.Y(n_744)
);

OAI322xp33_ASAP7_75t_SL g745 ( 
.A1(n_735),
.A2(n_741),
.A3(n_736),
.B1(n_738),
.B2(n_690),
.C1(n_646),
.C2(n_688),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_738),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_740),
.Y(n_747)
);

O2A1O1Ixp5_ASAP7_75t_L g748 ( 
.A1(n_737),
.A2(n_670),
.B(n_646),
.C(n_684),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_746),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_742),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_SL g751 ( 
.A1(n_747),
.A2(n_670),
.B1(n_650),
.B2(n_640),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_743),
.Y(n_752)
);

INVxp67_ASAP7_75t_SL g753 ( 
.A(n_744),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_745),
.A2(n_629),
.B1(n_670),
.B2(n_643),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_748),
.Y(n_755)
);

NOR4xp25_ASAP7_75t_L g756 ( 
.A(n_743),
.B(n_635),
.C(n_657),
.D(n_672),
.Y(n_756)
);

AO22x2_ASAP7_75t_L g757 ( 
.A1(n_743),
.A2(n_657),
.B1(n_635),
.B2(n_672),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_746),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_749),
.A2(n_697),
.B1(n_643),
.B2(n_688),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_758),
.B(n_695),
.Y(n_760)
);

OAI31xp33_ASAP7_75t_L g761 ( 
.A1(n_755),
.A2(n_695),
.A3(n_648),
.B(n_638),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_752),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_750),
.B(n_648),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_753),
.A2(n_643),
.B1(n_620),
.B2(n_633),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_757),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_757),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_765),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_762),
.A2(n_754),
.B1(n_751),
.B2(n_756),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_766),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_760),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_SL g771 ( 
.A1(n_763),
.A2(n_643),
.B1(n_492),
.B2(n_644),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_769),
.A2(n_764),
.B1(n_759),
.B2(n_761),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_767),
.A2(n_633),
.B1(n_644),
.B2(n_623),
.Y(n_773)
);

NOR2xp67_ASAP7_75t_SL g774 ( 
.A(n_772),
.B(n_770),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_774),
.A2(n_768),
.B1(n_771),
.B2(n_773),
.Y(n_775)
);

NAND2x1p5_ASAP7_75t_L g776 ( 
.A(n_775),
.B(n_492),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_776),
.A2(n_492),
.B1(n_644),
.B2(n_623),
.Y(n_777)
);


endmodule