module fake_jpeg_7010_n_334 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_38),
.B(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_7),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_14),
.B(n_7),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_26),
.Y(n_61)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_53),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_54),
.B(n_58),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_33),
.B1(n_27),
.B2(n_32),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_57),
.A2(n_92),
.B1(n_100),
.B2(n_14),
.Y(n_107)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_50),
.Y(n_59)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_61),
.B(n_62),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_27),
.B1(n_15),
.B2(n_19),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_81),
.B1(n_86),
.B2(n_30),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_35),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

CKINVDCx6p67_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_27),
.B1(n_15),
.B2(n_31),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_69),
.A2(n_99),
.B(n_23),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_70),
.Y(n_124)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_26),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_83),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_15),
.B1(n_32),
.B2(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_28),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_88),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_28),
.C(n_18),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_16),
.C(n_17),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_35),
.B1(n_32),
.B2(n_31),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_38),
.B(n_34),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_97),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_16),
.B1(n_29),
.B2(n_23),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_49),
.B(n_24),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_96),
.B(n_102),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_29),
.B(n_23),
.C(n_22),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_38),
.B(n_34),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_101),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_48),
.A2(n_30),
.B1(n_24),
.B2(n_28),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_50),
.A2(n_16),
.B1(n_29),
.B2(n_23),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_19),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_19),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_100),
.A3(n_53),
.B1(n_59),
.B2(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_104),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_104),
.A2(n_76),
.B(n_81),
.C(n_68),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_30),
.B(n_14),
.C(n_16),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_129),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_107),
.A2(n_55),
.B1(n_78),
.B2(n_74),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_16),
.B(n_29),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_110),
.A2(n_87),
.B(n_89),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_125),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_16),
.C(n_17),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_85),
.C(n_66),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_64),
.A2(n_16),
.B(n_17),
.C(n_34),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_21),
.B(n_1),
.Y(n_167)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_135),
.B(n_139),
.Y(n_185)
);

AOI22x1_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_59),
.B1(n_76),
.B2(n_77),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_136),
.A2(n_132),
.B1(n_121),
.B2(n_116),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_141),
.B1(n_150),
.B2(n_151),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_106),
.C(n_130),
.Y(n_195)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_140),
.A2(n_156),
.B1(n_122),
.B2(n_124),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_107),
.A2(n_69),
.B1(n_99),
.B2(n_90),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_60),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_143),
.B(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_56),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_155),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_68),
.B(n_58),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_153),
.B(n_158),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_113),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_147),
.Y(n_172)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_129),
.A2(n_90),
.B1(n_52),
.B2(n_88),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_128),
.A2(n_75),
.B1(n_84),
.B2(n_94),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_87),
.B1(n_89),
.B2(n_21),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_161),
.B1(n_165),
.B2(n_116),
.Y(n_194)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_157),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_117),
.B(n_0),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_55),
.B(n_22),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_78),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_79),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_171),
.Y(n_196)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_111),
.B(n_9),
.Y(n_164)
);

XNOR2x1_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_13),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_105),
.A2(n_22),
.B1(n_21),
.B2(n_79),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_22),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_165),
.B(n_158),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_133),
.B(n_0),
.Y(n_171)
);

AND2x4_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_119),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_175),
.A2(n_176),
.B(n_181),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_167),
.A2(n_125),
.B(n_113),
.Y(n_176)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_180),
.Y(n_211)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_182),
.B(n_164),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_122),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_6),
.Y(n_226)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_203),
.B1(n_206),
.B2(n_169),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_170),
.B(n_124),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_191),
.B(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_194),
.A2(n_148),
.B1(n_152),
.B2(n_155),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_173),
.C(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_168),
.B(n_106),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_130),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_157),
.Y(n_214)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_134),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_204),
.Y(n_232)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_179),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_136),
.A2(n_121),
.B1(n_120),
.B2(n_112),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_141),
.A2(n_109),
.B(n_108),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_207),
.A2(n_181),
.B(n_173),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_148),
.A2(n_121),
.B1(n_108),
.B2(n_112),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_135),
.B1(n_209),
.B2(n_207),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_146),
.B(n_120),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_209),
.B(n_145),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_212),
.A2(n_221),
.B1(n_228),
.B2(n_239),
.Y(n_257)
);

A2O1A1O1Ixp25_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_161),
.B(n_159),
.C(n_138),
.D(n_153),
.Y(n_213)
);

OAI322xp33_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_229),
.A3(n_224),
.B1(n_214),
.B2(n_216),
.C1(n_215),
.C2(n_196),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_220),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_217),
.C(n_235),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_161),
.C(n_151),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_222),
.A2(n_224),
.B(n_230),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_0),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_225),
.A2(n_233),
.B1(n_197),
.B2(n_178),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

BUFx4f_ASAP7_75t_SL g229 ( 
.A(n_175),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_229),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_6),
.B(n_1),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_193),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_231),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_174),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_2),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_13),
.C(n_4),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_238),
.C(n_196),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_3),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_182),
.B(n_184),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_189),
.B(n_184),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_260),
.B(n_233),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_253),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_178),
.B(n_200),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_255),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_213),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_246),
.B(n_212),
.Y(n_272)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_247),
.Y(n_281)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

OAI321xp33_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_203),
.A3(n_198),
.B1(n_183),
.B2(n_199),
.C(n_187),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_232),
.B(n_239),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_210),
.C(n_187),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_259),
.C(n_238),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_174),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_177),
.C(n_205),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_222),
.A2(n_177),
.B(n_5),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_172),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_262),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_230),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_278),
.C(n_242),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_280),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_241),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_279),
.B(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_235),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_277),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_225),
.B1(n_220),
.B2(n_219),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_247),
.B1(n_241),
.B2(n_259),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_226),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_221),
.C(n_224),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_254),
.A2(n_236),
.B1(n_180),
.B2(n_6),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_251),
.B(n_4),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_269),
.B(n_261),
.Y(n_284)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_273),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_243),
.B(n_259),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_244),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_296),
.B1(n_275),
.B2(n_271),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_295),
.C(n_240),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_257),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_293),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_294),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_270),
.B(n_244),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_269),
.B(n_256),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_240),
.C(n_252),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_264),
.A2(n_243),
.B1(n_255),
.B2(n_250),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_298),
.B(n_299),
.Y(n_312)
);

AOI21x1_ASAP7_75t_SL g299 ( 
.A1(n_290),
.A2(n_243),
.B(n_263),
.Y(n_299)
);

NAND4xp25_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_267),
.C(n_249),
.D(n_248),
.Y(n_300)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_295),
.C(n_282),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_307),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_281),
.B1(n_274),
.B2(n_251),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_281),
.B1(n_279),
.B2(n_252),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_267),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_274),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_283),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_310),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_304),
.B(n_287),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_314),
.C(n_315),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_282),
.C(n_278),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_301),
.C(n_293),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_322),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_301),
.C(n_242),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_299),
.C(n_288),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_323),
.B(n_324),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_311),
.B(n_297),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_310),
.A2(n_285),
.B1(n_258),
.B2(n_305),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_325),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_312),
.B(n_316),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_319),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_331),
.B(n_327),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_329),
.Y(n_331)
);

AOI321xp33_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_328),
.A3(n_312),
.B1(n_309),
.B2(n_314),
.C(n_318),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_262),
.B(n_248),
.Y(n_334)
);


endmodule