module fake_netlist_1_5356_n_15 (n_1, n_2, n_4, n_3, n_0, n_15);
input n_1;
input n_2;
input n_4;
input n_3;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_10;
wire n_8;
AND2x4_ASAP7_75t_L g5 ( .A(n_1), .B(n_3), .Y(n_5) );
AND2x4_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_3), .Y(n_7) );
OAI21x1_ASAP7_75t_SL g8 ( .A1(n_7), .A2(n_0), .B(n_1), .Y(n_8) );
AOI22xp33_ASAP7_75t_L g9 ( .A1(n_5), .A2(n_2), .B1(n_4), .B2(n_6), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_9), .B(n_6), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
INVx1_ASAP7_75t_SL g13 ( .A(n_12), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
XNOR2x1_ASAP7_75t_L g15 ( .A(n_14), .B(n_10), .Y(n_15) );
endmodule