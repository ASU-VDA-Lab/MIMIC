module fake_jpeg_20834_n_189 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_189);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_12),
.Y(n_36)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_22),
.Y(n_45)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_23),
.B1(n_21),
.B2(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_21),
.B1(n_23),
.B2(n_20),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_19),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_44),
.B1(n_27),
.B2(n_31),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_20),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_27),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_23),
.Y(n_42)
);

AOI32xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_27),
.A3(n_24),
.B1(n_30),
.B2(n_25),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_29),
.A2(n_19),
.B1(n_13),
.B2(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_50),
.Y(n_64)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_42),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_29),
.B1(n_24),
.B2(n_32),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_42),
.B1(n_43),
.B2(n_40),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_42),
.B(n_38),
.C(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_30),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_43),
.B1(n_37),
.B2(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_50),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_59),
.B(n_49),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_68),
.B1(n_76),
.B2(n_58),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_44),
.C(n_41),
.Y(n_67)
);

AOI31xp33_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_71),
.A3(n_56),
.B(n_55),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_43),
.B1(n_40),
.B2(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_31),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_18),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_28),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_70),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_86),
.B1(n_61),
.B2(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_79),
.Y(n_103)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_81),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_90),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_53),
.B1(n_57),
.B2(n_51),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_88),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_88),
.A2(n_65),
.B1(n_61),
.B2(n_71),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_93),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_75),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_86),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_75),
.B(n_64),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_87),
.B(n_79),
.Y(n_112)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_73),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_113),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_18),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_118),
.B(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_104),
.B(n_82),
.Y(n_113)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_76),
.B(n_82),
.Y(n_115)
);

AOI21x1_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_73),
.B(n_28),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_92),
.C(n_93),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_95),
.C(n_28),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_106),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_120),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_115),
.C(n_107),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_112),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_124),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_48),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_132),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_11),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_11),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_48),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_118),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_108),
.B1(n_109),
.B2(n_113),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_108),
.B1(n_120),
.B2(n_121),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_130),
.C(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_146),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_149),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_148),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_107),
.B1(n_114),
.B2(n_37),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_151),
.B(n_157),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_132),
.CI(n_133),
.CON(n_153),
.SN(n_153)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_144),
.A2(n_126),
.B1(n_134),
.B2(n_137),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_37),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_148),
.C(n_139),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_157),
.B(n_151),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_114),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_155),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_161),
.B(n_166),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_0),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_162),
.B(n_163),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_0),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_153),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_154),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_0),
.B(n_1),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_166),
.B(n_161),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_152),
.C(n_22),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_173),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_18),
.C(n_2),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_1),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_170),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_172),
.C(n_4),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_174),
.B(n_1),
.Y(n_180)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_172),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.C1(n_2),
.C2(n_9),
.Y(n_181)
);

OA21x2_ASAP7_75t_SL g186 ( 
.A1(n_181),
.A2(n_9),
.B(n_10),
.Y(n_186)
);

OAI21x1_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_184),
.B(n_8),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_3),
.C(n_6),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_186),
.B(n_183),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_9),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_10),
.Y(n_189)
);


endmodule