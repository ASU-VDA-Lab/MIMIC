module fake_jpeg_25764_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx12_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_20),
.Y(n_28)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_29),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_26),
.B(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_11),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_14),
.B1(n_9),
.B2(n_12),
.Y(n_30)
);

AO21x1_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_23),
.B(n_12),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_16),
.B1(n_9),
.B2(n_19),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_13),
.C(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

NAND2x1_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_21),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_2),
.B(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_27),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_25),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_22),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_41),
.B(n_42),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_49),
.B(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_51),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_22),
.B1(n_13),
.B2(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_5),
.Y(n_55)
);


endmodule