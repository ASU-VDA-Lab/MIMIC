module fake_ariane_607_n_188 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_188);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_188;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_178;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_28;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_26),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_8),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_31),
.B(n_0),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

NAND2x1_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_6),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_6),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_29),
.B(n_7),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_40),
.B(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_38),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_50),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

OAI221xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_46),
.B1(n_39),
.B2(n_50),
.C(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_37),
.B1(n_45),
.B2(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_31),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_37),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_56),
.B1(n_54),
.B2(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

OR2x6_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_39),
.B1(n_34),
.B2(n_35),
.Y(n_86)
);

OAI221xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_57),
.B1(n_58),
.B2(n_68),
.C(n_62),
.Y(n_87)
);

NAND2x1p5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_48),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_70),
.B1(n_64),
.B2(n_56),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_60),
.Y(n_99)
);

OA21x2_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_87),
.B(n_27),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_82),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

OR2x6_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_90),
.Y(n_108)
);

AND2x4_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_92),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_91),
.B1(n_89),
.B2(n_78),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_98),
.B(n_97),
.C(n_94),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_71),
.B1(n_88),
.B2(n_84),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_84),
.B1(n_111),
.B2(n_102),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_88),
.B1(n_84),
.B2(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

OR2x6_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_114),
.B(n_107),
.Y(n_130)
);

NOR2x1p5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_106),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_102),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_106),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_88),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_72),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_128),
.Y(n_138)
);

OAI221xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_123),
.B1(n_125),
.B2(n_124),
.C(n_73),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_128),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_135),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_78),
.B1(n_127),
.B2(n_128),
.Y(n_144)
);

NAND2x1_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_121),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_69),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_130),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_106),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_106),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_63),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_63),
.C(n_69),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_7),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_8),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_100),
.C(n_51),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_9),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

NAND5xp2_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_154),
.C(n_155),
.D(n_76),
.E(n_156),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_72),
.Y(n_165)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_51),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_161),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_100),
.B1(n_51),
.B2(n_86),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_86),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_10),
.Y(n_171)
);

AOI221xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_86),
.B1(n_73),
.B2(n_82),
.C(n_72),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_11),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_SL g174 ( 
.A1(n_159),
.A2(n_167),
.B(n_165),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_86),
.B(n_100),
.Y(n_175)
);

AND4x1_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_12),
.C(n_14),
.D(n_101),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_162),
.C(n_100),
.Y(n_177)
);

AOI211xp5_ASAP7_75t_SL g178 ( 
.A1(n_173),
.A2(n_162),
.B(n_14),
.C(n_12),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

NAND4xp75_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_100),
.C(n_107),
.D(n_98),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_174),
.B1(n_175),
.B2(n_169),
.Y(n_182)
);

OR5x1_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_172),
.C(n_100),
.D(n_82),
.E(n_18),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_100),
.B1(n_82),
.B2(n_97),
.Y(n_184)
);

OAI322xp33_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_178),
.A3(n_181),
.B1(n_180),
.B2(n_99),
.C1(n_44),
.C2(n_107),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_16),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_183),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_185),
.B1(n_105),
.B2(n_89),
.Y(n_188)
);


endmodule