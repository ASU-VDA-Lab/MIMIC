module fake_netlist_5_2401_n_2032 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2032);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2032;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2009;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_314;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_63),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_14),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_53),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_98),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_33),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_77),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_36),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_103),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_116),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_39),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_110),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_76),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_56),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_31),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_53),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_163),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_114),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_59),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_99),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_18),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_140),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_127),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_107),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_89),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_65),
.Y(n_220)
);

INVx4_ASAP7_75t_R g221 ( 
.A(n_18),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_27),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_142),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_112),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_8),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_46),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_52),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_11),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_75),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_187),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_94),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_130),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_82),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_38),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_21),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_86),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_56),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_81),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_8),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_109),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_23),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_73),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_128),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_96),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_156),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_172),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_102),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_126),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_117),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_27),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_79),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_50),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_88),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_178),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_22),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_32),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_135),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_141),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_14),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_164),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_175),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_121),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_123),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_51),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_69),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_2),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_165),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_49),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_16),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_168),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_35),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_66),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_6),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_158),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_185),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_84),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_28),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_183),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_40),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_177),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_145),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_60),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_108),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_16),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_12),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_36),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_166),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_139),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_111),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_115),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_153),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_46),
.Y(n_296)
);

BUFx2_ASAP7_75t_SL g297 ( 
.A(n_85),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_0),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_26),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_104),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_176),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_12),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_167),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_93),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_180),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_55),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_174),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_97),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_51),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_159),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_87),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_43),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_122),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_149),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_131),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_13),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_150),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_124),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_54),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_9),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_184),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_105),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_23),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_1),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_33),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_15),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_25),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_43),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_45),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_60),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_59),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_17),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_62),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_91),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_67),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_147),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_157),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_80),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_160),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_55),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_106),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_92),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_29),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_72),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_38),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_113),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_15),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_42),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_11),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_48),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_42),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_57),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_48),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_143),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_146),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_2),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_144),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_54),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_41),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_181),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_5),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_100),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_28),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_154),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_83),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_137),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_7),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_35),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_101),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_64),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_20),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_90),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_151),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_1),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_155),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_39),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_4),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_71),
.Y(n_378)
);

CKINVDCx12_ASAP7_75t_R g379 ( 
.A(n_5),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_190),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_136),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_30),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_74),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_47),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_13),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_288),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_230),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_288),
.Y(n_388)
);

BUFx5_ASAP7_75t_L g389 ( 
.A(n_199),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_214),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_288),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_288),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_242),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_288),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_233),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_210),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_301),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_288),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_288),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_379),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_353),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_194),
.B(n_0),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_288),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_348),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_236),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_244),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_346),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_246),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_348),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_348),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_261),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_348),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_247),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_348),
.Y(n_415)
);

INVxp33_ASAP7_75t_SL g416 ( 
.A(n_324),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_370),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_258),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_275),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_249),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_250),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_370),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_261),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_268),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_252),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_268),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_299),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_299),
.Y(n_429)
);

INVxp33_ASAP7_75t_SL g430 ( 
.A(n_198),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_261),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_255),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_370),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_285),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_384),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_384),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_384),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_384),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_274),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_257),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_345),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_345),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_384),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_285),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_286),
.Y(n_446)
);

INVxp33_ASAP7_75t_L g447 ( 
.A(n_195),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_286),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_326),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_326),
.Y(n_450)
);

INVxp33_ASAP7_75t_SL g451 ( 
.A(n_198),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_264),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_203),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_265),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_285),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_308),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_207),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_212),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_228),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_365),
.Y(n_460)
);

INVxp33_ASAP7_75t_SL g461 ( 
.A(n_200),
.Y(n_461)
);

INVxp33_ASAP7_75t_SL g462 ( 
.A(n_200),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_231),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_269),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_205),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_271),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_213),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_254),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_276),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_284),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_256),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_287),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_260),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_196),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_263),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_206),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_289),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_316),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_330),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_216),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_349),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_387),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_412),
.B(n_294),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_405),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_423),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_410),
.Y(n_488)
);

OR2x6_ASAP7_75t_L g489 ( 
.A(n_392),
.B(n_297),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_201),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_423),
.B(n_201),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_424),
.B(n_248),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_390),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_476),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_411),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_386),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_411),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_438),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_431),
.B(n_248),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_438),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_413),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_388),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_413),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_425),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_435),
.B(n_278),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_415),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_417),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_419),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_445),
.B(n_278),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_417),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_388),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_455),
.B(n_193),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_474),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_416),
.A2(n_302),
.B1(n_238),
.B2(n_327),
.Y(n_518)
);

XNOR2x2_ASAP7_75t_R g519 ( 
.A(n_403),
.B(n_3),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_391),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_391),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_394),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_420),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_393),
.A2(n_234),
.B(n_193),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_407),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_393),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_395),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_433),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_414),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_433),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_396),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_395),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_401),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_399),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_434),
.B(n_234),
.Y(n_535)
);

OA21x2_ASAP7_75t_L g536 ( 
.A1(n_399),
.A2(n_361),
.B(n_359),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_400),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_434),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_400),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_467),
.B(n_266),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_421),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_480),
.B(n_292),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_422),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_436),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_436),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_444),
.B(n_202),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_427),
.B(n_266),
.Y(n_547)
);

OA21x2_ASAP7_75t_L g548 ( 
.A1(n_404),
.A2(n_367),
.B(n_363),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_437),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_404),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_389),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_389),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_389),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_L g554 ( 
.A(n_389),
.B(n_356),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_437),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_439),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_389),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_426),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_432),
.Y(n_559)
);

OA21x2_ASAP7_75t_L g560 ( 
.A1(n_439),
.A2(n_295),
.B(n_291),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_516),
.A2(n_398),
.B1(n_397),
.B2(n_408),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_484),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_484),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_502),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_542),
.B(n_441),
.Y(n_565)
);

CKINVDCx6p67_ASAP7_75t_R g566 ( 
.A(n_496),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_484),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_502),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_L g569 ( 
.A1(n_542),
.A2(n_518),
.B1(n_489),
.B2(n_496),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_502),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_517),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_520),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_494),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_484),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_507),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_520),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_526),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_L g579 ( 
.A(n_483),
.B(n_452),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_526),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_482),
.B(n_454),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_526),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_522),
.B(n_464),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_527),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_527),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_527),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_532),
.Y(n_587)
);

AND3x2_ASAP7_75t_L g588 ( 
.A(n_511),
.B(n_343),
.C(n_340),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_507),
.B(n_466),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_484),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_484),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_532),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_532),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_537),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_525),
.B(n_469),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_518),
.A2(n_290),
.B1(n_331),
.B2(n_312),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_537),
.Y(n_597)
);

NOR2x1p5_ASAP7_75t_L g598 ( 
.A(n_529),
.B(n_206),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_537),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_485),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_485),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_507),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_504),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_486),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_504),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_541),
.B(n_470),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_507),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_504),
.Y(n_608)
);

INVxp33_ASAP7_75t_L g609 ( 
.A(n_517),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_504),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_543),
.B(n_472),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_484),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_504),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_521),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_483),
.B(n_430),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_486),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_558),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_507),
.B(n_389),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_512),
.B(n_389),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_488),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_492),
.B(n_451),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_488),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_521),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_484),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_512),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_498),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_490),
.B(n_362),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_493),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_493),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_521),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_490),
.B(n_428),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_497),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_490),
.B(n_429),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_497),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_512),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_516),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_492),
.B(n_461),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_499),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_512),
.B(n_516),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_498),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_521),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_521),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_499),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_516),
.A2(n_356),
.B1(n_462),
.B2(n_290),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_534),
.Y(n_645)
);

AND2x6_ASAP7_75t_L g646 ( 
.A(n_516),
.B(n_291),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_534),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_534),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_512),
.B(n_389),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_534),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_498),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_534),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_550),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_495),
.A2(n_333),
.B1(n_373),
.B2(n_383),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_503),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_494),
.Y(n_656)
);

INVxp33_ASAP7_75t_SL g657 ( 
.A(n_511),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_503),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_505),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_550),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_498),
.Y(n_661)
);

INVx8_ASAP7_75t_L g662 ( 
.A(n_489),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_559),
.B(n_251),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_505),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_508),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_508),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_509),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_501),
.B(n_389),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_501),
.B(n_447),
.Y(n_669)
);

BUFx6f_ASAP7_75t_SL g670 ( 
.A(n_489),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_559),
.B(n_251),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_540),
.B(n_197),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_489),
.B(n_295),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_509),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_510),
.Y(n_675)
);

AND3x2_ASAP7_75t_L g676 ( 
.A(n_559),
.B(n_351),
.C(n_311),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_540),
.B(n_225),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_531),
.Y(n_678)
);

BUFx6f_ASAP7_75t_SL g679 ( 
.A(n_489),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_498),
.Y(n_680)
);

NAND2xp33_ASAP7_75t_L g681 ( 
.A(n_540),
.B(n_362),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_536),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_498),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_510),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_498),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_533),
.B(n_442),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_513),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_495),
.B(n_251),
.Y(n_688)
);

AO21x2_ASAP7_75t_L g689 ( 
.A1(n_554),
.A2(n_219),
.B(n_218),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_533),
.B(n_406),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_SL g691 ( 
.A(n_546),
.B(n_208),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_550),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_489),
.A2(n_226),
.B1(n_222),
.B2(n_227),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_513),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_L g695 ( 
.A(n_546),
.B(n_362),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_515),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_531),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_506),
.B(n_202),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_515),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_550),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_498),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_523),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_523),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_528),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_489),
.B(n_443),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_506),
.B(n_311),
.Y(n_706)
);

XNOR2xp5_ASAP7_75t_L g707 ( 
.A(n_519),
.B(n_403),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_506),
.B(n_409),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_536),
.Y(n_709)
);

OR2x6_ASAP7_75t_L g710 ( 
.A(n_547),
.B(n_380),
.Y(n_710)
);

INVx5_ASAP7_75t_L g711 ( 
.A(n_514),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_550),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_528),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_713),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_713),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_575),
.B(n_554),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_600),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_600),
.Y(n_718)
);

NOR3xp33_ASAP7_75t_L g719 ( 
.A(n_569),
.B(n_547),
.C(n_253),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_669),
.B(n_547),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_575),
.B(n_536),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_602),
.B(n_536),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_571),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_564),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_602),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_607),
.B(n_536),
.Y(n_726)
);

OR2x6_ASAP7_75t_L g727 ( 
.A(n_571),
.B(n_453),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_607),
.B(n_536),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_636),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_625),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_625),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_601),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_682),
.A2(n_548),
.B1(n_560),
.B2(n_524),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_SL g734 ( 
.A(n_635),
.B(n_362),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_635),
.Y(n_735)
);

BUFx8_ASAP7_75t_L g736 ( 
.A(n_670),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_601),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_604),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_621),
.B(n_237),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_636),
.B(n_639),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_609),
.B(n_418),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_604),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_615),
.A2(n_565),
.B1(n_705),
.B2(n_637),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_616),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_693),
.A2(n_208),
.B1(n_352),
.B2(n_347),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_589),
.A2(n_440),
.B1(n_456),
.B2(n_460),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_668),
.B(n_548),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_616),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_682),
.A2(n_548),
.B1(n_560),
.B2(n_524),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_620),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_709),
.B(n_548),
.Y(n_751)
);

NOR2xp67_ASAP7_75t_L g752 ( 
.A(n_708),
.B(n_491),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_672),
.A2(n_380),
.B1(n_375),
.B2(n_279),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_620),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_622),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_636),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_566),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_618),
.B(n_514),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_709),
.B(n_548),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_677),
.B(n_548),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_646),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_619),
.B(n_514),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_603),
.B(n_514),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_L g764 ( 
.A(n_646),
.B(n_267),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_603),
.B(n_514),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_712),
.B(n_514),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_564),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_688),
.B(n_204),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_712),
.B(n_514),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_605),
.B(n_514),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_581),
.B(n_491),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_605),
.B(n_539),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_566),
.B(n_453),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_631),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_608),
.B(n_539),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_622),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_628),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_608),
.B(n_539),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_568),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_663),
.B(n_204),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_610),
.B(n_539),
.Y(n_781)
);

AO221x1_ASAP7_75t_L g782 ( 
.A1(n_562),
.A2(n_362),
.B1(n_337),
.B2(n_341),
.C(n_342),
.Y(n_782)
);

AO221x1_ASAP7_75t_L g783 ( 
.A1(n_562),
.A2(n_335),
.B1(n_355),
.B2(n_317),
.C(n_314),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_610),
.B(n_539),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_628),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_629),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_671),
.B(n_693),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_686),
.B(n_209),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_613),
.B(n_539),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_613),
.B(n_539),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_657),
.B(n_579),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_629),
.Y(n_792)
);

BUFx5_ASAP7_75t_L g793 ( 
.A(n_646),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_649),
.B(n_539),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_657),
.B(n_209),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_670),
.A2(n_318),
.B1(n_315),
.B2(n_321),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_R g797 ( 
.A(n_573),
.B(n_211),
.Y(n_797)
);

BUFx6f_ASAP7_75t_SL g798 ( 
.A(n_617),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_614),
.B(n_556),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_690),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_632),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_568),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_632),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_634),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_673),
.A2(n_262),
.B1(n_313),
.B2(n_310),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_678),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_634),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_638),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_638),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_614),
.B(n_267),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_646),
.A2(n_560),
.B1(n_524),
.B2(n_491),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_631),
.B(n_457),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_623),
.B(n_267),
.Y(n_813)
);

INVx8_ASAP7_75t_L g814 ( 
.A(n_662),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_643),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_623),
.B(n_556),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_630),
.B(n_556),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_643),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_561),
.B(n_241),
.C(n_239),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_583),
.B(n_211),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_662),
.B(n_673),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_595),
.B(n_217),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_630),
.B(n_556),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_655),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_641),
.B(n_267),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_574),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_681),
.A2(n_491),
.B(n_530),
.C(n_538),
.Y(n_827)
);

NOR2x1p5_ASAP7_75t_L g828 ( 
.A(n_573),
.B(n_215),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_641),
.B(n_491),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_655),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_642),
.B(n_535),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_697),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_658),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_633),
.B(n_617),
.Y(n_834)
);

O2A1O1Ixp5_ASAP7_75t_L g835 ( 
.A1(n_642),
.A2(n_535),
.B(n_530),
.C(n_538),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_645),
.B(n_267),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_645),
.B(n_535),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_606),
.B(n_217),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_647),
.B(n_267),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_647),
.A2(n_560),
.B(n_552),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_L g841 ( 
.A(n_644),
.B(n_245),
.C(n_243),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_648),
.B(n_535),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_611),
.B(n_280),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_648),
.B(n_535),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_633),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_650),
.B(n_551),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_658),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_691),
.B(n_280),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_650),
.B(n_551),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_698),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_659),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_646),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_652),
.B(n_551),
.Y(n_853)
);

CKINVDCx16_ASAP7_75t_R g854 ( 
.A(n_617),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_652),
.B(n_551),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_617),
.B(n_275),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_653),
.B(n_552),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_654),
.B(n_457),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_654),
.B(n_275),
.Y(n_859)
);

O2A1O1Ixp5_ASAP7_75t_L g860 ( 
.A1(n_653),
.A2(n_660),
.B(n_700),
.C(n_692),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_646),
.A2(n_560),
.B1(n_267),
.B2(n_224),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_659),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_646),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_660),
.B(n_552),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_598),
.B(n_350),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_692),
.B(n_552),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_700),
.B(n_553),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_627),
.B(n_553),
.Y(n_868)
);

AND2x6_ASAP7_75t_L g869 ( 
.A(n_562),
.B(n_223),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_598),
.B(n_350),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_664),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_664),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_689),
.B(n_553),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_689),
.B(n_553),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_665),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_689),
.B(n_557),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_673),
.A2(n_710),
.B1(n_679),
.B2(n_670),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_665),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_673),
.A2(n_560),
.B1(n_267),
.B2(n_366),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_666),
.B(n_557),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_666),
.B(n_557),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_676),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_667),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_667),
.B(n_232),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_674),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_674),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_743),
.B(n_662),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_739),
.B(n_710),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_714),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_739),
.B(n_710),
.Y(n_890)
);

NAND2xp33_ASAP7_75t_L g891 ( 
.A(n_814),
.B(n_662),
.Y(n_891)
);

AND2x6_ASAP7_75t_SL g892 ( 
.A(n_741),
.B(n_707),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_714),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_715),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_774),
.B(n_673),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_715),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_716),
.A2(n_680),
.B(n_612),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_720),
.B(n_710),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_717),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_788),
.B(n_710),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_723),
.B(n_806),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_814),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_787),
.A2(n_679),
.B1(n_662),
.B2(n_596),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_723),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_793),
.B(n_563),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_787),
.B(n_596),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_SL g907 ( 
.A(n_798),
.B(n_679),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_834),
.B(n_697),
.Y(n_908)
);

CKINVDCx8_ASAP7_75t_R g909 ( 
.A(n_854),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_717),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_718),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_845),
.B(n_812),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_718),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_727),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_788),
.B(n_725),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_730),
.B(n_675),
.Y(n_916)
);

AND2x6_ASAP7_75t_SL g917 ( 
.A(n_820),
.B(n_707),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_731),
.B(n_675),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_752),
.A2(n_760),
.B1(n_740),
.B2(n_791),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_736),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_732),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_773),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_732),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_727),
.B(n_856),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_812),
.B(n_706),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_727),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_753),
.A2(n_695),
.B(n_706),
.C(n_704),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_737),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_793),
.B(n_563),
.Y(n_929)
);

OR2x6_ASAP7_75t_L g930 ( 
.A(n_821),
.B(n_706),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_760),
.A2(n_706),
.B1(n_694),
.B2(n_704),
.Y(n_931)
);

AND2x6_ASAP7_75t_L g932 ( 
.A(n_761),
.B(n_563),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_793),
.B(n_756),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_736),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_798),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_832),
.B(n_656),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_SL g937 ( 
.A(n_757),
.B(n_656),
.Y(n_937)
);

NOR2x1p5_ASAP7_75t_L g938 ( 
.A(n_858),
.B(n_215),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_738),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_738),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_742),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_771),
.B(n_821),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_740),
.A2(n_791),
.B1(n_735),
.B2(n_719),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_742),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_776),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_793),
.B(n_567),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_776),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_797),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_785),
.Y(n_949)
);

NAND2xp33_ASAP7_75t_SL g950 ( 
.A(n_865),
.B(n_282),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_814),
.Y(n_951)
);

AND2x6_ASAP7_75t_SL g952 ( 
.A(n_820),
.B(n_458),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_800),
.B(n_588),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_785),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_729),
.B(n_684),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_850),
.B(n_684),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_792),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_729),
.B(n_687),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_793),
.B(n_567),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_797),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_792),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_745),
.A2(n_706),
.B1(n_687),
.B2(n_703),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_822),
.A2(n_696),
.B1(n_703),
.B2(n_702),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_756),
.B(n_694),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_807),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_821),
.Y(n_966)
);

INVx5_ASAP7_75t_L g967 ( 
.A(n_761),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_807),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_744),
.Y(n_969)
);

NOR2x2_ASAP7_75t_L g970 ( 
.A(n_745),
.B(n_859),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_808),
.Y(n_971)
);

O2A1O1Ixp5_ASAP7_75t_L g972 ( 
.A1(n_835),
.A2(n_696),
.B(n_702),
.C(n_699),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_808),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_873),
.A2(n_680),
.B(n_612),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_882),
.Y(n_975)
);

AND2x4_ASAP7_75t_SL g976 ( 
.A(n_756),
.B(n_350),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_783),
.A2(n_699),
.B1(n_585),
.B2(n_599),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_824),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_870),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_824),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_793),
.B(n_567),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_756),
.Y(n_982)
);

INVx5_ASAP7_75t_L g983 ( 
.A(n_761),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_828),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_795),
.B(n_822),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_746),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_830),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_830),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_795),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_869),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_838),
.A2(n_591),
.B1(n_661),
.B2(n_685),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_748),
.B(n_572),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_750),
.B(n_572),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_847),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_754),
.B(n_576),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_761),
.B(n_591),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_755),
.B(n_576),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_819),
.B(n_458),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_780),
.B(n_591),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_886),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_847),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_852),
.B(n_661),
.Y(n_1002)
);

NOR2x1_ASAP7_75t_L g1003 ( 
.A(n_838),
.B(n_661),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_751),
.A2(n_585),
.B1(n_582),
.B2(n_593),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_777),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_786),
.B(n_577),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_851),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_851),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_801),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_803),
.B(n_577),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_871),
.Y(n_1011)
);

INVx5_ASAP7_75t_L g1012 ( 
.A(n_852),
.Y(n_1012)
);

AND2x2_ASAP7_75t_SL g1013 ( 
.A(n_879),
.B(n_235),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_871),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_878),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_843),
.A2(n_685),
.B1(n_683),
.B2(n_580),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_878),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_804),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_809),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_815),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_759),
.A2(n_593),
.B1(n_599),
.B2(n_580),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_841),
.B(n_459),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_818),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_833),
.B(n_582),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_874),
.A2(n_680),
.B(n_612),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_862),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_843),
.B(n_459),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_863),
.B(n_463),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_852),
.B(n_683),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_863),
.B(n_852),
.Y(n_1030)
);

INVxp67_ASAP7_75t_SL g1031 ( 
.A(n_721),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_872),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_875),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_883),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_885),
.B(n_578),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_831),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_879),
.A2(n_240),
.B1(n_305),
.B2(n_304),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_724),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_837),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_876),
.A2(n_590),
.B(n_574),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_780),
.B(n_463),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_842),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_722),
.B(n_578),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_811),
.B(n_861),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_811),
.B(n_683),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_726),
.A2(n_303),
.B1(n_685),
.B2(n_584),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_728),
.B(n_584),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_877),
.B(n_468),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_767),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_SL g1050 ( 
.A(n_768),
.B(n_222),
.C(n_220),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_861),
.B(n_574),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_844),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_826),
.B(n_586),
.Y(n_1053)
);

AND2x6_ASAP7_75t_SL g1054 ( 
.A(n_768),
.B(n_468),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_829),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_869),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_796),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_747),
.B(n_574),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_733),
.B(n_574),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_884),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_SL g1061 ( 
.A1(n_848),
.A2(n_358),
.B1(n_377),
.B2(n_281),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_846),
.B(n_849),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_779),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_SL g1064 ( 
.A1(n_848),
.A2(n_805),
.B1(n_764),
.B2(n_782),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_869),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_884),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_799),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_853),
.B(n_586),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_802),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_869),
.A2(n_587),
.B1(n_592),
.B2(n_594),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_855),
.B(n_587),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_L g1072 ( 
.A(n_810),
.B(n_270),
.C(n_259),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_816),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_869),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_810),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_813),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_857),
.B(n_864),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_866),
.B(n_592),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_817),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_906),
.A2(n_1044),
.B1(n_1013),
.B2(n_903),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_985),
.B(n_880),
.Y(n_1081)
);

BUFx4f_ASAP7_75t_L g1082 ( 
.A(n_924),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_906),
.A2(n_827),
.B(n_860),
.C(n_823),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_982),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1044),
.A2(n_749),
.B(n_733),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_888),
.A2(n_839),
.B(n_825),
.C(n_836),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_889),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_989),
.A2(n_762),
.B1(n_758),
.B2(n_794),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_982),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_982),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_893),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_901),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_922),
.B(n_758),
.Y(n_1093)
);

AO32x1_ASAP7_75t_L g1094 ( 
.A1(n_1037),
.A2(n_479),
.A3(n_481),
.B1(n_478),
.B2(n_477),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1036),
.B(n_881),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_893),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1051),
.A2(n_749),
.B(n_762),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_890),
.A2(n_813),
.B(n_839),
.C(n_836),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_982),
.Y(n_1099)
);

NOR3xp33_ASAP7_75t_SL g1100 ( 
.A(n_1050),
.B(n_948),
.C(n_953),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_894),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1027),
.B(n_471),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1051),
.A2(n_794),
.B(n_868),
.Y(n_1103)
);

AO21x1_ASAP7_75t_L g1104 ( 
.A1(n_900),
.A2(n_825),
.B(n_765),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_904),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_986),
.B(n_867),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_899),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_899),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1062),
.A2(n_1077),
.B(n_1031),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_896),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1039),
.B(n_763),
.Y(n_1111)
);

O2A1O1Ixp5_ASAP7_75t_L g1112 ( 
.A1(n_887),
.A2(n_734),
.B(n_840),
.C(n_789),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_915),
.A2(n_898),
.B(n_979),
.C(n_1022),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_975),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_914),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_908),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_910),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1013),
.A2(n_790),
.B1(n_784),
.B2(n_781),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_911),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_L g1120 ( 
.A(n_1061),
.B(n_273),
.C(n_272),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1031),
.A2(n_769),
.B(n_766),
.Y(n_1121)
);

OAI22x1_ASAP7_75t_L g1122 ( 
.A1(n_938),
.A2(n_352),
.B1(n_226),
.B2(n_227),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_902),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_913),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_L g1125 ( 
.A(n_936),
.B(n_293),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_909),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1041),
.B(n_471),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_921),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_910),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1042),
.B(n_770),
.Y(n_1130)
);

OAI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1057),
.A2(n_368),
.B1(n_229),
.B2(n_281),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_960),
.B(n_952),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_974),
.A2(n_778),
.B(n_775),
.Y(n_1133)
);

BUFx12f_ASAP7_75t_L g1134 ( 
.A(n_935),
.Y(n_1134)
);

OAI22x1_ASAP7_75t_L g1135 ( 
.A1(n_926),
.A2(n_220),
.B1(n_229),
.B2(n_347),
.Y(n_1135)
);

INVxp67_ASAP7_75t_SL g1136 ( 
.A(n_1030),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_912),
.B(n_282),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_953),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_887),
.A2(n_300),
.B1(n_307),
.B2(n_322),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_1030),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_962),
.A2(n_919),
.B1(n_1052),
.B2(n_943),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_902),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1025),
.A2(n_1059),
.B(n_1045),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_912),
.B(n_772),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1055),
.B(n_594),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_925),
.A2(n_381),
.B1(n_378),
.B2(n_372),
.Y(n_1146)
);

BUFx5_ASAP7_75t_L g1147 ( 
.A(n_932),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_967),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_923),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_937),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_923),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_925),
.B(n_956),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_895),
.B(n_344),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_962),
.A2(n_374),
.B1(n_358),
.B2(n_368),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_920),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1055),
.B(n_1067),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_966),
.B(n_942),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1028),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1059),
.A2(n_701),
.B(n_651),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_928),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_895),
.A2(n_339),
.B1(n_338),
.B2(n_336),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_998),
.A2(n_481),
.B(n_475),
.C(n_477),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1060),
.A2(n_999),
.B(n_927),
.C(n_1076),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1054),
.B(n_277),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1045),
.A2(n_1040),
.B(n_891),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_933),
.A2(n_701),
.B(n_651),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1048),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1073),
.B(n_597),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_SL g1169 ( 
.A(n_990),
.B(n_344),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_969),
.A2(n_479),
.B(n_478),
.C(n_475),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_907),
.B(n_354),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1066),
.B(n_283),
.Y(n_1172)
);

AO22x1_ASAP7_75t_L g1173 ( 
.A1(n_966),
.A2(n_371),
.B1(n_382),
.B2(n_377),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_939),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_967),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_940),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_999),
.A2(n_1028),
.B(n_1072),
.C(n_950),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_933),
.A2(n_897),
.B(n_1043),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1009),
.B(n_296),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1047),
.A2(n_701),
.B(n_651),
.Y(n_1180)
);

INVx4_ASAP7_75t_L g1181 ( 
.A(n_902),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_969),
.A2(n_473),
.B(n_597),
.C(n_545),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1058),
.A2(n_626),
.B(n_701),
.Y(n_1183)
);

NOR3xp33_ASAP7_75t_SL g1184 ( 
.A(n_970),
.B(n_371),
.C(n_382),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_892),
.B(n_354),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_944),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_967),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_902),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_928),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1079),
.B(n_570),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_976),
.B(n_473),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1079),
.B(n_941),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1064),
.A2(n_376),
.B1(n_374),
.B2(n_332),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_963),
.A2(n_369),
.B(n_357),
.C(n_360),
.Y(n_1194)
);

AO21x2_ASAP7_75t_L g1195 ( 
.A1(n_931),
.A2(n_549),
.B(n_544),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1058),
.A2(n_626),
.B(n_701),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1018),
.B(n_357),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_941),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_945),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_917),
.B(n_298),
.Y(n_1200)
);

O2A1O1Ixp5_ASAP7_75t_SL g1201 ( 
.A1(n_1019),
.A2(n_446),
.B(n_448),
.C(n_449),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1005),
.A2(n_549),
.B(n_545),
.C(n_544),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_954),
.B(n_957),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_984),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_964),
.A2(n_651),
.B(n_590),
.Y(n_1205)
);

AOI33xp33_ASAP7_75t_L g1206 ( 
.A1(n_977),
.A2(n_450),
.A3(n_449),
.B1(n_448),
.B2(n_446),
.B3(n_376),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_967),
.B(n_364),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1004),
.A2(n_323),
.B1(n_328),
.B2(n_306),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_976),
.B(n_450),
.Y(n_1209)
);

OAI21xp33_ASAP7_75t_SL g1210 ( 
.A1(n_1070),
.A2(n_570),
.B(n_221),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1005),
.B(n_309),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_972),
.A2(n_557),
.B(n_711),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_954),
.B(n_590),
.Y(n_1213)
);

AND2x2_ASAP7_75t_SL g1214 ( 
.A(n_951),
.B(n_590),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1053),
.A2(n_651),
.B(n_626),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_955),
.A2(n_626),
.B(n_590),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1000),
.B(n_319),
.Y(n_1217)
);

NAND2x1p5_ASAP7_75t_L g1218 ( 
.A(n_951),
.B(n_626),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_958),
.A2(n_711),
.B(n_640),
.Y(n_1219)
);

BUFx10_ASAP7_75t_L g1220 ( 
.A(n_1048),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1000),
.B(n_320),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1075),
.A2(n_334),
.B1(n_381),
.B2(n_364),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_957),
.B(n_487),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1048),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_983),
.B(n_369),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_961),
.B(n_487),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_947),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_961),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_905),
.A2(n_711),
.B(n_640),
.Y(n_1229)
);

O2A1O1Ixp5_ASAP7_75t_SL g1230 ( 
.A1(n_1020),
.A2(n_500),
.B(n_487),
.C(n_385),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_965),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_949),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_968),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_905),
.A2(n_711),
.B(n_640),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_951),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1026),
.Y(n_1236)
);

NOR3xp33_ASAP7_75t_L g1237 ( 
.A(n_916),
.B(n_325),
.C(n_378),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1034),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_929),
.A2(n_711),
.B(n_640),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_929),
.A2(n_711),
.B(n_640),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1023),
.B(n_372),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_973),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_951),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1023),
.B(n_1032),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1140),
.Y(n_1245)
);

NOR2x1_ASAP7_75t_L g1246 ( 
.A(n_1181),
.B(n_920),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1092),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1109),
.A2(n_1065),
.B(n_1012),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1244),
.Y(n_1249)
);

AO21x1_ASAP7_75t_L g1250 ( 
.A1(n_1080),
.A2(n_1141),
.B(n_1113),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1114),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1159),
.A2(n_1196),
.B(n_1183),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1102),
.B(n_918),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1115),
.Y(n_1254)
);

AOI221xp5_ASAP7_75t_L g1255 ( 
.A1(n_1131),
.A2(n_977),
.B1(n_934),
.B2(n_1046),
.C(n_1033),
.Y(n_1255)
);

INVxp67_ASAP7_75t_SL g1256 ( 
.A(n_1136),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1165),
.A2(n_1065),
.B(n_1012),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1133),
.A2(n_1035),
.B(n_1024),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1080),
.A2(n_1003),
.B(n_1016),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1178),
.A2(n_1065),
.B(n_1012),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1163),
.A2(n_1065),
.B(n_1012),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1143),
.A2(n_992),
.B(n_1006),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1123),
.Y(n_1263)
);

OAI21xp33_ASAP7_75t_SL g1264 ( 
.A1(n_1141),
.A2(n_1070),
.B(n_1004),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1123),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1087),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1085),
.A2(n_983),
.B(n_1071),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1127),
.B(n_1032),
.Y(n_1268)
);

NAND3x1_ASAP7_75t_L g1269 ( 
.A(n_1132),
.B(n_934),
.C(n_1038),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1116),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1101),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1156),
.B(n_1033),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1121),
.A2(n_1103),
.B(n_1095),
.Y(n_1273)
);

CKINVDCx14_ASAP7_75t_R g1274 ( 
.A(n_1126),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1155),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1104),
.A2(n_991),
.B(n_946),
.Y(n_1276)
);

AOI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1097),
.A2(n_1010),
.B(n_997),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1166),
.A2(n_995),
.B(n_993),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1105),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1212),
.A2(n_965),
.B(n_980),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1156),
.B(n_980),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1212),
.A2(n_1180),
.B(n_1215),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1205),
.A2(n_988),
.B(n_1007),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1095),
.A2(n_983),
.B(n_1078),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1081),
.B(n_988),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_1123),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1083),
.A2(n_1007),
.A3(n_1068),
.B(n_1014),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1086),
.A2(n_983),
.B(n_981),
.Y(n_1288)
);

OAI21xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1206),
.A2(n_1021),
.B(n_946),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1118),
.A2(n_1008),
.A3(n_987),
.B(n_994),
.Y(n_1290)
);

INVxp67_ASAP7_75t_SL g1291 ( 
.A(n_1140),
.Y(n_1291)
);

CKINVDCx8_ASAP7_75t_R g1292 ( 
.A(n_1157),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1081),
.B(n_978),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1106),
.A2(n_930),
.B1(n_1017),
.B2(n_1011),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1110),
.Y(n_1295)
);

BUFx4f_ASAP7_75t_L g1296 ( 
.A(n_1134),
.Y(n_1296)
);

CKINVDCx11_ASAP7_75t_R g1297 ( 
.A(n_1220),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1142),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1177),
.A2(n_1074),
.B(n_1001),
.C(n_1038),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1093),
.A2(n_1074),
.B(n_1069),
.C(n_1063),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1144),
.B(n_971),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1118),
.A2(n_1015),
.A3(n_1063),
.B(n_1069),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1098),
.A2(n_959),
.B(n_981),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1192),
.B(n_1049),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1210),
.A2(n_1021),
.B(n_996),
.Y(n_1305)
);

AO32x2_ASAP7_75t_L g1306 ( 
.A1(n_1193),
.A2(n_930),
.A3(n_1049),
.B1(n_1029),
.B2(n_1002),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1216),
.A2(n_959),
.B(n_1029),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1112),
.A2(n_1002),
.B(n_996),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_SL g1309 ( 
.A1(n_1194),
.A2(n_930),
.B(n_932),
.C(n_1056),
.Y(n_1309)
);

AOI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1219),
.A2(n_932),
.B(n_1056),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1111),
.A2(n_1056),
.B(n_640),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1191),
.B(n_1056),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1119),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1237),
.A2(n_500),
.B(n_487),
.C(n_932),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1138),
.A2(n_932),
.B1(n_500),
.B2(n_487),
.Y(n_1315)
);

AO22x2_ASAP7_75t_L g1316 ( 
.A1(n_1193),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1236),
.A2(n_624),
.B1(n_500),
.B2(n_555),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1217),
.Y(n_1318)
);

OAI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1150),
.A2(n_624),
.B1(n_555),
.B2(n_500),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1111),
.A2(n_624),
.B(n_555),
.Y(n_1320)
);

AO32x2_ASAP7_75t_L g1321 ( 
.A1(n_1154),
.A2(n_9),
.A3(n_10),
.B1(n_17),
.B2(n_19),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1221),
.A2(n_555),
.B(n_624),
.C(n_20),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1130),
.A2(n_624),
.B(n_555),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1192),
.B(n_10),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1236),
.B(n_19),
.Y(n_1325)
);

NAND2x1p5_ASAP7_75t_L g1326 ( 
.A(n_1181),
.B(n_624),
.Y(n_1326)
);

NOR3xp33_ASAP7_75t_SL g1327 ( 
.A(n_1200),
.B(n_1164),
.C(n_1120),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1124),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1238),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1172),
.B(n_21),
.Y(n_1330)
);

NAND3x1_ASAP7_75t_L g1331 ( 
.A(n_1222),
.B(n_22),
.C(n_24),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1128),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1229),
.A2(n_555),
.B(n_192),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1088),
.A2(n_133),
.B(n_189),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1130),
.A2(n_555),
.B(n_188),
.Y(n_1335)
);

NOR2xp67_ASAP7_75t_L g1336 ( 
.A(n_1188),
.B(n_186),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1152),
.A2(n_555),
.B(n_173),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1238),
.B(n_24),
.Y(n_1338)
);

INVx4_ASAP7_75t_L g1339 ( 
.A(n_1142),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1142),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1224),
.B(n_170),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1168),
.A2(n_169),
.B(n_161),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1168),
.A2(n_152),
.B(n_148),
.Y(n_1343)
);

AO31x2_ASAP7_75t_L g1344 ( 
.A1(n_1230),
.A2(n_25),
.A3(n_26),
.B(n_29),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1241),
.B(n_30),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1184),
.A2(n_31),
.B(n_32),
.C(n_34),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1214),
.A2(n_134),
.B(n_132),
.Y(n_1347)
);

AOI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1145),
.A2(n_1190),
.B(n_1226),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1082),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1209),
.B(n_37),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1082),
.A2(n_1158),
.B1(n_1242),
.B2(n_1199),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1145),
.A2(n_129),
.B(n_125),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1203),
.A2(n_120),
.B(n_119),
.Y(n_1353)
);

BUFx12f_ASAP7_75t_L g1354 ( 
.A(n_1220),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1211),
.B(n_41),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1167),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_1356)
);

A2O1A1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1179),
.A2(n_44),
.B(n_49),
.C(n_50),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1157),
.B(n_1100),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1174),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1139),
.A2(n_52),
.B(n_57),
.C(n_58),
.Y(n_1360)
);

INVxp67_ASAP7_75t_SL g1361 ( 
.A(n_1084),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1235),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1203),
.A2(n_118),
.B(n_95),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1190),
.B(n_58),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1204),
.B(n_78),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1135),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1234),
.A2(n_68),
.B(n_70),
.Y(n_1367)
);

AO21x2_ASAP7_75t_L g1368 ( 
.A1(n_1195),
.A2(n_61),
.B(n_62),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1091),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1176),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1188),
.B(n_61),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1195),
.A2(n_63),
.B(n_64),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1208),
.B(n_65),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1096),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1208),
.B(n_1232),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1239),
.A2(n_1240),
.B(n_1213),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_1122),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1084),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1182),
.A2(n_1125),
.B(n_1161),
.C(n_1170),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1213),
.A2(n_1227),
.A3(n_1233),
.B(n_1186),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1223),
.A2(n_1226),
.B(n_1201),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1148),
.A2(n_1187),
.B(n_1175),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1223),
.A2(n_1225),
.B(n_1207),
.Y(n_1383)
);

AOI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1107),
.A2(n_1160),
.B(n_1189),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1185),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1148),
.A2(n_1187),
.B(n_1175),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1154),
.B(n_1146),
.Y(n_1387)
);

A2O1A1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1202),
.A2(n_1162),
.B(n_1153),
.C(n_1197),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1243),
.B(n_1099),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1218),
.A2(n_1094),
.B(n_1198),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1218),
.A2(n_1117),
.B(n_1151),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1169),
.B(n_1171),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1173),
.B(n_1169),
.C(n_1137),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1108),
.B(n_1129),
.C(n_1231),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1149),
.A2(n_1228),
.B(n_1089),
.C(n_1090),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1089),
.B(n_1090),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1147),
.A2(n_1094),
.B(n_1099),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1243),
.A2(n_1147),
.B1(n_1084),
.B2(n_1094),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1147),
.A2(n_739),
.B(n_985),
.C(n_906),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1243),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1147),
.A2(n_1159),
.B(n_1183),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1147),
.A2(n_1159),
.B(n_1183),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1102),
.B(n_985),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1114),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1244),
.Y(n_1405)
);

AO21x1_ASAP7_75t_L g1406 ( 
.A1(n_1080),
.A2(n_1141),
.B(n_900),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1092),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1080),
.A2(n_739),
.B(n_743),
.C(n_985),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1109),
.A2(n_1044),
.B(n_1165),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1159),
.A2(n_1196),
.B(n_1183),
.Y(n_1410)
);

NAND3xp33_ASAP7_75t_L g1411 ( 
.A(n_1080),
.B(n_739),
.C(n_743),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1109),
.A2(n_1044),
.B(n_1165),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1403),
.B(n_1253),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1266),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1411),
.A2(n_1408),
.B(n_1399),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1271),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_SL g1417 ( 
.A(n_1411),
.B(n_1393),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1268),
.B(n_1272),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1245),
.B(n_1312),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1350),
.B(n_1318),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1358),
.B(n_1249),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1405),
.B(n_1329),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1330),
.B(n_1327),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1259),
.A2(n_1412),
.B(n_1409),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1257),
.A2(n_1376),
.B(n_1333),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_SL g1426 ( 
.A1(n_1372),
.A2(n_1383),
.B(n_1334),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1252),
.A2(n_1410),
.B(n_1283),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1273),
.A2(n_1390),
.B(n_1305),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1302),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1282),
.A2(n_1258),
.B(n_1262),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1281),
.B(n_1387),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1295),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1267),
.A2(n_1307),
.B(n_1278),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1355),
.B(n_1407),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1316),
.A2(n_1373),
.B1(n_1406),
.B2(n_1250),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1313),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1302),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1324),
.B(n_1247),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1356),
.A2(n_1393),
.B1(n_1366),
.B2(n_1377),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1351),
.B(n_1261),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1301),
.B(n_1293),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1302),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1275),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1379),
.A2(n_1388),
.B(n_1299),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1328),
.Y(n_1445)
);

BUFx8_ASAP7_75t_L g1446 ( 
.A(n_1254),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1248),
.A2(n_1280),
.B(n_1310),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1332),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_SL g1449 ( 
.A1(n_1360),
.A2(n_1357),
.B(n_1322),
.C(n_1314),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1346),
.B(n_1356),
.C(n_1349),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1274),
.Y(n_1451)
);

AO31x2_ASAP7_75t_L g1452 ( 
.A1(n_1300),
.A2(n_1303),
.A3(n_1288),
.B(n_1395),
.Y(n_1452)
);

NAND3xp33_ASAP7_75t_SL g1453 ( 
.A(n_1345),
.B(n_1392),
.C(n_1255),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1375),
.B(n_1270),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1287),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1359),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1245),
.B(n_1396),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1370),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1389),
.B(n_1369),
.Y(n_1459)
);

AOI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1316),
.A2(n_1264),
.B1(n_1338),
.B2(n_1325),
.C(n_1289),
.Y(n_1460)
);

NOR2xp67_ASAP7_75t_L g1461 ( 
.A(n_1251),
.B(n_1404),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1289),
.A2(n_1294),
.B(n_1284),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1374),
.Y(n_1463)
);

CKINVDCx14_ASAP7_75t_R g1464 ( 
.A(n_1296),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1264),
.A2(n_1352),
.B1(n_1364),
.B2(n_1368),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1397),
.A2(n_1308),
.B(n_1277),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1389),
.B(n_1291),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1367),
.A2(n_1381),
.B(n_1348),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1380),
.Y(n_1469)
);

INVx8_ASAP7_75t_L g1470 ( 
.A(n_1263),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1294),
.A2(n_1347),
.B(n_1335),
.C(n_1342),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1309),
.A2(n_1279),
.B(n_1341),
.C(n_1365),
.Y(n_1472)
);

NAND2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1246),
.B(n_1339),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1304),
.B(n_1256),
.Y(n_1474)
);

AO21x2_ASAP7_75t_L g1475 ( 
.A1(n_1398),
.A2(n_1276),
.B(n_1311),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1341),
.A2(n_1285),
.B1(n_1292),
.B2(n_1354),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1400),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1380),
.Y(n_1478)
);

AO31x2_ASAP7_75t_L g1479 ( 
.A1(n_1317),
.A2(n_1323),
.A3(n_1320),
.B(n_1306),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1341),
.A2(n_1365),
.B(n_1371),
.C(n_1343),
.Y(n_1480)
);

AO31x2_ASAP7_75t_L g1481 ( 
.A1(n_1306),
.A2(n_1344),
.A3(n_1363),
.B(n_1353),
.Y(n_1481)
);

BUFx8_ASAP7_75t_L g1482 ( 
.A(n_1263),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1287),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1398),
.A2(n_1394),
.B(n_1391),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1337),
.A2(n_1386),
.B(n_1382),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1297),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1368),
.A2(n_1319),
.B(n_1331),
.C(n_1276),
.Y(n_1487)
);

INVx4_ASAP7_75t_SL g1488 ( 
.A(n_1263),
.Y(n_1488)
);

OAI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1394),
.A2(n_1315),
.B(n_1336),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1315),
.A2(n_1336),
.B(n_1290),
.Y(n_1490)
);

OA21x2_ASAP7_75t_L g1491 ( 
.A1(n_1306),
.A2(n_1290),
.B(n_1344),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1361),
.A2(n_1326),
.B(n_1378),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1269),
.A2(n_1287),
.B(n_1290),
.Y(n_1493)
);

AO31x2_ASAP7_75t_L g1494 ( 
.A1(n_1344),
.A2(n_1321),
.A3(n_1286),
.B(n_1339),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1378),
.A2(n_1265),
.B(n_1286),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1298),
.Y(n_1496)
);

A2O1A1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1321),
.A2(n_1296),
.B(n_1298),
.C(n_1340),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1298),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1265),
.A2(n_1340),
.B(n_1362),
.Y(n_1499)
);

OA21x2_ASAP7_75t_L g1500 ( 
.A1(n_1321),
.A2(n_1385),
.B(n_1340),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1362),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1362),
.A2(n_1260),
.B(n_1401),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1409),
.A2(n_1412),
.B(n_1259),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1411),
.A2(n_739),
.B(n_743),
.Y(n_1504)
);

AOI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1260),
.A2(n_1267),
.B(n_1165),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1411),
.A2(n_1408),
.B(n_906),
.C(n_1264),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1411),
.A2(n_739),
.B(n_743),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1409),
.A2(n_1412),
.B(n_1259),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1275),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1260),
.A2(n_1402),
.B(n_1401),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1350),
.B(n_908),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1403),
.B(n_1407),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1411),
.A2(n_739),
.B(n_743),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1245),
.B(n_1157),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1350),
.B(n_908),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1411),
.A2(n_906),
.B1(n_739),
.B2(n_1408),
.C(n_745),
.Y(n_1516)
);

NAND3xp33_ASAP7_75t_L g1517 ( 
.A(n_1411),
.B(n_739),
.C(n_743),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1409),
.A2(n_1412),
.B(n_1259),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1266),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1409),
.A2(n_1412),
.B(n_1259),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1275),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1403),
.B(n_985),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1273),
.A2(n_1109),
.B(n_1409),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1403),
.B(n_1407),
.Y(n_1524)
);

AO21x2_ASAP7_75t_L g1525 ( 
.A1(n_1259),
.A2(n_1412),
.B(n_1409),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1329),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1260),
.A2(n_1402),
.B(n_1401),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1263),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1266),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1411),
.B(n_739),
.Y(n_1530)
);

AOI21xp33_ASAP7_75t_L g1531 ( 
.A1(n_1411),
.A2(n_739),
.B(n_985),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1260),
.A2(n_1402),
.B(n_1401),
.Y(n_1532)
);

NAND2x1p5_ASAP7_75t_L g1533 ( 
.A(n_1245),
.B(n_982),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1403),
.B(n_985),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1411),
.A2(n_739),
.B(n_743),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1259),
.A2(n_1412),
.B(n_1409),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1409),
.A2(n_1412),
.B(n_1259),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1260),
.A2(n_1402),
.B(n_1401),
.Y(n_1538)
);

AOI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1260),
.A2(n_1267),
.B(n_1165),
.Y(n_1539)
);

AO32x2_ASAP7_75t_L g1540 ( 
.A1(n_1349),
.A2(n_1080),
.A3(n_1141),
.B1(n_1193),
.B2(n_1351),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1409),
.A2(n_1412),
.B(n_1259),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1403),
.B(n_985),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1384),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1329),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_SL g1545 ( 
.A(n_1296),
.B(n_697),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_SL g1546 ( 
.A1(n_1316),
.A2(n_906),
.B1(n_1411),
.B2(n_1080),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1260),
.A2(n_1402),
.B(n_1401),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1245),
.B(n_1157),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1403),
.B(n_1407),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1245),
.B(n_1157),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1260),
.A2(n_1402),
.B(n_1401),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1245),
.B(n_1157),
.Y(n_1552)
);

O2A1O1Ixp5_ASAP7_75t_L g1553 ( 
.A1(n_1250),
.A2(n_1411),
.B(n_1408),
.C(n_1406),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1274),
.Y(n_1554)
);

A2O1A1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1411),
.A2(n_1408),
.B(n_906),
.C(n_1264),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1389),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1351),
.B(n_1399),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1259),
.A2(n_1412),
.B(n_1409),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1350),
.B(n_908),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1329),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1260),
.A2(n_1402),
.B(n_1401),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1411),
.A2(n_906),
.B1(n_985),
.B2(n_1330),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1247),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1329),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1411),
.A2(n_739),
.B(n_743),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1411),
.A2(n_906),
.B1(n_985),
.B2(n_1330),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_SL g1567 ( 
.A(n_1296),
.B(n_697),
.Y(n_1567)
);

AOI221xp5_ASAP7_75t_L g1568 ( 
.A1(n_1411),
.A2(n_906),
.B1(n_739),
.B2(n_1408),
.C(n_745),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1415),
.B(n_1500),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1526),
.Y(n_1570)
);

OA22x2_ASAP7_75t_L g1571 ( 
.A1(n_1439),
.A2(n_1513),
.B1(n_1565),
.B2(n_1504),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1478),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1526),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1562),
.A2(n_1566),
.B1(n_1530),
.B2(n_1450),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1544),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1562),
.A2(n_1566),
.B1(n_1530),
.B2(n_1546),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1462),
.A2(n_1523),
.B(n_1468),
.Y(n_1577)
);

BUFx2_ASAP7_75t_SL g1578 ( 
.A(n_1461),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1413),
.B(n_1441),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1522),
.B(n_1534),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1531),
.A2(n_1507),
.B(n_1535),
.C(n_1453),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1421),
.B(n_1420),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1542),
.B(n_1418),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1512),
.B(n_1524),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1516),
.A2(n_1568),
.B(n_1444),
.C(n_1517),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1500),
.B(n_1546),
.Y(n_1586)
);

O2A1O1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1423),
.A2(n_1506),
.B(n_1555),
.C(n_1471),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1549),
.B(n_1454),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1431),
.B(n_1434),
.Y(n_1589)
);

BUFx12f_ASAP7_75t_L g1590 ( 
.A(n_1486),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1435),
.A2(n_1555),
.B1(n_1506),
.B2(n_1476),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1435),
.A2(n_1476),
.B1(n_1438),
.B2(n_1434),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1509),
.Y(n_1593)
);

BUFx4f_ASAP7_75t_SL g1594 ( 
.A(n_1486),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1422),
.B(n_1417),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1544),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1500),
.B(n_1497),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1497),
.B(n_1540),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1540),
.B(n_1455),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1560),
.B(n_1564),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1424),
.A2(n_1525),
.B(n_1558),
.Y(n_1601)
);

BUFx12f_ASAP7_75t_L g1602 ( 
.A(n_1451),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1540),
.B(n_1455),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1560),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1564),
.B(n_1474),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1451),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1554),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1465),
.A2(n_1557),
.B1(n_1460),
.B2(n_1511),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1424),
.A2(n_1525),
.B(n_1558),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1419),
.B(n_1457),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1528),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1414),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1416),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1540),
.B(n_1483),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1515),
.B(n_1559),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1419),
.B(n_1457),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1419),
.B(n_1457),
.Y(n_1617)
);

OA21x2_ASAP7_75t_L g1618 ( 
.A1(n_1466),
.A2(n_1553),
.B(n_1433),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1432),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1480),
.A2(n_1471),
.B(n_1472),
.Y(n_1620)
);

O2A1O1Ixp33_ASAP7_75t_L g1621 ( 
.A1(n_1449),
.A2(n_1426),
.B(n_1553),
.C(n_1557),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1463),
.B(n_1459),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1493),
.B(n_1469),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1459),
.B(n_1467),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1436),
.B(n_1445),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1448),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1465),
.A2(n_1557),
.B1(n_1464),
.B2(n_1563),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1467),
.B(n_1556),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1514),
.B(n_1548),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1548),
.B(n_1550),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1491),
.B(n_1456),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1458),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1536),
.A2(n_1518),
.B(n_1508),
.Y(n_1633)
);

OA21x2_ASAP7_75t_L g1634 ( 
.A1(n_1466),
.A2(n_1427),
.B(n_1430),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1489),
.A2(n_1487),
.B(n_1440),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1477),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1554),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1519),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1440),
.A2(n_1518),
.B(n_1537),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1552),
.B(n_1529),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1543),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1556),
.B(n_1552),
.Y(n_1642)
);

O2A1O1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1449),
.A2(n_1440),
.B(n_1567),
.C(n_1545),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1495),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1503),
.A2(n_1508),
.B(n_1541),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1494),
.B(n_1498),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1429),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1498),
.B(n_1501),
.Y(n_1648)
);

NOR2xp67_ASAP7_75t_L g1649 ( 
.A(n_1443),
.B(n_1499),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1509),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_SL g1651 ( 
.A1(n_1508),
.A2(n_1537),
.B(n_1520),
.Y(n_1651)
);

O2A1O1Ixp5_ASAP7_75t_L g1652 ( 
.A1(n_1505),
.A2(n_1539),
.B(n_1492),
.C(n_1437),
.Y(n_1652)
);

O2A1O1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1521),
.A2(n_1496),
.B(n_1473),
.C(n_1501),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1446),
.Y(n_1654)
);

A2O1A1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1442),
.A2(n_1485),
.B(n_1520),
.C(n_1541),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1446),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1488),
.B(n_1502),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1491),
.B(n_1494),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1452),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1541),
.A2(n_1447),
.B(n_1425),
.C(n_1452),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1446),
.B(n_1473),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1521),
.A2(n_1533),
.B1(n_1528),
.B2(n_1470),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1481),
.B(n_1452),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1481),
.B(n_1475),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1452),
.Y(n_1665)
);

O2A1O1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1428),
.A2(n_1490),
.B(n_1533),
.C(n_1475),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1528),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1484),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1482),
.B(n_1470),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1481),
.B(n_1479),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1484),
.A2(n_1482),
.B1(n_1479),
.B2(n_1510),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1479),
.B(n_1527),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1532),
.B(n_1538),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1561),
.B(n_1547),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1551),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1504),
.A2(n_1408),
.B(n_1399),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1414),
.Y(n_1677)
);

CKINVDCx20_ASAP7_75t_R g1678 ( 
.A(n_1451),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1446),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1504),
.A2(n_1408),
.B(n_1399),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1562),
.A2(n_1566),
.B1(n_906),
.B2(n_743),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1415),
.B(n_1500),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1512),
.B(n_1524),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1523),
.A2(n_1411),
.B(n_1408),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1523),
.A2(n_1411),
.B(n_1408),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1415),
.B(n_1500),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1509),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1414),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1631),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1569),
.B(n_1682),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1631),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1657),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1641),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1570),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1573),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1604),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1572),
.Y(n_1697)
);

INVx4_ASAP7_75t_L g1698 ( 
.A(n_1657),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1681),
.A2(n_1571),
.B1(n_1574),
.B2(n_1576),
.Y(n_1699)
);

OR2x6_ASAP7_75t_L g1700 ( 
.A(n_1620),
.B(n_1639),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1657),
.B(n_1569),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1682),
.B(n_1686),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1686),
.B(n_1586),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1586),
.B(n_1598),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1575),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1668),
.Y(n_1706)
);

OAI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1585),
.A2(n_1581),
.B1(n_1571),
.B2(n_1587),
.C(n_1643),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1596),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1579),
.B(n_1589),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1598),
.B(n_1597),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1647),
.Y(n_1711)
);

INVx4_ASAP7_75t_L g1712 ( 
.A(n_1611),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1597),
.B(n_1599),
.Y(n_1713)
);

AO21x2_ASAP7_75t_L g1714 ( 
.A1(n_1601),
.A2(n_1609),
.B(n_1633),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1605),
.B(n_1583),
.Y(n_1715)
);

BUFx4f_ASAP7_75t_SL g1716 ( 
.A(n_1590),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1604),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1588),
.B(n_1599),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1644),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1584),
.B(n_1683),
.Y(n_1720)
);

INVx4_ASAP7_75t_L g1721 ( 
.A(n_1611),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1600),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1636),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1603),
.B(n_1614),
.Y(n_1724)
);

OR2x6_ASAP7_75t_L g1725 ( 
.A(n_1635),
.B(n_1684),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1628),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1676),
.A2(n_1680),
.B(n_1685),
.Y(n_1727)
);

OA21x2_ASAP7_75t_L g1728 ( 
.A1(n_1655),
.A2(n_1660),
.B(n_1652),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1585),
.B(n_1688),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1646),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1663),
.B(n_1659),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1665),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1612),
.Y(n_1733)
);

AO21x1_ASAP7_75t_L g1734 ( 
.A1(n_1591),
.A2(n_1621),
.B(n_1608),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1580),
.B(n_1595),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1613),
.B(n_1619),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1626),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1623),
.B(n_1616),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1640),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1658),
.B(n_1664),
.Y(n_1740)
);

AOI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1592),
.A2(n_1627),
.B1(n_1582),
.B2(n_1615),
.C(n_1664),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1632),
.B(n_1638),
.Y(n_1742)
);

AO21x2_ASAP7_75t_L g1743 ( 
.A1(n_1660),
.A2(n_1651),
.B(n_1645),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1658),
.B(n_1677),
.Y(n_1744)
);

OAI211xp5_ASAP7_75t_L g1745 ( 
.A1(n_1653),
.A2(n_1622),
.B(n_1661),
.C(n_1666),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1628),
.A2(n_1616),
.B1(n_1642),
.B2(n_1624),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1625),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1733),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1706),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1706),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1699),
.A2(n_1734),
.B1(n_1707),
.B2(n_1727),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1690),
.B(n_1672),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1692),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1702),
.B(n_1670),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1702),
.B(n_1577),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1733),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1710),
.B(n_1577),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1737),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1718),
.B(n_1671),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1718),
.B(n_1577),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1710),
.B(n_1713),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1713),
.B(n_1740),
.Y(n_1762)
);

AND2x4_ASAP7_75t_SL g1763 ( 
.A(n_1700),
.B(n_1642),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1692),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1692),
.B(n_1674),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1740),
.B(n_1618),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1689),
.B(n_1618),
.Y(n_1767)
);

AOI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1699),
.A2(n_1661),
.B1(n_1656),
.B2(n_1654),
.C(n_1578),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1741),
.A2(n_1649),
.B(n_1679),
.C(n_1593),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1698),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1703),
.B(n_1675),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1703),
.B(n_1618),
.Y(n_1772)
);

BUFx3_ASAP7_75t_L g1773 ( 
.A(n_1719),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1698),
.B(n_1674),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1747),
.B(n_1648),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1732),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1744),
.B(n_1610),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1698),
.Y(n_1778)
);

BUFx4f_ASAP7_75t_L g1779 ( 
.A(n_1700),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1724),
.B(n_1673),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1691),
.B(n_1634),
.Y(n_1781)
);

CKINVDCx16_ASAP7_75t_R g1782 ( 
.A(n_1751),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1751),
.A2(n_1734),
.B1(n_1725),
.B2(n_1700),
.Y(n_1783)
);

O2A1O1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1769),
.A2(n_1725),
.B(n_1729),
.C(n_1700),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1780),
.B(n_1724),
.Y(n_1785)
);

AOI211xp5_ASAP7_75t_SL g1786 ( 
.A1(n_1768),
.A2(n_1745),
.B(n_1729),
.C(n_1716),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1777),
.B(n_1722),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1749),
.Y(n_1788)
);

NOR2x2_ASAP7_75t_L g1789 ( 
.A(n_1768),
.B(n_1725),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1779),
.A2(n_1725),
.B1(n_1700),
.B2(n_1735),
.C(n_1709),
.Y(n_1790)
);

AND2x4_ASAP7_75t_SL g1791 ( 
.A(n_1761),
.B(n_1726),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1773),
.Y(n_1792)
);

NOR2x1_ASAP7_75t_R g1793 ( 
.A(n_1753),
.B(n_1590),
.Y(n_1793)
);

AOI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1759),
.A2(n_1723),
.B1(n_1715),
.B2(n_1694),
.C(n_1708),
.Y(n_1794)
);

INVx4_ASAP7_75t_L g1795 ( 
.A(n_1779),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1765),
.B(n_1774),
.Y(n_1796)
);

OAI211xp5_ASAP7_75t_SL g1797 ( 
.A1(n_1759),
.A2(n_1715),
.B(n_1723),
.C(n_1720),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1775),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1765),
.B(n_1701),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_R g1800 ( 
.A(n_1779),
.B(n_1594),
.Y(n_1800)
);

NAND2xp33_ASAP7_75t_R g1801 ( 
.A(n_1778),
.B(n_1607),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1779),
.A2(n_1602),
.B1(n_1695),
.B2(n_1705),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1748),
.Y(n_1803)
);

OAI322xp33_ASAP7_75t_L g1804 ( 
.A1(n_1760),
.A2(n_1736),
.A3(n_1742),
.B1(n_1730),
.B2(n_1731),
.C1(n_1739),
.C2(n_1744),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1777),
.B(n_1704),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1760),
.B(n_1717),
.C(n_1746),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1775),
.A2(n_1742),
.B(n_1736),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1765),
.B(n_1701),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1780),
.B(n_1704),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1763),
.A2(n_1743),
.B(n_1728),
.Y(n_1810)
);

OAI31xp33_ASAP7_75t_L g1811 ( 
.A1(n_1763),
.A2(n_1662),
.A3(n_1617),
.B(n_1630),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_R g1812 ( 
.A(n_1770),
.B(n_1606),
.Y(n_1812)
);

OAI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1771),
.A2(n_1629),
.B1(n_1593),
.B2(n_1650),
.C(n_1687),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1748),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1756),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1761),
.B(n_1701),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1761),
.B(n_1738),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1756),
.Y(n_1818)
);

NOR4xp25_ASAP7_75t_SL g1819 ( 
.A(n_1778),
.B(n_1637),
.C(n_1607),
.D(n_1693),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1762),
.B(n_1738),
.Y(n_1820)
);

NAND3xp33_ASAP7_75t_L g1821 ( 
.A(n_1771),
.B(n_1728),
.C(n_1730),
.Y(n_1821)
);

AOI211xp5_ASAP7_75t_L g1822 ( 
.A1(n_1757),
.A2(n_1687),
.B(n_1650),
.C(n_1726),
.Y(n_1822)
);

AND2x6_ASAP7_75t_SL g1823 ( 
.A(n_1762),
.B(n_1669),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1758),
.A2(n_1602),
.B1(n_1606),
.B2(n_1678),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1750),
.Y(n_1825)
);

OA21x2_ASAP7_75t_L g1826 ( 
.A1(n_1767),
.A2(n_1697),
.B(n_1711),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1773),
.Y(n_1827)
);

NOR3xp33_ASAP7_75t_L g1828 ( 
.A(n_1782),
.B(n_1637),
.C(n_1667),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1803),
.Y(n_1829)
);

INVx4_ASAP7_75t_L g1830 ( 
.A(n_1795),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1826),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1814),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1815),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1784),
.A2(n_1743),
.B(n_1728),
.Y(n_1834)
);

NOR3xp33_ASAP7_75t_L g1835 ( 
.A(n_1783),
.B(n_1721),
.C(n_1712),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1818),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1821),
.B(n_1767),
.Y(n_1837)
);

OA21x2_ASAP7_75t_L g1838 ( 
.A1(n_1810),
.A2(n_1772),
.B(n_1767),
.Y(n_1838)
);

INVx2_ASAP7_75t_SL g1839 ( 
.A(n_1791),
.Y(n_1839)
);

INVx4_ASAP7_75t_L g1840 ( 
.A(n_1795),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1788),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1786),
.B(n_1728),
.C(n_1696),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1796),
.B(n_1757),
.Y(n_1843)
);

NOR2x1_ASAP7_75t_L g1844 ( 
.A(n_1797),
.B(n_1773),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1813),
.B(n_1678),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1800),
.B(n_1726),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1798),
.B(n_1754),
.Y(n_1847)
);

OA21x2_ASAP7_75t_L g1848 ( 
.A1(n_1825),
.A2(n_1772),
.B(n_1766),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1809),
.Y(n_1849)
);

AO21x2_ASAP7_75t_L g1850 ( 
.A1(n_1806),
.A2(n_1714),
.B(n_1743),
.Y(n_1850)
);

OA21x2_ASAP7_75t_L g1851 ( 
.A1(n_1807),
.A2(n_1772),
.B(n_1766),
.Y(n_1851)
);

INVxp67_ASAP7_75t_SL g1852 ( 
.A(n_1792),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1804),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1812),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1799),
.Y(n_1855)
);

INVx4_ASAP7_75t_SL g1856 ( 
.A(n_1800),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1799),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1854),
.B(n_1796),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1831),
.Y(n_1859)
);

OA21x2_ASAP7_75t_L g1860 ( 
.A1(n_1834),
.A2(n_1781),
.B(n_1776),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1856),
.B(n_1812),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1854),
.B(n_1796),
.Y(n_1862)
);

NAND2x1_ASAP7_75t_L g1863 ( 
.A(n_1844),
.B(n_1799),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1855),
.B(n_1857),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1855),
.B(n_1808),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1849),
.B(n_1785),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1829),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1829),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1853),
.B(n_1794),
.Y(n_1869)
);

AO22x2_ASAP7_75t_L g1870 ( 
.A1(n_1853),
.A2(n_1827),
.B1(n_1795),
.B2(n_1764),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1832),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1844),
.B(n_1805),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1849),
.B(n_1787),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1845),
.B(n_1830),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_R g1875 ( 
.A(n_1830),
.B(n_1801),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1855),
.B(n_1808),
.Y(n_1876)
);

INVxp67_ASAP7_75t_SL g1877 ( 
.A(n_1852),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1832),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1849),
.B(n_1762),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1833),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1857),
.B(n_1808),
.Y(n_1881)
);

NAND3xp33_ASAP7_75t_L g1882 ( 
.A(n_1842),
.B(n_1824),
.C(n_1802),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1833),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1857),
.B(n_1791),
.Y(n_1884)
);

NAND4xp25_ASAP7_75t_SL g1885 ( 
.A(n_1842),
.B(n_1824),
.C(n_1822),
.D(n_1802),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1839),
.B(n_1816),
.Y(n_1886)
);

AOI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1834),
.A2(n_1790),
.B(n_1846),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1836),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1839),
.B(n_1817),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1839),
.B(n_1820),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1831),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1843),
.B(n_1752),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1828),
.B(n_1823),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1852),
.Y(n_1894)
);

AND2x4_ASAP7_75t_L g1895 ( 
.A(n_1856),
.B(n_1765),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1837),
.B(n_1851),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1831),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1873),
.B(n_1847),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1885),
.A2(n_1835),
.B1(n_1828),
.B2(n_1830),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1858),
.B(n_1843),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1867),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1858),
.B(n_1851),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1873),
.B(n_1847),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1862),
.B(n_1851),
.Y(n_1904)
);

INVx1_ASAP7_75t_SL g1905 ( 
.A(n_1875),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1866),
.B(n_1830),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1866),
.B(n_1840),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1862),
.B(n_1851),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_SL g1909 ( 
.A(n_1882),
.B(n_1793),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1895),
.B(n_1851),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1867),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1895),
.B(n_1856),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1894),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1868),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1868),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1871),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1895),
.B(n_1856),
.Y(n_1917)
);

NOR2x1_ASAP7_75t_L g1918 ( 
.A(n_1863),
.B(n_1840),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1871),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1869),
.B(n_1835),
.Y(n_1920)
);

AND2x4_ASAP7_75t_L g1921 ( 
.A(n_1895),
.B(n_1856),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1872),
.B(n_1840),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_1863),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1861),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1878),
.Y(n_1925)
);

OAI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1882),
.A2(n_1840),
.B1(n_1819),
.B2(n_1837),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1877),
.B(n_1757),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1893),
.B(n_1856),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1894),
.B(n_1841),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1892),
.B(n_1841),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1878),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1879),
.B(n_1850),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1874),
.B(n_1755),
.Y(n_1933)
);

NAND2x1_ASAP7_75t_L g1934 ( 
.A(n_1870),
.B(n_1848),
.Y(n_1934)
);

AND3x2_ASAP7_75t_L g1935 ( 
.A(n_1909),
.B(n_1811),
.C(n_1884),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1898),
.B(n_1879),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1920),
.B(n_1886),
.Y(n_1937)
);

INVx2_ASAP7_75t_SL g1938 ( 
.A(n_1921),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1903),
.B(n_1913),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1913),
.Y(n_1940)
);

NOR3xp33_ASAP7_75t_L g1941 ( 
.A(n_1928),
.B(n_1887),
.C(n_1896),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1900),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1901),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1928),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1900),
.B(n_1870),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1924),
.B(n_1886),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1905),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1911),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1918),
.B(n_1892),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1899),
.B(n_1889),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1912),
.B(n_1870),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1922),
.B(n_1889),
.Y(n_1952)
);

AOI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1926),
.A2(n_1850),
.B1(n_1876),
.B2(n_1865),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_1923),
.Y(n_1954)
);

NOR2x1_ASAP7_75t_L g1955 ( 
.A(n_1923),
.B(n_1896),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1923),
.Y(n_1956)
);

INVx1_ASAP7_75t_SL g1957 ( 
.A(n_1912),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1906),
.B(n_1890),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1907),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1914),
.B(n_1890),
.Y(n_1960)
);

XNOR2x1_ASAP7_75t_L g1961 ( 
.A(n_1947),
.B(n_1921),
.Y(n_1961)
);

AOI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1941),
.A2(n_1921),
.B1(n_1917),
.B2(n_1801),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1940),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1953),
.A2(n_1934),
.B(n_1917),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1949),
.B(n_1902),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1946),
.B(n_1937),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1942),
.B(n_1884),
.Y(n_1967)
);

OAI21xp33_ASAP7_75t_L g1968 ( 
.A1(n_1950),
.A2(n_1933),
.B(n_1927),
.Y(n_1968)
);

A2O1A1Ixp33_ASAP7_75t_L g1969 ( 
.A1(n_1955),
.A2(n_1902),
.B(n_1904),
.C(n_1908),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1944),
.A2(n_1870),
.B1(n_1931),
.B2(n_1916),
.C(n_1915),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1957),
.B(n_1919),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1940),
.Y(n_1972)
);

INVx1_ASAP7_75t_SL g1973 ( 
.A(n_1939),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1942),
.B(n_1865),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1959),
.B(n_1925),
.Y(n_1975)
);

O2A1O1Ixp33_ASAP7_75t_L g1976 ( 
.A1(n_1938),
.A2(n_1932),
.B(n_1904),
.C(n_1908),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_SL g1977 ( 
.A1(n_1938),
.A2(n_1860),
.B1(n_1789),
.B2(n_1838),
.Y(n_1977)
);

AOI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1952),
.A2(n_1910),
.B1(n_1850),
.B2(n_1929),
.C(n_1930),
.Y(n_1978)
);

O2A1O1Ixp33_ASAP7_75t_L g1979 ( 
.A1(n_1955),
.A2(n_1850),
.B(n_1910),
.C(n_1860),
.Y(n_1979)
);

OAI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1939),
.A2(n_1860),
.B(n_1929),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1973),
.B(n_1958),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1963),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1966),
.B(n_1960),
.Y(n_1983)
);

INVx2_ASAP7_75t_SL g1984 ( 
.A(n_1961),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1972),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1970),
.A2(n_1935),
.B1(n_1954),
.B2(n_1948),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1975),
.Y(n_1987)
);

NAND2xp33_ASAP7_75t_SL g1988 ( 
.A(n_1965),
.B(n_1954),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1971),
.Y(n_1989)
);

OA21x2_ASAP7_75t_L g1990 ( 
.A1(n_1980),
.A2(n_1956),
.B(n_1948),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1967),
.Y(n_1991)
);

OAI21xp33_ASAP7_75t_L g1992 ( 
.A1(n_1986),
.A2(n_1962),
.B(n_1968),
.Y(n_1992)
);

NOR3xp33_ASAP7_75t_L g1993 ( 
.A(n_1984),
.B(n_1964),
.C(n_1978),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1986),
.B(n_1949),
.Y(n_1994)
);

OAI221xp5_ASAP7_75t_L g1995 ( 
.A1(n_1988),
.A2(n_1964),
.B1(n_1977),
.B2(n_1969),
.C(n_1980),
.Y(n_1995)
);

AOI21xp33_ASAP7_75t_L g1996 ( 
.A1(n_1981),
.A2(n_1990),
.B(n_1983),
.Y(n_1996)
);

A2O1A1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1985),
.A2(n_1979),
.B(n_1976),
.C(n_1949),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1991),
.A2(n_1974),
.B1(n_1951),
.B2(n_1945),
.Y(n_1998)
);

NAND3xp33_ASAP7_75t_SL g1999 ( 
.A(n_1989),
.B(n_1951),
.C(n_1956),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1987),
.B(n_1982),
.Y(n_2000)
);

OAI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_1995),
.A2(n_1990),
.B1(n_1985),
.B2(n_1936),
.Y(n_2001)
);

INVx1_ASAP7_75t_SL g2002 ( 
.A(n_1994),
.Y(n_2002)
);

OAI21xp33_ASAP7_75t_SL g2003 ( 
.A1(n_1996),
.A2(n_1998),
.B(n_1945),
.Y(n_2003)
);

OAI221xp5_ASAP7_75t_L g2004 ( 
.A1(n_1997),
.A2(n_1990),
.B1(n_1943),
.B2(n_1936),
.C(n_1860),
.Y(n_2004)
);

NOR2x1_ASAP7_75t_L g2005 ( 
.A(n_1999),
.B(n_1943),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_2002),
.B(n_1992),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_2005),
.Y(n_2007)
);

NOR2xp67_ASAP7_75t_L g2008 ( 
.A(n_2004),
.B(n_2000),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_2003),
.B(n_1993),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_2001),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_2002),
.B(n_1876),
.Y(n_2011)
);

AOI221xp5_ASAP7_75t_L g2012 ( 
.A1(n_2010),
.A2(n_1929),
.B1(n_1859),
.B2(n_1891),
.C(n_1897),
.Y(n_2012)
);

AOI221x1_ASAP7_75t_L g2013 ( 
.A1(n_2007),
.A2(n_2009),
.B1(n_2011),
.B2(n_2008),
.C(n_2006),
.Y(n_2013)
);

INVx1_ASAP7_75t_SL g2014 ( 
.A(n_2008),
.Y(n_2014)
);

INVx1_ASAP7_75t_SL g2015 ( 
.A(n_2011),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_2009),
.A2(n_1864),
.B1(n_1930),
.B2(n_1881),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_SL g2017 ( 
.A(n_2015),
.B(n_1864),
.Y(n_2017)
);

AOI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_2014),
.A2(n_1891),
.B(n_1859),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2013),
.B(n_1930),
.Y(n_2019)
);

AND2x4_ASAP7_75t_L g2020 ( 
.A(n_2019),
.B(n_2016),
.Y(n_2020)
);

NOR3xp33_ASAP7_75t_L g2021 ( 
.A(n_2020),
.B(n_2018),
.C(n_2012),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2021),
.Y(n_2022)
);

NOR2xp67_ASAP7_75t_L g2023 ( 
.A(n_2021),
.B(n_2017),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2023),
.Y(n_2024)
);

BUFx2_ASAP7_75t_L g2025 ( 
.A(n_2022),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_2025),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_2026),
.Y(n_2027)
);

OA21x2_ASAP7_75t_L g2028 ( 
.A1(n_2027),
.A2(n_2024),
.B(n_1859),
.Y(n_2028)
);

OAI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_2028),
.A2(n_1891),
.B(n_1897),
.Y(n_2029)
);

XNOR2xp5_ASAP7_75t_L g2030 ( 
.A(n_2029),
.B(n_1881),
.Y(n_2030)
);

AOI221xp5_ASAP7_75t_L g2031 ( 
.A1(n_2030),
.A2(n_1897),
.B1(n_1880),
.B2(n_1883),
.C(n_1888),
.Y(n_2031)
);

AOI211xp5_ASAP7_75t_L g2032 ( 
.A1(n_2031),
.A2(n_1880),
.B(n_1888),
.C(n_1883),
.Y(n_2032)
);


endmodule