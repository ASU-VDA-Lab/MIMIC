module real_jpeg_1132_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_2),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_2),
.A2(n_51),
.B1(n_52),
.B2(n_80),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_2),
.A2(n_37),
.B1(n_43),
.B2(n_80),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_30),
.B1(n_33),
.B2(n_61),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_3),
.A2(n_37),
.B1(n_43),
.B2(n_61),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_6),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_6),
.A2(n_42),
.B1(n_51),
.B2(n_52),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_7),
.A2(n_37),
.B1(n_43),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_7),
.Y(n_109)
);

BUFx16f_ASAP7_75t_L g86 ( 
.A(n_8),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_10),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_83),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_10),
.A2(n_37),
.B1(n_43),
.B2(n_83),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_11),
.B(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_11),
.A2(n_32),
.B(n_33),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_11),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_11),
.B(n_50),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_11),
.A2(n_24),
.B(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_11),
.B(n_37),
.C(n_86),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_126),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_11),
.B(n_40),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_11),
.B(n_91),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_13),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_14),
.A2(n_30),
.B1(n_33),
.B2(n_58),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_14),
.A2(n_51),
.B1(n_52),
.B2(n_58),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_14),
.A2(n_37),
.B1(n_43),
.B2(n_58),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_15),
.A2(n_37),
.B1(n_43),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_15),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_15),
.A2(n_51),
.B1(n_52),
.B2(n_69),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_115),
.B1(n_187),
.B2(n_188),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_19),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_94),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_21),
.B(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_21),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_21),
.B(n_117),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_47),
.CI(n_70),
.CON(n_21),
.SN(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_23),
.B(n_35),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.A3(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_24),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_24),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_65)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_24),
.A2(n_52),
.A3(n_54),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_25),
.B(n_126),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_36),
.A2(n_40),
.B1(n_41),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_36),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_36),
.A2(n_40),
.B1(n_130),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_36),
.A2(n_40),
.B1(n_126),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_36),
.A2(n_40),
.B1(n_167),
.B2(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_37),
.A2(n_43),
.B1(n_86),
.B2(n_87),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_37),
.B(n_165),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_39),
.A2(n_45),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_39),
.A2(n_107),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_39),
.A2(n_107),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_62),
.C(n_66),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_48),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_59),
.B1(n_60),
.B2(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_49),
.A2(n_59),
.B1(n_79),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_49),
.A2(n_57),
.B1(n_59),
.B2(n_146),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

AO22x2_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_52),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_51),
.B(n_55),
.Y(n_127)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_52),
.B(n_155),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_119)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_65),
.A2(n_72),
.B1(n_76),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_78),
.C(n_93),
.Y(n_113)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_92),
.B2(n_93),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_89),
.B2(n_91),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_84),
.B1(n_91),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_84),
.A2(n_91),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_84),
.A2(n_91),
.B1(n_137),
.B2(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_90),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_88),
.A2(n_111),
.B1(n_122),
.B2(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_113),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_132),
.B(n_186),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.C(n_123),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_118),
.B(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_123),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_181),
.B(n_185),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_150),
.B(n_180),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_142),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_142),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_140),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_139),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_145),
.C(n_148),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_161),
.B(n_179),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_159),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_173),
.B(n_178),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_168),
.B(n_172),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_177),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_184),
.Y(n_185)
);


endmodule