module fake_jpeg_13460_n_171 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_4),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_37),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_31),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_3),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_2),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_0),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_71),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_97),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_54),
.B1(n_72),
.B2(n_49),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_87),
.B1(n_94),
.B2(n_64),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_54),
.B1(n_72),
.B2(n_49),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_67),
.B1(n_69),
.B2(n_57),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_64),
.B1(n_51),
.B2(n_4),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_68),
.B1(n_70),
.B2(n_53),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_98),
.B1(n_51),
.B2(n_5),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_75),
.A2(n_53),
.B1(n_51),
.B2(n_64),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_85),
.B1(n_91),
.B2(n_84),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_101),
.B1(n_110),
.B2(n_114),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_112),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_76),
.B1(n_77),
.B2(n_65),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_106),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_56),
.B(n_55),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_18),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_0),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_111),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_1),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_2),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_3),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_119),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_9),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_8),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_23),
.A3(n_46),
.B1(n_44),
.B2(n_43),
.Y(n_124)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_9),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_21),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

CKINVDCx12_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_20),
.C(n_42),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_137),
.C(n_139),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_22),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_139),
.B(n_12),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_118),
.B1(n_10),
.B2(n_11),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_138),
.B1(n_123),
.B2(n_127),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_17),
.B1(n_41),
.B2(n_39),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_151),
.B(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_124),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_149),
.C(n_132),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_47),
.C(n_26),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_130),
.C(n_125),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_157),
.C(n_161),
.Y(n_163)
);

XNOR2x2_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_134),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_158),
.A2(n_159),
.B(n_160),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

OA21x2_ASAP7_75t_SL g165 ( 
.A1(n_162),
.A2(n_147),
.B(n_142),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_166),
.C(n_152),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_164),
.A2(n_152),
.B1(n_120),
.B2(n_159),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_145),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_150),
.A3(n_140),
.B1(n_163),
.B2(n_154),
.C1(n_155),
.C2(n_149),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_148),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_35),
.Y(n_171)
);


endmodule