module fake_netlist_1_4686_n_522 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_522);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_522;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g68 ( .A(n_52), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_61), .Y(n_69) );
CKINVDCx5p33_ASAP7_75t_R g70 ( .A(n_42), .Y(n_70) );
INVxp67_ASAP7_75t_SL g71 ( .A(n_18), .Y(n_71) );
INVxp67_ASAP7_75t_SL g72 ( .A(n_67), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_29), .Y(n_73) );
INVx2_ASAP7_75t_L g74 ( .A(n_47), .Y(n_74) );
CKINVDCx5p33_ASAP7_75t_R g75 ( .A(n_55), .Y(n_75) );
BUFx3_ASAP7_75t_L g76 ( .A(n_35), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_56), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_53), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_57), .Y(n_79) );
BUFx3_ASAP7_75t_L g80 ( .A(n_39), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_48), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_2), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_58), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_33), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_62), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_1), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_41), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_6), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_37), .Y(n_89) );
CKINVDCx14_ASAP7_75t_R g90 ( .A(n_46), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_28), .Y(n_91) );
BUFx2_ASAP7_75t_L g92 ( .A(n_23), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_16), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_34), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_20), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_66), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_9), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_36), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_65), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_38), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_63), .Y(n_101) );
INVx3_ASAP7_75t_L g102 ( .A(n_59), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_3), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_40), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_21), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_68), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_92), .B(n_0), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_92), .B(n_0), .Y(n_108) );
INVx3_ASAP7_75t_L g109 ( .A(n_102), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_102), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_102), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_68), .Y(n_112) );
AND2x4_ASAP7_75t_L g113 ( .A(n_102), .B(n_1), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_69), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_74), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_76), .Y(n_116) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_69), .A2(n_24), .B(n_64), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
INVx2_ASAP7_75t_SL g119 ( .A(n_76), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_74), .Y(n_120) );
INVx4_ASAP7_75t_L g121 ( .A(n_76), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_73), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_105), .B(n_2), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_90), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_81), .B(n_3), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_81), .B(n_4), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_82), .B(n_4), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_78), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_83), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_78), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_109), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_124), .B(n_70), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_109), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_113), .Y(n_138) );
BUFx4f_ASAP7_75t_L g139 ( .A(n_113), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_124), .B(n_96), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_116), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_108), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_109), .B(n_75), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_108), .B(n_88), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
BUFx4f_ASAP7_75t_L g146 ( .A(n_113), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_113), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_109), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_116), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_106), .B(n_88), .Y(n_150) );
INVx1_ASAP7_75t_SL g151 ( .A(n_107), .Y(n_151) );
OAI22xp33_ASAP7_75t_L g152 ( .A1(n_106), .A2(n_86), .B1(n_82), .B2(n_103), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_112), .Y(n_153) );
OR2x2_ASAP7_75t_L g154 ( .A(n_134), .B(n_103), .Y(n_154) );
INVx4_ASAP7_75t_SL g155 ( .A(n_116), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_116), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_116), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_121), .B(n_80), .Y(n_158) );
BUFx2_ASAP7_75t_L g159 ( .A(n_121), .Y(n_159) );
INVxp67_ASAP7_75t_SL g160 ( .A(n_110), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_110), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_129), .A2(n_86), .B1(n_91), .B2(n_89), .Y(n_162) );
HB1xp67_ASAP7_75t_SL g163 ( .A(n_129), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_112), .B(n_80), .Y(n_164) );
AND2x6_ASAP7_75t_L g165 ( .A(n_110), .B(n_93), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_114), .B(n_83), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_151), .A2(n_123), .B1(n_134), .B2(n_114), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_153), .B(n_133), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_161), .Y(n_171) );
OR2x2_ASAP7_75t_L g172 ( .A(n_142), .B(n_133), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_139), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_135), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_139), .A2(n_131), .B1(n_118), .B2(n_127), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
BUFx8_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
OR2x2_ASAP7_75t_SL g178 ( .A(n_163), .B(n_117), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_147), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_147), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
OAI22xp33_ASAP7_75t_L g182 ( .A1(n_142), .A2(n_97), .B1(n_131), .B2(n_127), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_136), .B(n_122), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_146), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_146), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_165), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_165), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_135), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_150), .B(n_160), .Y(n_191) );
NOR2xp33_ASAP7_75t_R g192 ( .A(n_140), .B(n_119), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_137), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_137), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_148), .Y(n_195) );
NOR2xp67_ASAP7_75t_L g196 ( .A(n_162), .B(n_111), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_138), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_154), .A2(n_118), .B1(n_125), .B2(n_122), .Y(n_198) );
INVx5_ASAP7_75t_L g199 ( .A(n_165), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_141), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_152), .B(n_125), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_165), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_145), .Y(n_203) );
NOR2x1p5_ASAP7_75t_L g204 ( .A(n_154), .B(n_126), .Y(n_204) );
BUFx2_ASAP7_75t_L g205 ( .A(n_165), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_165), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_150), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_143), .B(n_121), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_199), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_172), .B(n_159), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_168), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_181), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_177), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_181), .Y(n_214) );
BUFx12f_ASAP7_75t_L g215 ( .A(n_177), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_184), .A2(n_164), .B1(n_166), .B2(n_119), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_171), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_171), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_177), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_181), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_186), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_186), .B(n_128), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_168), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_172), .B(n_159), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_174), .Y(n_225) );
AOI21x1_ASAP7_75t_L g226 ( .A1(n_197), .A2(n_158), .B(n_149), .Y(n_226) );
NAND2x1p5_ASAP7_75t_L g227 ( .A(n_186), .B(n_111), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_185), .Y(n_228) );
INVx1_ASAP7_75t_SL g229 ( .A(n_183), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_204), .A2(n_121), .B1(n_111), .B2(n_115), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_179), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_196), .A2(n_115), .B1(n_132), .B2(n_120), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_199), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_207), .B(n_132), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_207), .A2(n_120), .B1(n_72), .B2(n_94), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_170), .B(n_120), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_191), .Y(n_237) );
OR2x6_ASAP7_75t_L g238 ( .A(n_187), .B(n_101), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_187), .B(n_71), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_187), .B(n_105), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_185), .Y(n_241) );
BUFx2_ASAP7_75t_SL g242 ( .A(n_199), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_188), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_199), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_179), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_237), .A2(n_182), .B1(n_201), .B2(n_173), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_240), .A2(n_197), .B(n_176), .C(n_180), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_229), .B(n_173), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_213), .B(n_198), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_223), .B(n_169), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_213), .B(n_176), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_223), .B(n_175), .Y(n_252) );
INVx1_ASAP7_75t_SL g253 ( .A(n_238), .Y(n_253) );
OAI22xp33_ASAP7_75t_L g254 ( .A1(n_215), .A2(n_176), .B1(n_180), .B2(n_174), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_217), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_215), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_217), .B(n_180), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_218), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_238), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_238), .A2(n_194), .B1(n_190), .B2(n_193), .Y(n_260) );
AOI21x1_ASAP7_75t_L g261 ( .A1(n_226), .A2(n_141), .B(n_149), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_212), .Y(n_262) );
OAI22xp5_ASAP7_75t_SL g263 ( .A1(n_219), .A2(n_178), .B1(n_117), .B2(n_84), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_211), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_238), .A2(n_194), .B1(n_190), .B2(n_193), .Y(n_265) );
AOI222xp33_ASAP7_75t_L g266 ( .A1(n_219), .A2(n_195), .B1(n_100), .B2(n_99), .C1(n_85), .C2(n_79), .Y(n_266) );
AOI22xp33_ASAP7_75t_SL g267 ( .A1(n_210), .A2(n_192), .B1(n_205), .B2(n_195), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_224), .B(n_205), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_211), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_218), .B(n_189), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_212), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_266), .B(n_234), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_246), .A2(n_232), .B1(n_235), .B2(n_234), .C(n_230), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_268), .A2(n_238), .B1(n_222), .B2(n_239), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_250), .A2(n_225), .B1(n_239), .B2(n_235), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_264), .Y(n_276) );
OAI21xp33_ASAP7_75t_L g277 ( .A1(n_266), .A2(n_216), .B(n_236), .Y(n_277) );
BUFx2_ASAP7_75t_R g278 ( .A(n_256), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_250), .A2(n_225), .B1(n_239), .B2(n_216), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_249), .B(n_239), .Y(n_280) );
OAI33xp33_ASAP7_75t_L g281 ( .A1(n_263), .A2(n_99), .A3(n_84), .B1(n_85), .B2(n_87), .B3(n_93), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_255), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_249), .B(n_222), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_264), .Y(n_284) );
OAI22xp33_ASAP7_75t_L g285 ( .A1(n_253), .A2(n_227), .B1(n_245), .B2(n_231), .Y(n_285) );
AOI22xp33_ASAP7_75t_SL g286 ( .A1(n_253), .A2(n_220), .B1(n_221), .B2(n_214), .Y(n_286) );
AOI221x1_ASAP7_75t_SL g287 ( .A1(n_255), .A2(n_101), .B1(n_100), .B2(n_98), .C(n_95), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_248), .B(n_227), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g289 ( .A1(n_251), .A2(n_222), .B1(n_214), .B2(n_220), .C(n_221), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_252), .A2(n_222), .B1(n_214), .B2(n_220), .C(n_221), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_258), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_264), .Y(n_292) );
INVx8_ASAP7_75t_L g293 ( .A(n_262), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_282), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_283), .B(n_258), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_276), .B(n_269), .Y(n_296) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_275), .A2(n_267), .B(n_259), .C(n_95), .Y(n_297) );
INVx11_ASAP7_75t_L g298 ( .A(n_278), .Y(n_298) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_285), .A2(n_261), .B(n_226), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_291), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_277), .A2(n_252), .B1(n_263), .B2(n_265), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_272), .A2(n_260), .B1(n_254), .B2(n_257), .Y(n_302) );
INVx4_ASAP7_75t_L g303 ( .A(n_293), .Y(n_303) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_287), .A2(n_257), .B1(n_247), .B2(n_270), .C(n_98), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_279), .A2(n_270), .B(n_227), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_293), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_276), .Y(n_307) );
NAND3xp33_ASAP7_75t_L g308 ( .A(n_275), .B(n_87), .C(n_130), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_280), .B(n_269), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_274), .A2(n_269), .B1(n_271), .B2(n_262), .Y(n_310) );
OR2x6_ASAP7_75t_L g311 ( .A(n_293), .B(n_242), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_288), .B(n_271), .Y(n_312) );
AOI33xp33_ASAP7_75t_L g313 ( .A1(n_279), .A2(n_104), .A3(n_6), .B1(n_7), .B2(n_8), .B3(n_9), .Y(n_313) );
CKINVDCx14_ASAP7_75t_R g314 ( .A(n_284), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_292), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_292), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_290), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_284), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_273), .A2(n_271), .B1(n_262), .B2(n_228), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_294), .B(n_284), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_307), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_312), .B(n_284), .Y(n_322) );
INVx4_ASAP7_75t_L g323 ( .A(n_311), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_313), .B(n_285), .Y(n_324) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_313), .B(n_104), .C(n_289), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_304), .A2(n_281), .B1(n_130), .B2(n_271), .C(n_262), .Y(n_326) );
OAI31xp33_ASAP7_75t_SL g327 ( .A1(n_297), .A2(n_286), .A3(n_178), .B(n_8), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_315), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_317), .A2(n_220), .B1(n_221), .B2(n_212), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_300), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_316), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_309), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_296), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
NAND3xp33_ASAP7_75t_SL g335 ( .A(n_303), .B(n_5), .C(n_7), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_318), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_311), .B(n_305), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_306), .Y(n_338) );
INVx2_ASAP7_75t_SL g339 ( .A(n_298), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_295), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_295), .B(n_5), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_299), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_314), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_299), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_314), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_301), .A2(n_130), .B1(n_212), .B2(n_214), .C(n_245), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_302), .B(n_10), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_311), .B(n_261), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_308), .A2(n_310), .B1(n_319), .B2(n_306), .C(n_130), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_299), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_311), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_306), .Y(n_352) );
OAI31xp33_ASAP7_75t_SL g353 ( .A1(n_298), .A2(n_10), .A3(n_11), .B(n_12), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_303), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_303), .A2(n_228), .B1(n_241), .B2(n_231), .Y(n_355) );
NOR2x1_ASAP7_75t_R g356 ( .A(n_303), .B(n_242), .Y(n_356) );
NAND3xp33_ASAP7_75t_L g357 ( .A(n_313), .B(n_130), .C(n_167), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_330), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_321), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_331), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_340), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_348), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_328), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_337), .B(n_60), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_333), .B(n_12), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_334), .B(n_13), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_332), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_342), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_336), .B(n_13), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_336), .B(n_14), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_337), .B(n_117), .Y(n_372) );
AO21x2_ASAP7_75t_L g373 ( .A1(n_342), .A2(n_156), .B(n_157), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_354), .Y(n_374) );
AND2x4_ASAP7_75t_SL g375 ( .A(n_323), .B(n_244), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g376 ( .A(n_323), .B(n_241), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_322), .Y(n_377) );
NAND4xp25_ASAP7_75t_L g378 ( .A(n_353), .B(n_156), .C(n_157), .D(n_14), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_320), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_344), .Y(n_380) );
OAI21xp33_ASAP7_75t_L g381 ( .A1(n_327), .A2(n_145), .B(n_167), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_338), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_343), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_337), .B(n_117), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_341), .B(n_167), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_344), .B(n_167), .Y(n_386) );
INVx2_ASAP7_75t_SL g387 ( .A(n_323), .Y(n_387) );
NAND3xp33_ASAP7_75t_SL g388 ( .A(n_357), .B(n_206), .C(n_202), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_356), .Y(n_389) );
AND4x1_ASAP7_75t_L g390 ( .A(n_325), .B(n_15), .C(n_17), .D(n_19), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_350), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_345), .B(n_145), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_338), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_348), .B(n_145), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_351), .B(n_145), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_352), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_347), .B(n_241), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_324), .B(n_22), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_324), .B(n_228), .Y(n_399) );
AOI21xp33_ASAP7_75t_SL g400 ( .A1(n_339), .A2(n_25), .B(n_26), .Y(n_400) );
AND4x1_ASAP7_75t_L g401 ( .A(n_326), .B(n_27), .C(n_30), .D(n_31), .Y(n_401) );
NOR2x1_ASAP7_75t_L g402 ( .A(n_335), .B(n_233), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_329), .B(n_32), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_383), .B(n_355), .Y(n_404) );
NOR3xp33_ASAP7_75t_L g405 ( .A(n_378), .B(n_349), .C(n_346), .Y(n_405) );
NAND2x1_ASAP7_75t_L g406 ( .A(n_389), .B(n_244), .Y(n_406) );
NOR4xp75_ASAP7_75t_L g407 ( .A(n_381), .B(n_43), .C(n_44), .D(n_45), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_361), .B(n_49), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_358), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_382), .B(n_244), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_377), .B(n_50), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_360), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_393), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_368), .B(n_51), .Y(n_414) );
INVxp33_ASAP7_75t_L g415 ( .A(n_366), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_374), .B(n_54), .Y(n_416) );
OR2x6_ASAP7_75t_L g417 ( .A(n_387), .B(n_244), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_364), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_379), .B(n_206), .Y(n_419) );
OAI21xp5_ASAP7_75t_L g420 ( .A1(n_402), .A2(n_202), .B(n_208), .Y(n_420) );
NAND2xp33_ASAP7_75t_R g421 ( .A(n_365), .B(n_188), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_359), .B(n_155), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_396), .B(n_155), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_396), .B(n_155), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_363), .B(n_366), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_370), .B(n_243), .Y(n_426) );
NAND2xp33_ASAP7_75t_SL g427 ( .A(n_387), .B(n_244), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_370), .B(n_371), .C(n_398), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_388), .A2(n_244), .B(n_233), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_371), .B(n_203), .C(n_199), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_369), .Y(n_431) );
AND3x2_ASAP7_75t_L g432 ( .A(n_365), .B(n_200), .C(n_209), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_394), .B(n_203), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_367), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_392), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_369), .B(n_200), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_362), .B(n_391), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_380), .B(n_188), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_397), .B(n_243), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_395), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_365), .B(n_243), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_398), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
O2A1O1Ixp33_ASAP7_75t_L g444 ( .A1(n_405), .A2(n_400), .B(n_399), .C(n_385), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_412), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_413), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_418), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_425), .Y(n_448) );
XOR2x2_ASAP7_75t_L g449 ( .A(n_428), .B(n_390), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_413), .B(n_362), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_435), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_431), .Y(n_452) );
XNOR2xp5_ASAP7_75t_L g453 ( .A(n_415), .B(n_401), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_434), .B(n_362), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_427), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_404), .B(n_375), .Y(n_456) );
INVx2_ASAP7_75t_SL g457 ( .A(n_417), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_437), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_440), .B(n_372), .Y(n_459) );
OAI21xp5_ASAP7_75t_SL g460 ( .A1(n_432), .A2(n_375), .B(n_376), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_442), .B(n_384), .Y(n_461) );
NAND2x1_ASAP7_75t_L g462 ( .A(n_417), .B(n_391), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_417), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_410), .B(n_376), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_421), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_436), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_436), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_411), .Y(n_468) );
OAI32xp33_ASAP7_75t_L g469 ( .A1(n_416), .A2(n_403), .A3(n_386), .B1(n_373), .B2(n_189), .Y(n_469) );
OAI22xp33_ASAP7_75t_L g470 ( .A1(n_430), .A2(n_403), .B1(n_373), .B2(n_209), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_406), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_426), .A2(n_373), .B1(n_189), .B2(n_209), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_408), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_408), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_438), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_438), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_419), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_414), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_433), .Y(n_479) );
OAI21xp5_ASAP7_75t_SL g480 ( .A1(n_420), .A2(n_209), .B(n_233), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_420), .A2(n_439), .B(n_422), .C(n_441), .Y(n_481) );
AO22x2_ASAP7_75t_L g482 ( .A1(n_423), .A2(n_233), .B1(n_424), .B2(n_429), .Y(n_482) );
XOR2x2_ASAP7_75t_L g483 ( .A(n_407), .B(n_233), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_427), .B(n_233), .Y(n_484) );
NAND2xp33_ASAP7_75t_SL g485 ( .A(n_421), .B(n_406), .Y(n_485) );
AOI31xp33_ASAP7_75t_L g486 ( .A1(n_421), .A2(n_356), .A3(n_354), .B(n_415), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_413), .B(n_377), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_409), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_427), .B(n_413), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_449), .A2(n_456), .B1(n_454), .B2(n_465), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_449), .A2(n_456), .B1(n_453), .B2(n_457), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_443), .Y(n_492) );
OAI221xp5_ASAP7_75t_R g493 ( .A1(n_486), .A2(n_489), .B1(n_485), .B2(n_472), .C(n_450), .Y(n_493) );
NAND3xp33_ASAP7_75t_L g494 ( .A(n_446), .B(n_489), .C(n_444), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_446), .B(n_478), .C(n_450), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_487), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_455), .A2(n_471), .B1(n_484), .B2(n_462), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_448), .B(n_451), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_454), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_452), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_485), .A2(n_482), .B1(n_463), .B2(n_459), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_452), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_496), .Y(n_503) );
NAND5xp2_ASAP7_75t_L g504 ( .A(n_491), .B(n_460), .C(n_481), .D(n_480), .E(n_473), .Y(n_504) );
XOR2x2_ASAP7_75t_L g505 ( .A(n_490), .B(n_494), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_499), .B(n_474), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_492), .B(n_495), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_501), .A2(n_484), .B1(n_468), .B2(n_482), .Y(n_508) );
OAI211xp5_ASAP7_75t_L g509 ( .A1(n_497), .A2(n_464), .B(n_469), .C(n_461), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_503), .Y(n_510) );
OR5x1_ASAP7_75t_L g511 ( .A(n_509), .B(n_493), .C(n_498), .D(n_482), .E(n_470), .Y(n_511) );
INVxp67_ASAP7_75t_SL g512 ( .A(n_507), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g513 ( .A(n_504), .B(n_493), .C(n_464), .Y(n_513) );
NOR3xp33_ASAP7_75t_SL g514 ( .A(n_512), .B(n_508), .C(n_505), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_513), .A2(n_506), .B1(n_476), .B2(n_467), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_510), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_514), .A2(n_511), .B1(n_445), .B2(n_488), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_516), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_518), .A2(n_515), .B(n_483), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_519), .A2(n_517), .B1(n_477), .B2(n_502), .Y(n_520) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_520), .A2(n_500), .B1(n_447), .B2(n_458), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_521), .A2(n_479), .B1(n_475), .B2(n_466), .Y(n_522) );
endmodule