module fake_jpeg_31499_n_502 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_502);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_502;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_SL g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_56),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_58),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_59),
.Y(n_139)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_14),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_79),
.Y(n_127)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_14),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_96),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_14),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_103),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_18),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_16),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g130 ( 
.A(n_104),
.Y(n_130)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_105),
.B(n_44),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_39),
.B1(n_48),
.B2(n_25),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_121),
.B(n_74),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_52),
.A2(n_18),
.B1(n_36),
.B2(n_31),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_155),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_61),
.A2(n_18),
.B1(n_36),
.B2(n_46),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_132),
.A2(n_140),
.B1(n_165),
.B2(n_25),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_67),
.A2(n_36),
.B1(n_50),
.B2(n_31),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_80),
.A2(n_34),
.B1(n_50),
.B2(n_22),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_136),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_58),
.B(n_26),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_138),
.B(n_29),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_93),
.A2(n_46),
.B1(n_39),
.B2(n_20),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_81),
.A2(n_22),
.B1(n_34),
.B2(n_26),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_83),
.A2(n_46),
.B1(n_39),
.B2(n_20),
.Y(n_165)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_167),
.Y(n_240)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_169),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_170),
.B(n_184),
.Y(n_227)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_171),
.Y(n_217)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_175),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_44),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_176),
.B(n_183),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_120),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_149),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_186),
.B(n_192),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_109),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_196),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_29),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_212),
.Y(n_236)
);

BUFx4f_ASAP7_75t_SL g189 ( 
.A(n_123),
.Y(n_189)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_127),
.A2(n_46),
.B(n_49),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_98),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_193),
.Y(n_241)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_152),
.B(n_159),
.C(n_162),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_108),
.B(n_100),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_205),
.B1(n_210),
.B2(n_213),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_130),
.A2(n_57),
.B1(n_49),
.B2(n_104),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_198),
.A2(n_199),
.B1(n_202),
.B2(n_204),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_139),
.A2(n_49),
.B1(n_94),
.B2(n_54),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_200),
.B(n_201),
.Y(n_242)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_207),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_139),
.A2(n_62),
.B1(n_65),
.B2(n_75),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_146),
.A2(n_89),
.B1(n_102),
.B2(n_92),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_209),
.Y(n_249)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_118),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_L g211 ( 
.A1(n_106),
.A2(n_85),
.B1(n_84),
.B2(n_90),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_211),
.A2(n_214),
.B1(n_137),
.B2(n_112),
.Y(n_225)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_146),
.A2(n_87),
.B1(n_19),
.B2(n_86),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_181),
.A2(n_213),
.B1(n_165),
.B2(n_132),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_216),
.A2(n_225),
.B1(n_233),
.B2(n_244),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_181),
.A2(n_140),
.B1(n_112),
.B2(n_153),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_176),
.A2(n_107),
.B1(n_119),
.B2(n_153),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_176),
.B(n_107),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_192),
.Y(n_253)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_236),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_268),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_192),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_220),
.A2(n_206),
.B1(n_191),
.B2(n_197),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_255),
.A2(n_257),
.B(n_218),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_235),
.B1(n_234),
.B2(n_229),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_256),
.A2(n_279),
.B1(n_152),
.B2(n_217),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_197),
.B(n_196),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_236),
.B(n_188),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_259),
.B(n_265),
.Y(n_294)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_233),
.A2(n_211),
.B1(n_168),
.B2(n_175),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_263),
.A2(n_224),
.B1(n_218),
.B2(n_240),
.Y(n_285)
);

OAI32xp33_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_178),
.A3(n_195),
.B1(n_201),
.B2(n_212),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_270),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_242),
.B(n_190),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_248),
.A2(n_174),
.B1(n_203),
.B2(n_172),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_266),
.A2(n_267),
.B(n_271),
.C(n_274),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_189),
.B(n_17),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_223),
.B(n_186),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_208),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_247),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_237),
.A2(n_171),
.B1(n_133),
.B2(n_110),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_272),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_273),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g274 ( 
.A1(n_225),
.A2(n_189),
.B(n_99),
.C(n_58),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_180),
.C(n_154),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_280),
.C(n_141),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_216),
.B(n_17),
.Y(n_276)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_276),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_245),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_277),
.A2(n_238),
.B1(n_222),
.B2(n_145),
.Y(n_299)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_278),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_223),
.A2(n_119),
.B1(n_126),
.B2(n_122),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_228),
.B(n_46),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_285),
.A2(n_296),
.B1(n_297),
.B2(n_279),
.Y(n_315)
);

OAI32xp33_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_237),
.A3(n_228),
.B1(n_224),
.B2(n_158),
.Y(n_288)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_288),
.Y(n_324)
);

OAI32xp33_ASAP7_75t_L g290 ( 
.A1(n_256),
.A2(n_241),
.A3(n_226),
.B1(n_221),
.B2(n_147),
.Y(n_290)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_291),
.A2(n_298),
.B(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_128),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_257),
.A2(n_221),
.B1(n_167),
.B2(n_240),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_293),
.A2(n_300),
.B1(n_304),
.B2(n_307),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_262),
.A2(n_263),
.B1(n_255),
.B2(n_253),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_260),
.A2(n_221),
.B1(n_240),
.B2(n_239),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_254),
.A2(n_217),
.B(n_238),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_272),
.B(n_274),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_126),
.B1(n_231),
.B2(n_207),
.Y(n_300)
);

XNOR2x1_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_275),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_252),
.A2(n_231),
.B1(n_202),
.B2(n_226),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_254),
.A2(n_222),
.B(n_243),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_270),
.A2(n_231),
.B1(n_241),
.B2(n_194),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_269),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_326),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_291),
.A2(n_265),
.B(n_267),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_311),
.A2(n_317),
.B(n_319),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_307),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_337),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_318),
.C(n_302),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_277),
.B1(n_267),
.B2(n_251),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_314),
.A2(n_315),
.B1(n_328),
.B2(n_306),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_SL g316 ( 
.A1(n_289),
.A2(n_267),
.B(n_274),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_316),
.A2(n_333),
.B1(n_285),
.B2(n_298),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_268),
.B(n_274),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_280),
.C(n_259),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_287),
.A2(n_258),
.B(n_274),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_321),
.A2(n_289),
.B(n_182),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_283),
.B(n_278),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_322),
.B(n_327),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_282),
.B(n_264),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_325),
.B(n_105),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_261),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_294),
.B(n_243),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_283),
.B(n_309),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_329),
.B(n_35),
.Y(n_359)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_331),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_219),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_336),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_300),
.A2(n_193),
.B1(n_185),
.B2(n_230),
.Y(n_333)
);

INVx13_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_334),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_287),
.A2(n_230),
.B(n_173),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_335),
.A2(n_219),
.B(n_232),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_296),
.B(n_219),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_32),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_339),
.A2(n_352),
.B1(n_360),
.B2(n_319),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_304),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_342),
.Y(n_372)
);

FAx1_ASAP7_75t_SL g345 ( 
.A(n_310),
.B(n_293),
.CI(n_292),
.CON(n_345),
.SN(n_345)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_345),
.B(n_349),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_305),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_346),
.B(n_351),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_290),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_349),
.B(n_350),
.C(n_358),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_299),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_323),
.A2(n_289),
.B1(n_288),
.B2(n_295),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_353),
.A2(n_320),
.B1(n_334),
.B2(n_42),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_308),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_354),
.B(n_367),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_306),
.Y(n_355)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_355),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g356 ( 
.A1(n_330),
.A2(n_289),
.B(n_295),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_356),
.A2(n_357),
.B(n_365),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_179),
.C(n_289),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_359),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_330),
.A2(n_124),
.B1(n_72),
.B2(n_60),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_361),
.B(n_311),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_324),
.A2(n_35),
.B1(n_51),
.B2(n_32),
.Y(n_362)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_232),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_336),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_331),
.B(n_51),
.Y(n_367)
);

BUFx5_ASAP7_75t_L g368 ( 
.A(n_364),
.Y(n_368)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_368),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_369),
.A2(n_379),
.B1(n_366),
.B2(n_346),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_324),
.Y(n_370)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_375),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_338),
.Y(n_373)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g413 ( 
.A(n_376),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_321),
.Y(n_378)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_352),
.A2(n_315),
.B1(n_312),
.B2(n_317),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_347),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_387),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_391),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_341),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_348),
.A2(n_335),
.B(n_328),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_388),
.B(n_232),
.Y(n_405)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_363),
.Y(n_389)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_389),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_334),
.Y(n_390)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_390),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_339),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_323),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_392),
.B(n_393),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_356),
.B(n_333),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_394),
.A2(n_358),
.B1(n_357),
.B2(n_356),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_369),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_391),
.A2(n_348),
.B(n_345),
.Y(n_397)
);

NAND3xp33_ASAP7_75t_SL g435 ( 
.A(n_397),
.B(n_381),
.C(n_390),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_383),
.A2(n_345),
.B1(n_350),
.B2(n_351),
.Y(n_399)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_399),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_400),
.A2(n_415),
.B1(n_376),
.B2(n_388),
.Y(n_421)
);

XNOR2x1_ASAP7_75t_SL g401 ( 
.A(n_386),
.B(n_361),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_405),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_343),
.C(n_340),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_414),
.C(n_375),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_391),
.A2(n_320),
.B1(n_343),
.B2(n_340),
.Y(n_404)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_380),
.A2(n_42),
.B1(n_91),
.B2(n_11),
.Y(n_412)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_412),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_386),
.C(n_384),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_379),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_395),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_419),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_411),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_421),
.B(n_423),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_386),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_401),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_395),
.Y(n_426)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_426),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_368),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_431),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_428),
.A2(n_433),
.B1(n_403),
.B2(n_406),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_372),
.C(n_378),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_429),
.B(n_404),
.C(n_416),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_403),
.A2(n_393),
.B1(n_370),
.B2(n_392),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_430),
.A2(n_432),
.B1(n_434),
.B2(n_409),
.Y(n_442)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_385),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_408),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_410),
.Y(n_434)
);

XOR2x1_ASAP7_75t_SL g447 ( 
.A(n_435),
.B(n_397),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_418),
.A2(n_410),
.B(n_414),
.Y(n_437)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_437),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_443),
.Y(n_465)
);

OAI321xp33_ASAP7_75t_L g439 ( 
.A1(n_427),
.A2(n_373),
.A3(n_377),
.B1(n_368),
.B2(n_409),
.C(n_380),
.Y(n_439)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_439),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_416),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_436),
.Y(n_453)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_442),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_425),
.C(n_422),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_444),
.B(n_448),
.C(n_434),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_424),
.A2(n_382),
.B1(n_407),
.B2(n_406),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_445),
.B(n_449),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_421),
.A2(n_396),
.B1(n_407),
.B2(n_405),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_446),
.A2(n_430),
.B1(n_433),
.B2(n_382),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_447),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_377),
.C(n_371),
.Y(n_448)
);

OAI321xp33_ASAP7_75t_L g449 ( 
.A1(n_419),
.A2(n_370),
.A3(n_385),
.B1(n_381),
.B2(n_394),
.C(n_415),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_420),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_453),
.B(n_457),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_447),
.B(n_387),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_460),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_420),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_462),
.A2(n_464),
.B(n_440),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_463),
.A2(n_455),
.B1(n_456),
.B2(n_446),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_444),
.A2(n_433),
.B(n_389),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_450),
.A2(n_166),
.B(n_99),
.Y(n_466)
);

O2A1O1Ixp33_ASAP7_75t_L g477 ( 
.A1(n_466),
.A2(n_21),
.B(n_12),
.C(n_11),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_451),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_0),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_471),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_465),
.B(n_438),
.C(n_448),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_469),
.B(n_470),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_454),
.Y(n_471)
);

AOI221xp5_ASAP7_75t_L g472 ( 
.A1(n_459),
.A2(n_452),
.B1(n_443),
.B2(n_441),
.C(n_74),
.Y(n_472)
);

NOR2x1_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_478),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_461),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_475),
.B(n_476),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_21),
.C(n_13),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_477),
.B(n_479),
.Y(n_481)
);

AND2x2_ASAP7_75t_SL g478 ( 
.A(n_461),
.B(n_0),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_478),
.A2(n_466),
.B1(n_467),
.B2(n_463),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_474),
.B(n_453),
.C(n_460),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_480),
.B(n_484),
.C(n_21),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_482),
.B(n_3),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_483),
.A2(n_0),
.B(n_2),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_21),
.C(n_2),
.Y(n_484)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_487),
.B(n_473),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_491),
.C(n_485),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_489),
.B(n_490),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_486),
.A2(n_5),
.B(n_6),
.Y(n_492)
);

AOI21xp33_ASAP7_75t_L g493 ( 
.A1(n_492),
.A2(n_481),
.B(n_482),
.Y(n_493)
);

NAND4xp25_ASAP7_75t_L g496 ( 
.A(n_493),
.B(n_494),
.C(n_5),
.D(n_6),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_496),
.A2(n_497),
.B(n_5),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_495),
.B(n_21),
.C(n_6),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_498),
.B(n_9),
.C(n_5),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_7),
.C(n_9),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_7),
.B(n_9),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_7),
.B(n_450),
.Y(n_502)
);


endmodule