module real_jpeg_19633_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_335, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_335;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_323;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_1),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_1),
.A2(n_26),
.B1(n_32),
.B2(n_50),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_2),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_130),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_130),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_2),
.A2(n_26),
.B1(n_32),
.B2(n_130),
.Y(n_267)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_3),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_28),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_3),
.A2(n_8),
.B(n_63),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_133),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_3),
.A2(n_105),
.B1(n_112),
.B2(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_3),
.B(n_87),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_3),
.B(n_30),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_3),
.A2(n_30),
.B(n_219),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_4),
.A2(n_26),
.B1(n_32),
.B2(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_4),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_57),
.Y(n_117)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_6),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_6),
.A2(n_26),
.B1(n_32),
.B2(n_128),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_128),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_128),
.Y(n_208)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_7),
.Y(n_108)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_8),
.A2(n_45),
.B(n_60),
.C(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_8),
.B(n_45),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_10),
.A2(n_26),
.B1(n_32),
.B2(n_135),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_10),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_135),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_135),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_135),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_12),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_12),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_12),
.A2(n_33),
.B1(n_62),
.B2(n_63),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_283)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_14),
.A2(n_26),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_14),
.A2(n_35),
.B1(n_62),
.B2(n_63),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_14),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_259)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_15),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_78),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_73),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_20),
.A2(n_21),
.B1(n_70),
.B2(n_321),
.Y(n_327)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_37),
.B1(n_38),
.B2(n_69),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_23),
.A2(n_36),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_23),
.A2(n_36),
.B1(n_147),
.B2(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_23),
.A2(n_267),
.B(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_23),
.A2(n_84),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_24),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_24),
.A2(n_28),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_26),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_25),
.B(n_30),
.Y(n_139)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g132 ( 
.A(n_26),
.B(n_133),
.CON(n_132),
.SN(n_132)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_27),
.A2(n_29),
.B1(n_132),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_28),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_28),
.B(n_287),
.Y(n_286)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g218 ( 
.A1(n_29),
.A2(n_45),
.A3(n_48),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_42),
.B(n_43),
.C(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_43),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_31),
.A2(n_36),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_51),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_41),
.A2(n_52),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_49),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_42),
.A2(n_53),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_42),
.A2(n_53),
.B1(n_166),
.B2(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_42),
.A2(n_51),
.B(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_42),
.A2(n_53),
.B1(n_76),
.B2(n_283),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_42)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g220 ( 
.A(n_43),
.B(n_46),
.Y(n_220)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_46),
.A2(n_64),
.B(n_133),
.C(n_184),
.Y(n_183)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_75),
.B(n_77),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_52),
.A2(n_87),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_52),
.A2(n_77),
.B(n_88),
.Y(n_269)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_68),
.C(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_58),
.A2(n_67),
.B1(n_74),
.B2(n_324),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_61),
.B(n_65),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_59),
.A2(n_65),
.B(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_59),
.A2(n_61),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_59),
.A2(n_61),
.B1(n_188),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_59),
.A2(n_61),
.B1(n_208),
.B2(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_59),
.A2(n_226),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_59),
.A2(n_61),
.B1(n_115),
.B2(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_59),
.A2(n_123),
.B(n_259),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_61),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_61),
.B(n_133),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_62),
.B(n_197),
.Y(n_196)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_66),
.B(n_124),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_70),
.C(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_70),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_70),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_73),
.B(n_327),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_74),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_318),
.A3(n_328),
.B1(n_331),
.B2(n_332),
.C(n_335),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_298),
.B(n_317),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_274),
.B(n_297),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_168),
.B(n_250),
.C(n_273),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_152),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_99),
.B(n_152),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_136),
.B2(n_151),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_120),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_102),
.B(n_120),
.C(n_151),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_114),
.B2(n_119),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_103),
.B(n_119),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B(n_110),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_105),
.A2(n_109),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_105),
.A2(n_108),
.B1(n_177),
.B2(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_105),
.A2(n_180),
.B(n_210),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_105),
.A2(n_108),
.B(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_106),
.B(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_106),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_106),
.A2(n_111),
.B(n_211),
.Y(n_217)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_107),
.B(n_211),
.Y(n_210)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_141),
.B(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_112),
.B(n_133),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_116),
.B(n_242),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.C(n_131),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_127),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_137),
.B(n_144),
.C(n_149),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_140),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_157),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_153),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.C(n_164),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_161),
.B(n_210),
.Y(n_257)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_163),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_164),
.B(n_236),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_249),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_244),
.B(n_248),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_231),
.B(n_243),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_213),
.B(n_230),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_200),
.B(n_212),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_189),
.B(n_199),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_181),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_181),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_183),
.B(n_185),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_194),
.B(n_198),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_192),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_202),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_209),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_207),
.C(n_209),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_211),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_215),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_221),
.B1(n_228),
.B2(n_229),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_222),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_227),
.C(n_228),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_233),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_238),
.B2(n_239),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_240),
.C(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_252),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_271),
.B2(n_272),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_260),
.B2(n_261),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_261),
.C(n_272),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_270),
.Y(n_261)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_269),
.C(n_270),
.Y(n_296)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_275),
.B(n_276),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_296),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_289),
.B2(n_290),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_290),
.C(n_296),
.Y(n_299)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_284),
.C(n_288),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_284),
.B1(n_285),
.B2(n_288),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_282),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_287),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_292),
.B1(n_312),
.B2(n_314),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_291),
.A2(n_308),
.B(n_312),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_294),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_300),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_315),
.B2(n_316),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_307),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_307),
.C(n_316),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_305),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_320),
.C(n_325),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g330 ( 
.A(n_306),
.B(n_320),
.CI(n_325),
.CON(n_330),
.SN(n_330)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_312),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_315),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_326),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_326),
.Y(n_332)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_330),
.Y(n_334)
);


endmodule