module fake_jpeg_31087_n_167 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_39),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_14),
.B1(n_15),
.B2(n_25),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_45),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_38),
.B1(n_25),
.B2(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_62),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_51),
.A2(n_27),
.B1(n_30),
.B2(n_29),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_28),
.Y(n_59)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_21),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_63),
.Y(n_100)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_27),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_69),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_26),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_16),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_80),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_16),
.B(n_34),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_31),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_80),
.B1(n_57),
.B2(n_62),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_97),
.B1(n_90),
.B2(n_86),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_17),
.B1(n_22),
.B2(n_34),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_37),
.B1(n_78),
.B2(n_17),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_22),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_95),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_34),
.B(n_37),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_77),
.C(n_70),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_13),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_9),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_9),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_1),
.B(n_2),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_107),
.Y(n_121)
);

XNOR2x1_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_69),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_64),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_106),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_58),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_79),
.C(n_60),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_60),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_114),
.B(n_105),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_116),
.B1(n_100),
.B2(n_83),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_115),
.B(n_89),
.C(n_81),
.D(n_117),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_55),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_97),
.B(n_86),
.C(n_93),
.D(n_88),
.Y(n_124)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_109),
.C(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_95),
.B1(n_83),
.B2(n_85),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_116),
.B1(n_110),
.B2(n_100),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_114),
.B1(n_101),
.B2(n_108),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_119),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_140),
.B(n_120),
.Y(n_142)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_84),
.B(n_61),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_144),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_130),
.C(n_127),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_147),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_128),
.B1(n_123),
.B2(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_146),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_124),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_122),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_136),
.B(n_137),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_151),
.B(n_152),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_138),
.B(n_84),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_55),
.B(n_37),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_147),
.B1(n_141),
.B2(n_148),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_158),
.C(n_3),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_2),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_150),
.B(n_63),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_156),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_162),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_165)
);

OAI21x1_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_3),
.B(n_4),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_4),
.Y(n_167)
);


endmodule