module fake_netlist_1_6578_n_43 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_43);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_43;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_30;
wire n_16;
wire n_26;
wire n_25;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
NAND2xp33_ASAP7_75t_L g14 ( .A(n_5), .B(n_4), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_1), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_9), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_10), .B(n_13), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_3), .Y(n_21) );
AND2x4_ASAP7_75t_L g22 ( .A(n_15), .B(n_0), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_21), .B(n_1), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_18), .B(n_2), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_17), .Y(n_25) );
BUFx3_ASAP7_75t_L g26 ( .A(n_22), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_22), .Y(n_27) );
INVx2_ASAP7_75t_SL g28 ( .A(n_26), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_27), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_16), .Y(n_31) );
O2A1O1Ixp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_23), .B(n_25), .C(n_24), .Y(n_32) );
INVx2_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
AOI21xp33_ASAP7_75t_SL g34 ( .A1(n_33), .A2(n_20), .B(n_19), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
NAND5xp2_ASAP7_75t_L g37 ( .A(n_35), .B(n_14), .C(n_7), .D(n_8), .E(n_12), .Y(n_37) );
INVx3_ASAP7_75t_SL g38 ( .A(n_36), .Y(n_38) );
CKINVDCx5p33_ASAP7_75t_R g39 ( .A(n_34), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
INVx1_ASAP7_75t_L g41 ( .A(n_38), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_40), .Y(n_42) );
AOI22x1_ASAP7_75t_L g43 ( .A1(n_42), .A2(n_39), .B1(n_41), .B2(n_37), .Y(n_43) );
endmodule