module fake_jpeg_19250_n_284 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_38),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_20),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_61),
.C(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_56),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_56),
.Y(n_73)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

CKINVDCx10_ASAP7_75t_R g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_30),
.B1(n_28),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_54),
.B1(n_58),
.B2(n_63),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_64),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_30),
.B1(n_28),
.B2(n_21),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_27),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_28),
.B1(n_21),
.B2(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_22),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_20),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_37),
.B1(n_38),
.B2(n_17),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_76),
.B1(n_58),
.B2(n_41),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_38),
.B1(n_18),
.B2(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_43),
.A2(n_15),
.B1(n_23),
.B2(n_22),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_33),
.C(n_45),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_92),
.B(n_108),
.Y(n_132)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_46),
.B(n_60),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_100),
.B(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_111),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_42),
.B1(n_44),
.B2(n_61),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_100),
.B1(n_97),
.B2(n_96),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_65),
.B(n_61),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_71),
.B(n_69),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_42),
.B(n_57),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_64),
.C(n_86),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_62),
.B1(n_55),
.B2(n_59),
.Y(n_105)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_109),
.B(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_62),
.B1(n_43),
.B2(n_45),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_49),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_15),
.B(n_23),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_126),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_82),
.B1(n_73),
.B2(n_57),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_122),
.Y(n_156)
);

NAND2x1p5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_73),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_125),
.B(n_109),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_106),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_127),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_113),
.B1(n_92),
.B2(n_89),
.Y(n_119)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_43),
.B1(n_80),
.B2(n_68),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_74),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_103),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_89),
.A2(n_68),
.B1(n_87),
.B2(n_79),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_102),
.B1(n_91),
.B2(n_94),
.Y(n_128)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_69),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_134),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_77),
.B1(n_86),
.B2(n_55),
.Y(n_130)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_31),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_109),
.C(n_90),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_29),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_138),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_143),
.C(n_146),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_144),
.B(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_11),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_141),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_109),
.C(n_104),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_90),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_48),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_64),
.C(n_48),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_152),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_29),
.C(n_22),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_159),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_120),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_162),
.A2(n_159),
.B(n_152),
.Y(n_180)
);

OAI22x1_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_119),
.B1(n_118),
.B2(n_135),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_135),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_177),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_R g172 ( 
.A1(n_144),
.A2(n_118),
.B(n_123),
.C(n_134),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_175),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_160),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_174),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_129),
.B(n_125),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_178),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_143),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_151),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_180),
.B(n_162),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_136),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_181),
.B(n_182),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_123),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_153),
.A2(n_140),
.B1(n_158),
.B2(n_147),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_185),
.B1(n_186),
.B2(n_0),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_153),
.A2(n_118),
.B1(n_130),
.B2(n_117),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_125),
.B1(n_121),
.B2(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_149),
.B1(n_154),
.B2(n_141),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_188),
.A2(n_190),
.B1(n_191),
.B2(n_185),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_164),
.A2(n_154),
.B1(n_155),
.B2(n_148),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_175),
.A2(n_157),
.B1(n_131),
.B2(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_31),
.C(n_22),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_199),
.C(n_169),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_168),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_204),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_29),
.C(n_7),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_200),
.A2(n_171),
.B1(n_169),
.B2(n_174),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_166),
.Y(n_215)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_14),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_165),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_7),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_13),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_215),
.B1(n_191),
.B2(n_189),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_209),
.A2(n_211),
.B1(n_221),
.B2(n_200),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_183),
.B1(n_186),
.B2(n_167),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_220),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_179),
.C(n_166),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_199),
.C(n_197),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_6),
.B1(n_12),
.B2(n_10),
.Y(n_221)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_223),
.B(n_192),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_6),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_224),
.B(n_225),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_204),
.B(n_8),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_195),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_233),
.C(n_234),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

NAND2x1_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_212),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_195),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_236),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_198),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_238),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_206),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_221),
.B1(n_220),
.B2(n_13),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_222),
.B(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_226),
.A2(n_209),
.B(n_208),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_3),
.B(n_4),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_234),
.A2(n_213),
.B1(n_223),
.B2(n_215),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_227),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_250),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_9),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_252),
.B(n_1),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_256),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_228),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_257),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_233),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_238),
.B(n_228),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_249),
.B(n_245),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_237),
.C(n_4),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_251),
.C(n_250),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_263),
.B(n_266),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_241),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_269),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_4),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_256),
.C(n_254),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_274),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_258),
.C(n_4),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_258),
.Y(n_275)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_265),
.B(n_5),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_276),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_272),
.B(n_5),
.CI(n_271),
.CON(n_277),
.SN(n_277)
);

O2A1O1Ixp33_ASAP7_75t_SL g281 ( 
.A1(n_277),
.A2(n_5),
.B(n_278),
.C(n_279),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_277),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_282),
.B(n_280),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_283),
.Y(n_284)
);


endmodule