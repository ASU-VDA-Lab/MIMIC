module fake_jpeg_24128_n_267 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_1),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_39),
.B(n_2),
.Y(n_89)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_41),
.B(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_60),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_55),
.A2(n_84),
.B1(n_28),
.B2(n_22),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_67),
.B1(n_71),
.B2(n_80),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_61),
.Y(n_92)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_27),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_65),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_25),
.B(n_24),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_63),
.A2(n_30),
.B(n_29),
.C(n_28),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_17),
.B1(n_23),
.B2(n_26),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_48),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_17),
.B1(n_23),
.B2(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_38),
.Y(n_72)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_87),
.Y(n_95)
);

CKINVDCx12_ASAP7_75t_R g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_79),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_42),
.A2(n_36),
.B1(n_19),
.B2(n_32),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_83),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g84 ( 
.A1(n_37),
.A2(n_33),
.B1(n_3),
.B2(n_4),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_32),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_77),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_33),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_117),
.Y(n_120)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_111),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_33),
.B1(n_4),
.B2(n_5),
.Y(n_110)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_118),
.B(n_22),
.Y(n_124)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_119),
.B1(n_20),
.B2(n_52),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_20),
.B1(n_72),
.B2(n_53),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_3),
.Y(n_117)
);

AO22x1_ASAP7_75t_L g118 ( 
.A1(n_55),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_122),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_71),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_123),
.B(n_130),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_127),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_86),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_128),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_76),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_135),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_69),
.CI(n_81),
.CON(n_130),
.SN(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_52),
.B1(n_58),
.B2(n_88),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_134),
.B1(n_143),
.B2(n_101),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_133),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_82),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_137),
.Y(n_159)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_141),
.B1(n_144),
.B2(n_146),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_147),
.B(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_50),
.Y(n_140)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_78),
.B1(n_62),
.B2(n_73),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_148),
.B1(n_107),
.B2(n_109),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_73),
.B1(n_64),
.B2(n_54),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_82),
.B(n_7),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_99),
.B(n_104),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_92),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_64),
.B(n_54),
.C(n_66),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_118),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_148)
);

AOI32xp33_ASAP7_75t_L g149 ( 
.A1(n_96),
.A2(n_6),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_154),
.A2(n_163),
.B1(n_171),
.B2(n_173),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_156),
.A2(n_176),
.B(n_138),
.Y(n_195)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_158),
.B(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_136),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_168),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_104),
.C(n_95),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_101),
.B1(n_107),
.B2(n_111),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_175),
.B1(n_109),
.B2(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_178),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_120),
.A2(n_107),
.B1(n_94),
.B2(n_102),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_96),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_132),
.A2(n_97),
.B(n_94),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_187),
.Y(n_201)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_130),
.B(n_124),
.C(n_149),
.D(n_122),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_170),
.C(n_165),
.Y(n_209)
);

NAND2xp33_ASAP7_75t_SL g182 ( 
.A(n_176),
.B(n_178),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_182),
.A2(n_152),
.B(n_168),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_121),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_194),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_196),
.B1(n_158),
.B2(n_154),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_124),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_192),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_146),
.B1(n_150),
.B2(n_148),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_163),
.B1(n_172),
.B2(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_195),
.A2(n_156),
.B(n_164),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_90),
.B1(n_91),
.B2(n_135),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_129),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_197),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_198),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_166),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_209),
.C(n_215),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_184),
.A2(n_173),
.B1(n_171),
.B2(n_166),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_204),
.A2(n_208),
.B1(n_213),
.B2(n_190),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_207),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_174),
.B1(n_151),
.B2(n_164),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_210),
.A2(n_192),
.B1(n_183),
.B2(n_180),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_184),
.A2(n_165),
.B1(n_169),
.B2(n_177),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_182),
.B(n_180),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_189),
.C(n_197),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_152),
.C(n_127),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_222),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_221),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_206),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_219),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_199),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_196),
.B1(n_199),
.B2(n_191),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_226),
.B(n_228),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_179),
.B1(n_181),
.B2(n_187),
.Y(n_226)
);

BUFx12_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_230),
.B(n_215),
.Y(n_235)
);

AOI31xp67_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_214),
.A3(n_200),
.B(n_202),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_205),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_227),
.A2(n_207),
.B(n_200),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_238),
.B(n_208),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_228),
.Y(n_249)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_204),
.B(n_210),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_241),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_203),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_240),
.A2(n_229),
.B1(n_218),
.B2(n_221),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_234),
.B(n_232),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_240),
.A2(n_224),
.B1(n_226),
.B2(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_246),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_217),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_249),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_238),
.B(n_228),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_228),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_242),
.C(n_220),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_233),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_253),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_255),
.A2(n_245),
.B(n_244),
.Y(n_257)
);

OAI21x1_ASAP7_75t_SL g258 ( 
.A1(n_256),
.A2(n_243),
.B(n_241),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_257),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_258),
.A2(n_254),
.B1(n_137),
.B2(n_141),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_90),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_259),
.B(n_11),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_262),
.A3(n_260),
.B1(n_259),
.B2(n_16),
.C1(n_15),
.C2(n_14),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_12),
.C(n_13),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_265),
.Y(n_267)
);


endmodule