module fake_netlist_6_1460_n_951 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_951);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_951;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_842;
wire n_720;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_63),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_183),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_85),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_36),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_149),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_175),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_38),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_89),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_30),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_133),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_10),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_28),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_47),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_156),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_119),
.Y(n_203)
);

BUFx2_ASAP7_75t_SL g204 ( 
.A(n_158),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_74),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_152),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_46),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_75),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_26),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_19),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_2),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_59),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_138),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_157),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_102),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_132),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_49),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_9),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_21),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_55),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_65),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_18),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_66),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_58),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_82),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_146),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_166),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_141),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_136),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_43),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_126),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_45),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_129),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_180),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_53),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_94),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_16),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_31),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_12),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_177),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_105),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_34),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_125),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_100),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_137),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_135),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_16),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_76),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_32),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_99),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_174),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_22),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_116),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_140),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_72),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_14),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_122),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_91),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_187),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_211),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_220),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_259),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_186),
.B(n_0),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_203),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_194),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_189),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_195),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_236),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_188),
.B(n_0),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_199),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_201),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_208),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_219),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_253),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_190),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_191),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_260),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_233),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_238),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_207),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_192),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_245),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_193),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_196),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_249),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_252),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_207),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_188),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_197),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_198),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_213),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_224),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_207),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_207),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_202),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_263),
.B(n_185),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_312),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_307),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_296),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_296),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_185),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_200),
.Y(n_323)
);

AND3x1_ASAP7_75t_L g324 ( 
.A(n_268),
.B(n_250),
.C(n_237),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_216),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_265),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

OAI21x1_ASAP7_75t_L g329 ( 
.A1(n_306),
.A2(n_204),
.B(n_231),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_287),
.B(n_206),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_276),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_266),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_269),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_280),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g339 ( 
.A(n_283),
.B(n_209),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_270),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_285),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_262),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_295),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_301),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_302),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_271),
.B(n_209),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_264),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_309),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_272),
.B(n_261),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_297),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_299),
.B(n_209),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_278),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_310),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_310),
.B(n_237),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_273),
.B(n_237),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_277),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_290),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_291),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_284),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_284),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_286),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_328),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_341),
.B(n_210),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_361),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_343),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

BUFx4f_ASAP7_75t_L g376 ( 
.A(n_361),
.Y(n_376)
);

INVx8_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_325),
.B(n_286),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_345),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_318),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_354),
.B(n_212),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_325),
.B(n_323),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_361),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_214),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_215),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_348),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_217),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_317),
.B(n_218),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_318),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_357),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_354),
.B(n_222),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_357),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_325),
.B(n_223),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_350),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_321),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_319),
.B(n_320),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_321),
.Y(n_403)
);

AND2x6_ASAP7_75t_L g404 ( 
.A(n_358),
.B(n_27),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_321),
.Y(n_405)
);

OR2x6_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_267),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g407 ( 
.A(n_358),
.B(n_29),
.Y(n_407)
);

AND3x4_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_282),
.C(n_267),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_326),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_352),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_352),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_325),
.B(n_225),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_327),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_361),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_337),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_323),
.B(n_226),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_323),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_319),
.B(n_227),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_337),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_327),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_320),
.B(n_229),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_339),
.A2(n_243),
.B1(n_257),
.B2(n_256),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_323),
.B(n_230),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g425 ( 
.A(n_331),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_351),
.B(n_234),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_337),
.Y(n_427)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_354),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_316),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_337),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_337),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_358),
.B(n_235),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_355),
.Y(n_434)
);

AO22x2_ASAP7_75t_L g435 ( 
.A1(n_363),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g436 ( 
.A(n_356),
.B(n_33),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_364),
.B(n_239),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_369),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_335),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_354),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_316),
.Y(n_441)
);

NAND3x1_ASAP7_75t_L g442 ( 
.A(n_364),
.B(n_282),
.C(n_3),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_324),
.A2(n_248),
.B1(n_247),
.B2(n_246),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_355),
.Y(n_444)
);

NAND2x1p5_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_355),
.Y(n_445)
);

AO22x2_ASAP7_75t_L g446 ( 
.A1(n_408),
.A2(n_362),
.B1(n_368),
.B2(n_370),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_355),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_371),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_383),
.B(n_356),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_412),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_360),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_371),
.B(n_342),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_375),
.Y(n_455)
);

AO22x2_ASAP7_75t_L g456 ( 
.A1(n_383),
.A2(n_362),
.B1(n_368),
.B2(n_370),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_360),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_380),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_387),
.Y(n_460)
);

OR2x2_ASAP7_75t_SL g461 ( 
.A(n_442),
.B(n_367),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_393),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_428),
.A2(n_339),
.B1(n_314),
.B2(n_322),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_398),
.B(n_332),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_409),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_394),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_410),
.Y(n_467)
);

AO22x2_ASAP7_75t_L g468 ( 
.A1(n_378),
.A2(n_365),
.B1(n_324),
.B2(n_359),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_438),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_406),
.Y(n_470)
);

AO22x2_ASAP7_75t_L g471 ( 
.A1(n_435),
.A2(n_365),
.B1(n_359),
.B2(n_340),
.Y(n_471)
);

AO22x2_ASAP7_75t_L g472 ( 
.A1(n_435),
.A2(n_336),
.B1(n_340),
.B2(n_5),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_381),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_414),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_421),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_424),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_372),
.B(n_339),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_429),
.Y(n_479)
);

AO22x2_ASAP7_75t_L g480 ( 
.A1(n_435),
.A2(n_336),
.B1(n_4),
.B2(n_5),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_428),
.Y(n_481)
);

AO22x2_ASAP7_75t_L g482 ( 
.A1(n_392),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_384),
.B(n_330),
.Y(n_483)
);

NAND2x1p5_ASAP7_75t_L g484 ( 
.A(n_415),
.B(n_329),
.Y(n_484)
);

NAND2x1p5_ASAP7_75t_L g485 ( 
.A(n_388),
.B(n_329),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_390),
.B(n_353),
.Y(n_486)
);

NAND2x1p5_ASAP7_75t_L g487 ( 
.A(n_388),
.B(n_330),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_439),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_372),
.B(n_339),
.Y(n_489)
);

BUFx6f_ASAP7_75t_SL g490 ( 
.A(n_406),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_381),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

AO22x2_ASAP7_75t_L g494 ( 
.A1(n_413),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_391),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_391),
.Y(n_496)
);

AO22x2_ASAP7_75t_L g497 ( 
.A1(n_417),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_497)
);

AO22x2_ASAP7_75t_L g498 ( 
.A1(n_382),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

AO22x2_ASAP7_75t_L g500 ( 
.A1(n_382),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_500)
);

AO22x2_ASAP7_75t_L g501 ( 
.A1(n_396),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_SL g502 ( 
.A(n_426),
.B(n_241),
.Y(n_502)
);

AO22x2_ASAP7_75t_L g503 ( 
.A1(n_396),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_395),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_403),
.Y(n_506)
);

OR2x2_ASAP7_75t_SL g507 ( 
.A(n_437),
.B(n_349),
.Y(n_507)
);

NAND2x1p5_ASAP7_75t_L g508 ( 
.A(n_399),
.B(n_349),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_403),
.Y(n_509)
);

OAI22xp33_ASAP7_75t_SL g510 ( 
.A1(n_437),
.A2(n_251),
.B1(n_344),
.B2(n_333),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_405),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_428),
.A2(n_339),
.B1(n_346),
.B2(n_344),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_390),
.B(n_333),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_385),
.B(n_339),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_430),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_385),
.A2(n_346),
.B1(n_338),
.B2(n_334),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_441),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_443),
.B(n_334),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_376),
.B(n_338),
.Y(n_520)
);

AO22x2_ASAP7_75t_L g521 ( 
.A1(n_443),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_406),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_401),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_425),
.B(n_337),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_386),
.A2(n_389),
.B1(n_423),
.B2(n_376),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_454),
.B(n_373),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_444),
.B(n_373),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_464),
.B(n_423),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_SL g529 ( 
.A(n_477),
.B(n_386),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_514),
.B(n_389),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_447),
.B(n_422),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_SL g532 ( 
.A(n_469),
.B(n_422),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_449),
.B(n_419),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_458),
.B(n_419),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_510),
.B(n_377),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_SL g536 ( 
.A(n_493),
.B(n_490),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_492),
.B(n_404),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_486),
.B(n_377),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_448),
.B(n_315),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_499),
.B(n_404),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_524),
.B(n_377),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_445),
.B(n_401),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_450),
.B(n_404),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_451),
.B(n_436),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_525),
.B(n_416),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_SL g546 ( 
.A(n_453),
.B(n_416),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_455),
.B(n_404),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_457),
.B(n_416),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_459),
.B(n_420),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_460),
.B(n_436),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_463),
.B(n_420),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_462),
.B(n_420),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_SL g553 ( 
.A(n_466),
.B(n_431),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_470),
.B(n_35),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_SL g555 ( 
.A(n_473),
.B(n_431),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_SL g556 ( 
.A(n_475),
.B(n_431),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_476),
.B(n_407),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_479),
.B(n_432),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_488),
.B(n_407),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_481),
.B(n_517),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_502),
.B(n_432),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_SL g562 ( 
.A(n_478),
.B(n_489),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_495),
.B(n_407),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_474),
.B(n_491),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_496),
.B(n_432),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_504),
.B(n_427),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_512),
.B(n_427),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_456),
.B(n_407),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_SL g569 ( 
.A(n_515),
.B(n_436),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_523),
.B(n_347),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_452),
.B(n_436),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_513),
.B(n_347),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_456),
.B(n_347),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_505),
.B(n_506),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_509),
.B(n_347),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_511),
.B(n_347),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_487),
.B(n_347),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_452),
.B(n_316),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_508),
.B(n_316),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_452),
.B(n_519),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_SL g581 ( 
.A(n_520),
.B(n_20),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_465),
.B(n_37),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_467),
.B(n_39),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_516),
.B(n_40),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_519),
.B(n_22),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_519),
.B(n_41),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_483),
.B(n_23),
.Y(n_587)
);

AOI211x1_ASAP7_75t_L g588 ( 
.A1(n_528),
.A2(n_480),
.B(n_472),
.C(n_494),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_545),
.A2(n_484),
.B(n_485),
.Y(n_589)
);

NAND3xp33_ASAP7_75t_L g590 ( 
.A(n_529),
.B(n_522),
.C(n_518),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_526),
.B(n_471),
.Y(n_591)
);

AO22x2_ASAP7_75t_L g592 ( 
.A1(n_585),
.A2(n_472),
.B1(n_480),
.B2(n_471),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_562),
.A2(n_483),
.B(n_507),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_537),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_530),
.B(n_483),
.Y(n_595)
);

OAI21x1_ASAP7_75t_L g596 ( 
.A1(n_551),
.A2(n_468),
.B(n_109),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_586),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_531),
.B(n_468),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_540),
.A2(n_497),
.B(n_494),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_534),
.B(n_446),
.Y(n_600)
);

OA21x2_ASAP7_75t_L g601 ( 
.A1(n_551),
.A2(n_497),
.B(n_521),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_586),
.B(n_580),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_539),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_544),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_533),
.A2(n_446),
.B(n_521),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_569),
.A2(n_503),
.B(n_501),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_532),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_573),
.B(n_498),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_559),
.B(n_498),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_544),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_564),
.Y(n_611)
);

AO31x2_ASAP7_75t_L g612 ( 
.A1(n_543),
.A2(n_503),
.A3(n_501),
.B(n_500),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_541),
.A2(n_500),
.B(n_482),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_550),
.B(n_574),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_563),
.A2(n_482),
.B(n_106),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_554),
.B(n_461),
.Y(n_616)
);

AO31x2_ASAP7_75t_L g617 ( 
.A1(n_547),
.A2(n_23),
.A3(n_24),
.B(n_25),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_538),
.A2(n_104),
.B(n_182),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_557),
.A2(n_24),
.B(n_25),
.C(n_42),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_560),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_578),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_568),
.B(n_550),
.Y(n_622)
);

OA21x2_ASAP7_75t_L g623 ( 
.A1(n_527),
.A2(n_572),
.B(n_575),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_571),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_624)
);

OAI21x1_ASAP7_75t_L g625 ( 
.A1(n_570),
.A2(n_566),
.B(n_567),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_587),
.Y(n_626)
);

INVxp33_ASAP7_75t_L g627 ( 
.A(n_561),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_527),
.B(n_184),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_576),
.A2(n_51),
.B(n_52),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_542),
.B(n_54),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_536),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_535),
.A2(n_56),
.B(n_57),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_577),
.A2(n_60),
.B(n_61),
.Y(n_633)
);

AOI21xp33_ASAP7_75t_L g634 ( 
.A1(n_548),
.A2(n_62),
.B(n_64),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_579),
.A2(n_67),
.B(n_68),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_565),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_549),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_581),
.B(n_69),
.Y(n_638)
);

AOI211x1_ASAP7_75t_L g639 ( 
.A1(n_584),
.A2(n_70),
.B(n_71),
.C(n_73),
.Y(n_639)
);

NAND2x1p5_ASAP7_75t_L g640 ( 
.A(n_597),
.B(n_552),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_631),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_603),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_611),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_589),
.A2(n_558),
.B(n_582),
.Y(n_644)
);

AO21x2_ASAP7_75t_L g645 ( 
.A1(n_593),
.A2(n_583),
.B(n_556),
.Y(n_645)
);

BUFx8_ASAP7_75t_L g646 ( 
.A(n_597),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_625),
.A2(n_555),
.B(n_553),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_626),
.Y(n_648)
);

A2O1A1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_638),
.A2(n_546),
.B(n_78),
.C(n_79),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_622),
.Y(n_650)
);

OAI21x1_ASAP7_75t_L g651 ( 
.A1(n_596),
.A2(n_77),
.B(n_80),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_620),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_597),
.Y(n_653)
);

AO21x2_ASAP7_75t_L g654 ( 
.A1(n_632),
.A2(n_81),
.B(n_83),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_636),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_591),
.B(n_84),
.Y(n_656)
);

OA21x2_ASAP7_75t_L g657 ( 
.A1(n_599),
.A2(n_86),
.B(n_87),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_629),
.A2(n_88),
.B(n_90),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_607),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_602),
.B(n_92),
.Y(n_660)
);

OAI22xp33_ASAP7_75t_L g661 ( 
.A1(n_608),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_610),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_600),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_618),
.A2(n_97),
.B(n_98),
.Y(n_664)
);

AOI21xp33_ASAP7_75t_L g665 ( 
.A1(n_598),
.A2(n_101),
.B(n_103),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_588),
.B(n_108),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_628),
.A2(n_110),
.B(n_111),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_621),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_594),
.Y(n_669)
);

AOI222xp33_ASAP7_75t_L g670 ( 
.A1(n_616),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.C1(n_115),
.C2(n_117),
.Y(n_670)
);

BUFx12f_ASAP7_75t_L g671 ( 
.A(n_604),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_604),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_609),
.B(n_120),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_590),
.B(n_123),
.C(n_124),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_637),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_623),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_588),
.B(n_127),
.Y(n_677)
);

OAI21x1_ASAP7_75t_L g678 ( 
.A1(n_615),
.A2(n_128),
.B(n_130),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_595),
.A2(n_131),
.B(n_134),
.Y(n_679)
);

OAI221xp5_ASAP7_75t_L g680 ( 
.A1(n_605),
.A2(n_139),
.B1(n_142),
.B2(n_143),
.C(n_144),
.Y(n_680)
);

AO21x2_ASAP7_75t_L g681 ( 
.A1(n_613),
.A2(n_145),
.B(n_147),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_601),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_623),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_601),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_614),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_592),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_592),
.A2(n_148),
.B1(n_150),
.B2(n_153),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_610),
.A2(n_154),
.B1(n_155),
.B2(n_159),
.Y(n_688)
);

OA21x2_ASAP7_75t_L g689 ( 
.A1(n_619),
.A2(n_160),
.B(n_161),
.Y(n_689)
);

AOI21x1_ASAP7_75t_L g690 ( 
.A1(n_606),
.A2(n_162),
.B(n_163),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_630),
.A2(n_164),
.B(n_165),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_668),
.B(n_686),
.Y(n_692)
);

OAI21xp33_ASAP7_75t_SL g693 ( 
.A1(n_687),
.A2(n_634),
.B(n_627),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_682),
.Y(n_694)
);

O2A1O1Ixp5_ASAP7_75t_L g695 ( 
.A1(n_649),
.A2(n_624),
.B(n_633),
.C(n_635),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_669),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_684),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_668),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_676),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_683),
.Y(n_700)
);

CKINVDCx11_ASAP7_75t_R g701 ( 
.A(n_648),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_650),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_651),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_683),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_652),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_643),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_671),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_647),
.A2(n_678),
.B(n_658),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_663),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_669),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_675),
.Y(n_711)
);

CKINVDCx11_ASAP7_75t_R g712 ( 
.A(n_671),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_657),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_666),
.B(n_612),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_685),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_657),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_657),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_678),
.A2(n_639),
.B(n_617),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_655),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_690),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_664),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_664),
.B(n_639),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_681),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_642),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_656),
.B(n_612),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_646),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_681),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_677),
.B(n_612),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_644),
.A2(n_617),
.B(n_614),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_679),
.Y(n_730)
);

INVx4_ASAP7_75t_SL g731 ( 
.A(n_687),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_673),
.B(n_610),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_667),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_667),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_689),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_670),
.A2(n_617),
.B1(n_170),
.B2(n_171),
.Y(n_736)
);

OAI21x1_ASAP7_75t_L g737 ( 
.A1(n_689),
.A2(n_169),
.B(n_172),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_689),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_645),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_691),
.A2(n_173),
.B(n_176),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_680),
.A2(n_178),
.B1(n_179),
.B2(n_661),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_662),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_645),
.A2(n_654),
.B(n_649),
.Y(n_743)
);

AO21x2_ASAP7_75t_L g744 ( 
.A1(n_665),
.A2(n_661),
.B(n_654),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_640),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_653),
.B(n_640),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_659),
.B(n_641),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_672),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_701),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_R g750 ( 
.A(n_747),
.B(n_659),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_715),
.B(n_653),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_712),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_702),
.B(n_660),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_746),
.B(n_672),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_710),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_707),
.Y(n_756)
);

INVxp33_ASAP7_75t_L g757 ( 
.A(n_742),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_707),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_726),
.B(n_688),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_726),
.B(n_674),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_726),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_709),
.B(n_646),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_724),
.Y(n_763)
);

BUFx10_ASAP7_75t_L g764 ( 
.A(n_707),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_724),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_694),
.Y(n_766)
);

OR2x6_ASAP7_75t_L g767 ( 
.A(n_696),
.B(n_646),
.Y(n_767)
);

XNOR2xp5_ASAP7_75t_L g768 ( 
.A(n_746),
.B(n_641),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_709),
.B(n_732),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_R g770 ( 
.A(n_707),
.B(n_748),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_706),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_731),
.B(n_693),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_707),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_692),
.B(n_728),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_706),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_745),
.B(n_692),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_748),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_711),
.B(n_710),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_R g779 ( 
.A(n_748),
.B(n_696),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_711),
.B(n_705),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_705),
.B(n_719),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_R g782 ( 
.A(n_714),
.B(n_728),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_705),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_719),
.B(n_698),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_745),
.B(n_698),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_R g786 ( 
.A(n_714),
.B(n_725),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_731),
.B(n_725),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_731),
.B(n_748),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_748),
.B(n_731),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_694),
.Y(n_790)
);

BUFx10_ASAP7_75t_L g791 ( 
.A(n_697),
.Y(n_791)
);

OR2x4_ASAP7_75t_L g792 ( 
.A(n_697),
.B(n_704),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_693),
.B(n_740),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_700),
.B(n_704),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_722),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_766),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_776),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_SL g798 ( 
.A(n_752),
.B(n_743),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_774),
.B(n_766),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_769),
.B(n_700),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_790),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_787),
.B(n_739),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_776),
.B(n_739),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_792),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_789),
.B(n_733),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_772),
.B(n_717),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_755),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_781),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_763),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_794),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_751),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_765),
.B(n_699),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_791),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_778),
.B(n_738),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_795),
.B(n_783),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_780),
.Y(n_816)
);

NAND4xp25_ASAP7_75t_L g817 ( 
.A(n_793),
.B(n_736),
.C(n_741),
.D(n_695),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_758),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_784),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_753),
.B(n_723),
.C(n_727),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_785),
.B(n_713),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_791),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_779),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_771),
.B(n_738),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_775),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_754),
.B(n_727),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_785),
.B(n_717),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_789),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_796),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_799),
.B(n_735),
.Y(n_830)
);

OAI222xp33_ASAP7_75t_L g831 ( 
.A1(n_804),
.A2(n_760),
.B1(n_759),
.B2(n_788),
.C1(n_767),
.C2(n_722),
.Y(n_831)
);

AO21x2_ASAP7_75t_L g832 ( 
.A1(n_820),
.A2(n_723),
.B(n_735),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_806),
.B(n_716),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_796),
.Y(n_834)
);

AO21x2_ASAP7_75t_L g835 ( 
.A1(n_820),
.A2(n_716),
.B(n_713),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_806),
.B(n_734),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_802),
.B(n_734),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_809),
.B(n_757),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_802),
.B(n_733),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_807),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_811),
.B(n_754),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_801),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_804),
.Y(n_843)
);

NOR2x1_ASAP7_75t_L g844 ( 
.A(n_822),
.B(n_768),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_807),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_801),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_825),
.B(n_762),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_799),
.B(n_729),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_825),
.B(n_699),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_840),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_838),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_840),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_843),
.B(n_828),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_829),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_848),
.B(n_814),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_848),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_844),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_834),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_834),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_845),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_833),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_830),
.B(n_814),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_829),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_847),
.A2(n_817),
.B1(n_798),
.B2(n_744),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_843),
.B(n_833),
.Y(n_865)
);

OAI221xp5_ASAP7_75t_L g866 ( 
.A1(n_857),
.A2(n_817),
.B1(n_841),
.B2(n_749),
.C(n_823),
.Y(n_866)
);

AND2x4_ASAP7_75t_SL g867 ( 
.A(n_853),
.B(n_761),
.Y(n_867)
);

AO221x2_ASAP7_75t_L g868 ( 
.A1(n_860),
.A2(n_831),
.B1(n_822),
.B2(n_846),
.C(n_842),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_851),
.B(n_836),
.Y(n_869)
);

OAI22xp33_ASAP7_75t_L g870 ( 
.A1(n_861),
.A2(n_782),
.B1(n_786),
.B2(n_767),
.Y(n_870)
);

NAND2xp33_ASAP7_75t_SL g871 ( 
.A(n_853),
.B(n_750),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_862),
.B(n_836),
.Y(n_872)
);

OAI22xp33_ASAP7_75t_L g873 ( 
.A1(n_862),
.A2(n_760),
.B1(n_759),
.B2(n_828),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_855),
.B(n_846),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_855),
.B(n_839),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_869),
.B(n_865),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_874),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_867),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_872),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_875),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_868),
.B(n_865),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_873),
.B(n_864),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_870),
.B(n_856),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_871),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_866),
.Y(n_885)
);

NAND2x1_ASAP7_75t_L g886 ( 
.A(n_874),
.B(n_859),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_885),
.B(n_850),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_886),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_882),
.A2(n_826),
.B(n_756),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_884),
.B(n_852),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_884),
.B(n_852),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_878),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_892),
.B(n_881),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_887),
.B(n_889),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_890),
.B(n_877),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_891),
.B(n_880),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_895),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_893),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_896),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_894),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_SL g901 ( 
.A(n_900),
.B(n_888),
.C(n_883),
.Y(n_901)
);

NOR2x1p5_ASAP7_75t_L g902 ( 
.A(n_898),
.B(n_879),
.Y(n_902)
);

AOI211xp5_ASAP7_75t_L g903 ( 
.A1(n_897),
.A2(n_876),
.B(n_773),
.C(n_770),
.Y(n_903)
);

NOR2x1_ASAP7_75t_L g904 ( 
.A(n_899),
.B(n_818),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_899),
.B(n_813),
.Y(n_905)
);

NOR2x1_ASAP7_75t_L g906 ( 
.A(n_900),
.B(n_818),
.Y(n_906)
);

OAI21xp33_ASAP7_75t_L g907 ( 
.A1(n_898),
.A2(n_815),
.B(n_813),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_900),
.B(n_842),
.Y(n_908)
);

AOI211xp5_ASAP7_75t_L g909 ( 
.A1(n_901),
.A2(n_740),
.B(n_815),
.C(n_737),
.Y(n_909)
);

AOI221xp5_ASAP7_75t_L g910 ( 
.A1(n_907),
.A2(n_863),
.B1(n_854),
.B2(n_858),
.C(n_859),
.Y(n_910)
);

OAI211xp5_ASAP7_75t_SL g911 ( 
.A1(n_906),
.A2(n_854),
.B(n_859),
.C(n_858),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_902),
.Y(n_912)
);

AOI221x1_ASAP7_75t_L g913 ( 
.A1(n_904),
.A2(n_810),
.B1(n_819),
.B2(n_808),
.C(n_849),
.Y(n_913)
);

AOI221xp5_ASAP7_75t_L g914 ( 
.A1(n_905),
.A2(n_819),
.B1(n_810),
.B2(n_744),
.C(n_808),
.Y(n_914)
);

AOI221xp5_ASAP7_75t_L g915 ( 
.A1(n_903),
.A2(n_744),
.B1(n_832),
.B2(n_835),
.C(n_800),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_912),
.Y(n_916)
);

AND3x4_ASAP7_75t_L g917 ( 
.A(n_909),
.B(n_908),
.C(n_805),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_913),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_911),
.B(n_830),
.Y(n_919)
);

NAND2x1p5_ASAP7_75t_L g920 ( 
.A(n_910),
.B(n_737),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_915),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_914),
.B(n_839),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_R g923 ( 
.A(n_916),
.B(n_764),
.Y(n_923)
);

NAND2xp33_ASAP7_75t_SL g924 ( 
.A(n_918),
.B(n_917),
.Y(n_924)
);

NAND2xp33_ASAP7_75t_SL g925 ( 
.A(n_919),
.B(n_777),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_921),
.B(n_764),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_R g927 ( 
.A(n_922),
.B(n_812),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_920),
.B(n_805),
.Y(n_928)
);

XNOR2xp5_ASAP7_75t_L g929 ( 
.A(n_916),
.B(n_797),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_929),
.B(n_816),
.Y(n_930)
);

AOI21xp33_ASAP7_75t_SL g931 ( 
.A1(n_926),
.A2(n_832),
.B(n_835),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_924),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_928),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_925),
.A2(n_730),
.B(n_720),
.C(n_816),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_923),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_932),
.B(n_927),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_933),
.Y(n_937)
);

O2A1O1Ixp5_ASAP7_75t_L g938 ( 
.A1(n_935),
.A2(n_730),
.B(n_720),
.C(n_703),
.Y(n_938)
);

AO22x2_ASAP7_75t_L g939 ( 
.A1(n_937),
.A2(n_931),
.B1(n_934),
.B2(n_930),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_936),
.B(n_938),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_937),
.A2(n_824),
.B1(n_805),
.B2(n_722),
.Y(n_941)
);

AOI31xp33_ASAP7_75t_L g942 ( 
.A1(n_940),
.A2(n_824),
.A3(n_837),
.B(n_805),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_941),
.A2(n_832),
.B1(n_835),
.B2(n_837),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_942),
.A2(n_939),
.B(n_722),
.C(n_721),
.Y(n_944)
);

OAI322xp33_ASAP7_75t_L g945 ( 
.A1(n_943),
.A2(n_721),
.A3(n_703),
.B1(n_821),
.B2(n_827),
.C1(n_803),
.C2(n_718),
.Y(n_945)
);

AOI21x1_ASAP7_75t_L g946 ( 
.A1(n_944),
.A2(n_827),
.B(n_821),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_945),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_947),
.Y(n_948)
);

INVxp67_ASAP7_75t_SL g949 ( 
.A(n_946),
.Y(n_949)
);

AOI221xp5_ASAP7_75t_L g950 ( 
.A1(n_948),
.A2(n_949),
.B1(n_721),
.B2(n_703),
.C(n_803),
.Y(n_950)
);

AOI211xp5_ASAP7_75t_L g951 ( 
.A1(n_950),
.A2(n_729),
.B(n_718),
.C(n_708),
.Y(n_951)
);


endmodule