module fake_jpeg_3256_n_183 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_183);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_68),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_0),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_61),
.B1(n_59),
.B2(n_55),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_59),
.B1(n_49),
.B2(n_60),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_72),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_56),
.B1(n_51),
.B2(n_58),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_76),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_56),
.B1(n_51),
.B2(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_61),
.B1(n_57),
.B2(n_60),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_68),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_89),
.Y(n_102)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_2),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_54),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_45),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_50),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_70),
.B1(n_71),
.B2(n_50),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_103),
.B1(n_111),
.B2(n_113),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_76),
.B(n_74),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_7),
.B(n_9),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_45),
.B1(n_47),
.B2(n_3),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_102),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_82),
.A2(n_94),
.B1(n_81),
.B2(n_96),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_4),
.B(n_5),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_7),
.B(n_8),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_6),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_31),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_125),
.Y(n_137)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_20),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_SL g151 ( 
.A(n_122),
.B(n_32),
.C(n_42),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_130),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_90),
.C(n_86),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_110),
.C(n_103),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_127),
.C(n_132),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_6),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_19),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_11),
.Y(n_152)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_134),
.B(n_23),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_113),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_33),
.C(n_41),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_147),
.Y(n_160)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_156)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_10),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_149),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_152),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_127),
.B(n_122),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_155),
.B(n_157),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_128),
.B(n_13),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_15),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_15),
.B(n_16),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_34),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_161),
.Y(n_165)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_162),
.A2(n_150),
.B1(n_139),
.B2(n_135),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_135),
.B1(n_144),
.B2(n_140),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_141),
.B1(n_152),
.B2(n_151),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_170),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_161),
.C(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_172),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_163),
.C(n_157),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_176),
.A2(n_16),
.B(n_17),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_175),
.B1(n_177),
.B2(n_18),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_180),
.A2(n_24),
.B(n_38),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_39),
.C(n_40),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_43),
.Y(n_183)
);


endmodule