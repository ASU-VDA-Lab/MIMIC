module fake_jpeg_17564_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_68),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_17),
.B1(n_21),
.B2(n_27),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_27),
.B1(n_24),
.B2(n_56),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_17),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_17),
.B1(n_21),
.B2(n_27),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_20),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_87),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_90),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_43),
.B1(n_21),
.B2(n_44),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_79),
.B1(n_86),
.B2(n_88),
.Y(n_124)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_44),
.C(n_45),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_64),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_44),
.B1(n_24),
.B2(n_39),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_56),
.A2(n_34),
.B1(n_33),
.B2(n_20),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_33),
.B1(n_15),
.B2(n_11),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_99),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_93)
);

OAI22x1_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_102),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_48),
.A2(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_13),
.B1(n_12),
.B2(n_14),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_60),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_75),
.Y(n_123)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_40),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_100),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_37),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_13),
.B1(n_12),
.B2(n_14),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_100),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_106),
.C(n_108),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_63),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_117),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_23),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_50),
.B(n_23),
.C(n_31),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_111),
.B(n_19),
.C(n_31),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_23),
.B(n_31),
.C(n_15),
.Y(n_111)
);

NAND2x1_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_67),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_113),
.A2(n_19),
.B(n_84),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_63),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_80),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_101),
.B(n_85),
.Y(n_143)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_77),
.Y(n_157)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_67),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_63),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_63),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_63),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_86),
.B1(n_94),
.B2(n_79),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_142),
.B1(n_146),
.B2(n_149),
.Y(n_173)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_71),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_143),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_78),
.B(n_96),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_148),
.B(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_122),
.B(n_71),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_138),
.B(n_141),
.Y(n_193)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_90),
.B1(n_54),
.B2(n_62),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_101),
.C(n_36),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_130),
.C(n_107),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_62),
.B1(n_54),
.B2(n_97),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_111),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_0),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_124),
.A2(n_81),
.B1(n_72),
.B2(n_69),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx2_ASAP7_75t_R g151 ( 
.A(n_113),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_69),
.B1(n_35),
.B2(n_37),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_152),
.A2(n_156),
.B1(n_125),
.B2(n_77),
.Y(n_190)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_159),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_105),
.A2(n_35),
.B1(n_36),
.B2(n_61),
.Y(n_156)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_103),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_112),
.B(n_15),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_84),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_19),
.B(n_28),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_118),
.B1(n_103),
.B2(n_121),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_177),
.B1(n_182),
.B2(n_185),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_184),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_167),
.B(n_2),
.Y(n_223)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_103),
.Y(n_169)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_113),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_28),
.B1(n_22),
.B2(n_59),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_105),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_176),
.C(n_178),
.Y(n_207)
);

CKINVDCx10_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_121),
.B1(n_126),
.B2(n_112),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_104),
.C(n_128),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_126),
.B(n_128),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_181),
.A2(n_139),
.B1(n_153),
.B2(n_148),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_146),
.B1(n_162),
.B2(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_115),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_156),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_131),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_119),
.B1(n_125),
.B2(n_120),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_137),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_187),
.B(n_190),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_140),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_143),
.A2(n_35),
.B1(n_36),
.B2(n_73),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_185),
.B1(n_188),
.B2(n_163),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_196),
.B(n_19),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_199),
.A2(n_204),
.B(n_209),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_148),
.B1(n_147),
.B2(n_152),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_200),
.A2(n_202),
.B1(n_210),
.B2(n_211),
.Y(n_245)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_135),
.B1(n_154),
.B2(n_131),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_160),
.B1(n_133),
.B2(n_150),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_167),
.A2(n_73),
.B1(n_129),
.B2(n_3),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_171),
.B1(n_175),
.B2(n_182),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_216),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_181),
.A2(n_129),
.B1(n_28),
.B2(n_22),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_214),
.A2(n_224),
.B1(n_188),
.B2(n_186),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_1),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

A2O1A1O1Ixp25_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_28),
.B(n_22),
.C(n_11),
.D(n_4),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_196),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_22),
.B1(n_11),
.B2(n_3),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_219),
.B(n_220),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_1),
.Y(n_221)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_193),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_171),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_174),
.C(n_176),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_236),
.C(n_243),
.Y(n_259)
);

AND2x6_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_180),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_223),
.B1(n_218),
.B2(n_212),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_178),
.C(n_166),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_168),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_241),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_210),
.B1(n_214),
.B2(n_206),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_166),
.C(n_191),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_246),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_165),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_165),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_249),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_179),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_228),
.A2(n_217),
.B1(n_197),
.B2(n_200),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_258),
.B1(n_266),
.B2(n_232),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_199),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_251),
.B(n_237),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_208),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_260),
.C(n_261),
.Y(n_277)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_245),
.B1(n_232),
.B2(n_225),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_228),
.A2(n_209),
.B1(n_194),
.B2(n_224),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_204),
.C(n_179),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_195),
.C(n_194),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_215),
.B1(n_190),
.B2(n_170),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_59),
.C(n_6),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_269),
.C(n_247),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_59),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_278),
.B1(n_281),
.B2(n_279),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_235),
.Y(n_274)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_248),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_280),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_254),
.B1(n_263),
.B2(n_265),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_283),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_259),
.C(n_260),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_234),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_258),
.B(n_227),
.Y(n_282)
);

OAI321xp33_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_249),
.A3(n_238),
.B1(n_233),
.B2(n_242),
.C(n_5),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_252),
.C(n_262),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_268),
.Y(n_284)
);

NOR3xp33_ASAP7_75t_SL g287 ( 
.A(n_284),
.B(n_229),
.C(n_234),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_250),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_299),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_226),
.B1(n_253),
.B2(n_264),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_294),
.B1(n_277),
.B2(n_280),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_285),
.A2(n_226),
.B1(n_269),
.B2(n_240),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_8),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_293),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_283),
.A2(n_253),
.B1(n_264),
.B2(n_241),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_7),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_59),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_296),
.B(n_8),
.Y(n_309)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_5),
.B(n_6),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_302),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_6),
.C(n_7),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_7),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_303),
.B(n_304),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_7),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_306),
.B(n_308),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_309),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_8),
.C(n_294),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_287),
.B(n_296),
.Y(n_317)
);

INVx11_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_307),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_288),
.Y(n_319)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_320),
.B(n_322),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_314),
.A2(n_298),
.B1(n_290),
.B2(n_305),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_323),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_293),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

AOI322xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_315),
.A3(n_324),
.B1(n_311),
.B2(n_312),
.C1(n_321),
.C2(n_316),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_327),
.B(n_313),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_328),
.Y(n_329)
);


endmodule