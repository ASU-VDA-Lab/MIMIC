module fake_jpeg_12753_n_534 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_534);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_54),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_58),
.Y(n_150)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_59),
.Y(n_135)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_61),
.B(n_94),
.Y(n_113)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_34),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_63),
.B(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_65),
.B(n_70),
.Y(n_131)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_68),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_33),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_52),
.B1(n_23),
.B2(n_43),
.Y(n_123)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_40),
.B(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_95),
.Y(n_121)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_104),
.Y(n_134)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_97),
.Y(n_124)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_42),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_22),
.B(n_2),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_100),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_22),
.B(n_39),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_47),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_49),
.B1(n_25),
.B2(n_44),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_105),
.A2(n_148),
.B1(n_152),
.B2(n_50),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_56),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_111),
.B(n_127),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_60),
.A2(n_33),
.B1(n_47),
.B2(n_48),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_112),
.A2(n_114),
.B1(n_122),
.B2(n_149),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_75),
.A2(n_33),
.B1(n_47),
.B2(n_48),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_26),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_137),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_83),
.A2(n_48),
.B1(n_47),
.B2(n_37),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_123),
.A2(n_38),
.B1(n_27),
.B2(n_43),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_56),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_66),
.B(n_26),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_68),
.B(n_25),
.C(n_44),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_24),
.C(n_50),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_53),
.A2(n_37),
.B1(n_44),
.B2(n_32),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_101),
.A2(n_47),
.B1(n_48),
.B2(n_32),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_55),
.A2(n_37),
.B1(n_44),
.B2(n_32),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_104),
.A2(n_39),
.B1(n_37),
.B2(n_32),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_43),
.B1(n_35),
.B2(n_31),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_92),
.B(n_52),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_157),
.B(n_160),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_121),
.A2(n_131),
.B1(n_118),
.B2(n_134),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_163),
.A2(n_202),
.B1(n_203),
.B2(n_217),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_165),
.B(n_170),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_166),
.B(n_188),
.C(n_209),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_167),
.Y(n_267)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_171),
.Y(n_256)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_174),
.A2(n_196),
.B1(n_206),
.B2(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_176),
.Y(n_271)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_177),
.Y(n_241)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_178),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_105),
.A2(n_24),
.B1(n_50),
.B2(n_148),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_152),
.A2(n_24),
.B1(n_52),
.B2(n_35),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_182),
.B(n_189),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_35),
.B(n_23),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_184),
.A2(n_128),
.B(n_5),
.Y(n_265)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_113),
.A2(n_59),
.B(n_3),
.Y(n_187)
);

HAxp5_ASAP7_75t_SL g262 ( 
.A(n_187),
.B(n_2),
.CON(n_262),
.SN(n_262)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_102),
.C(n_98),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_116),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_110),
.B(n_58),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_190),
.B(n_194),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_135),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_191),
.B(n_198),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_192),
.Y(n_227)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_193),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_142),
.B(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_126),
.B(n_89),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_195),
.B(n_208),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_116),
.A2(n_57),
.B1(n_91),
.B2(n_79),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_197),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_117),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_133),
.A2(n_27),
.B1(n_23),
.B2(n_30),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_199),
.A2(n_200),
.B1(n_218),
.B2(n_158),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_133),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_125),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_201),
.B(n_207),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_115),
.A2(n_78),
.B1(n_71),
.B2(n_69),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_204),
.A2(n_216),
.B1(n_154),
.B2(n_144),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_145),
.B(n_31),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_210),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_145),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_125),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_109),
.A2(n_28),
.B(n_63),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_76),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_108),
.B(n_151),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_108),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_214),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_106),
.A2(n_38),
.B1(n_73),
.B2(n_102),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_151),
.B(n_48),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_107),
.A2(n_38),
.B1(n_132),
.B2(n_130),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_159),
.A2(n_38),
.B1(n_48),
.B2(n_74),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_129),
.A2(n_74),
.B1(n_3),
.B2(n_4),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_129),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_219),
.Y(n_247)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_107),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_215),
.B(n_167),
.C(n_172),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_222),
.A2(n_265),
.B(n_207),
.Y(n_305)
);

O2A1O1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_117),
.B(n_158),
.C(n_155),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_224),
.B(n_262),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_234),
.A2(n_169),
.B1(n_168),
.B2(n_171),
.Y(n_287)
);

OAI22x1_ASAP7_75t_SL g235 ( 
.A1(n_164),
.A2(n_155),
.B1(n_150),
.B2(n_138),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_235),
.A2(n_264),
.B1(n_217),
.B2(n_211),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_165),
.B(n_159),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_243),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_183),
.B(n_153),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_163),
.A2(n_119),
.B1(n_153),
.B2(n_146),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_245),
.A2(n_252),
.B1(n_266),
.B2(n_14),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_170),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_183),
.B(n_146),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_254),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_194),
.B(n_138),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_195),
.C(n_210),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_215),
.B(n_147),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_250),
.B(n_258),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_202),
.A2(n_132),
.B1(n_130),
.B2(n_119),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_128),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_186),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_188),
.B(n_147),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_175),
.A2(n_154),
.B1(n_144),
.B2(n_6),
.Y(n_266)
);

OAI32xp33_ASAP7_75t_L g270 ( 
.A1(n_214),
.A2(n_4),
.A3(n_5),
.B1(n_7),
.B2(n_10),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_204),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_273),
.B(n_247),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_221),
.A2(n_184),
.B(n_186),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_274),
.A2(n_265),
.B(n_267),
.Y(n_331)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_222),
.A2(n_166),
.B(n_190),
.C(n_177),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_277),
.B(n_290),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_278),
.B(n_292),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_251),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_279),
.B(n_282),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_244),
.B(n_178),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_280),
.B(n_237),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_221),
.B(n_185),
.C(n_211),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_303),
.C(n_306),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_268),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_283),
.B(n_312),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_284),
.Y(n_338)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_240),
.A2(n_204),
.B1(n_189),
.B2(n_201),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_296),
.B1(n_308),
.B2(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_231),
.B(n_208),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_182),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_231),
.B(n_212),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_293),
.B(n_300),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_227),
.Y(n_294)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_294),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_240),
.A2(n_264),
.B1(n_228),
.B2(n_253),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_297),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_258),
.A2(n_220),
.B1(n_180),
.B2(n_197),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_298),
.A2(n_302),
.B1(n_316),
.B2(n_238),
.Y(n_333)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_299),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_243),
.B(n_219),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_263),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_314),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_229),
.A2(n_220),
.B1(n_180),
.B2(n_176),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_249),
.B(n_173),
.C(n_193),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_248),
.B(n_4),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_304),
.B(n_307),
.Y(n_355)
);

AO21x1_ASAP7_75t_SL g339 ( 
.A1(n_305),
.A2(n_259),
.B(n_270),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_223),
.B(n_192),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_233),
.B(n_5),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_228),
.A2(n_5),
.B1(n_7),
.B2(n_10),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_253),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_242),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_310),
.A2(n_245),
.B1(n_252),
.B2(n_266),
.Y(n_344)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_241),
.Y(n_311)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_250),
.B(n_13),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_313),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_257),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_236),
.B(n_14),
.C(n_15),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_317),
.C(n_227),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_236),
.B(n_14),
.C(n_16),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_254),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_233),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_237),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_319),
.B(n_350),
.C(n_360),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_305),
.A2(n_295),
.B(n_288),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_323),
.A2(n_332),
.B(n_339),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_314),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_327),
.B(n_18),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_290),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_329),
.B(n_356),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_331),
.B(n_307),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_295),
.A2(n_224),
.B(n_235),
.Y(n_332)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_333),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_302),
.A2(n_259),
.B1(n_224),
.B2(n_229),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_334),
.A2(n_347),
.B1(n_354),
.B2(n_308),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_232),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_337),
.B(n_341),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_291),
.A2(n_271),
.B(n_239),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_340),
.A2(n_293),
.B(n_282),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_280),
.B(n_232),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_344),
.A2(n_353),
.B1(n_298),
.B2(n_299),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_316),
.A2(n_239),
.B1(n_226),
.B2(n_247),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_279),
.B(n_269),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_348),
.B(n_315),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_296),
.A2(n_226),
.B1(n_225),
.B2(n_230),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_318),
.A2(n_225),
.B1(n_230),
.B2(n_256),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_SL g357 ( 
.A1(n_295),
.A2(n_256),
.B(n_16),
.C(n_18),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_300),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_297),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_281),
.B(n_16),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_322),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_361),
.B(n_367),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_324),
.B(n_272),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_362),
.B(n_392),
.Y(n_398)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_354),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_365),
.B(n_368),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_274),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_366),
.B(n_375),
.C(n_326),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_352),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_370),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_320),
.A2(n_303),
.B1(n_273),
.B2(n_277),
.Y(n_371)
);

OAI21xp33_ASAP7_75t_L g426 ( 
.A1(n_371),
.A2(n_357),
.B(n_330),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_352),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_373),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_342),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_342),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_374),
.B(n_376),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_326),
.B(n_306),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_320),
.A2(n_275),
.B1(n_286),
.B2(n_283),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_329),
.B(n_275),
.Y(n_378)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_342),
.A2(n_286),
.B1(n_304),
.B2(n_311),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_379),
.B(n_386),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_355),
.Y(n_416)
);

A2O1A1O1Ixp25_ASAP7_75t_L g382 ( 
.A1(n_328),
.A2(n_276),
.B(n_285),
.C(n_289),
.D(n_312),
.Y(n_382)
);

NOR3xp33_ASAP7_75t_L g410 ( 
.A(n_382),
.B(n_385),
.C(n_349),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_384),
.A2(n_336),
.B1(n_333),
.B2(n_327),
.Y(n_413)
);

OAI32xp33_ASAP7_75t_L g386 ( 
.A1(n_328),
.A2(n_294),
.A3(n_309),
.B1(n_310),
.B2(n_284),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_347),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_387),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_388),
.B(n_391),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_355),
.Y(n_389)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_389),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_344),
.A2(n_18),
.B1(n_317),
.B2(n_353),
.Y(n_390)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_390),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_321),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_340),
.A2(n_336),
.B1(n_339),
.B2(n_334),
.Y(n_394)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_394),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_321),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_395),
.B(n_359),
.Y(n_397)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_397),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_370),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_372),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_401),
.B(n_408),
.C(n_415),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_402),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_364),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_410),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_360),
.C(n_319),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_413),
.A2(n_383),
.B1(n_376),
.B2(n_387),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_366),
.B(n_323),
.C(n_331),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_416),
.B(n_381),
.Y(n_431)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_396),
.Y(n_418)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_418),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_381),
.B(n_356),
.C(n_332),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_380),
.C(n_367),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_393),
.A2(n_343),
.B(n_351),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_422),
.A2(n_427),
.B(n_373),
.Y(n_430)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_378),
.Y(n_424)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_424),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_369),
.Y(n_438)
);

A2O1A1Ixp33_ASAP7_75t_SL g427 ( 
.A1(n_393),
.A2(n_357),
.B(n_330),
.C(n_346),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_422),
.A2(n_394),
.B(n_374),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_432),
.Y(n_464)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_430),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_431),
.B(n_424),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_400),
.A2(n_383),
.B(n_371),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_434),
.A2(n_425),
.B1(n_417),
.B2(n_421),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_453),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_404),
.B(n_389),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_436),
.B(n_440),
.Y(n_462)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_437),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_451),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_398),
.B(n_392),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_401),
.B(n_379),
.C(n_368),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_442),
.C(n_445),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_384),
.C(n_382),
.Y(n_442)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_407),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_448),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_403),
.A2(n_365),
.B1(n_395),
.B2(n_391),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_446),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_408),
.B(n_351),
.C(n_346),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_386),
.B1(n_363),
.B2(n_390),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_420),
.A2(n_335),
.B1(n_345),
.B2(n_343),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_409),
.B(n_345),
.Y(n_450)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_450),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_357),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_357),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_439),
.Y(n_455)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_455),
.Y(n_475)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_450),
.Y(n_461)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_461),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_400),
.C(n_420),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_463),
.B(n_465),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_421),
.C(n_412),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_452),
.Y(n_466)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_466),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_471),
.C(n_473),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_433),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_468),
.A2(n_470),
.B1(n_474),
.B2(n_448),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_414),
.C(n_425),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_435),
.B(n_413),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_433),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_464),
.A2(n_428),
.B(n_432),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_476),
.A2(n_479),
.B(n_486),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g478 ( 
.A(n_462),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_478),
.B(n_458),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_454),
.A2(n_430),
.B(n_414),
.Y(n_479)
);

NOR3xp33_ASAP7_75t_SL g480 ( 
.A(n_457),
.B(n_405),
.C(n_406),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_488),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_485),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_454),
.A2(n_411),
.B(n_446),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_484),
.A2(n_449),
.B1(n_397),
.B2(n_427),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_471),
.A2(n_429),
.B(n_442),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_460),
.A2(n_439),
.B(n_447),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_487),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_431),
.C(n_451),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_444),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_491),
.Y(n_501)
);

NOR3xp33_ASAP7_75t_SL g491 ( 
.A(n_456),
.B(n_405),
.C(n_406),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_465),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_492),
.B(n_497),
.Y(n_511)
);

AOI21xp33_ASAP7_75t_SL g494 ( 
.A1(n_476),
.A2(n_463),
.B(n_472),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_500),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_487),
.A2(n_470),
.B1(n_456),
.B2(n_452),
.Y(n_496)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_496),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_477),
.B(n_473),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_483),
.A2(n_417),
.B1(n_411),
.B2(n_449),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_505),
.C(n_503),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_477),
.B(n_458),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_479),
.A2(n_438),
.B(n_472),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_502),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_484),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_338),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_453),
.Y(n_505)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_507),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_510),
.A2(n_493),
.B1(n_502),
.B2(n_494),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_495),
.B(n_488),
.C(n_475),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_514),
.Y(n_524)
);

AOI322xp5_ASAP7_75t_L g514 ( 
.A1(n_496),
.A2(n_491),
.A3(n_484),
.B1(n_480),
.B2(n_489),
.C1(n_418),
.C2(n_423),
.Y(n_514)
);

A2O1A1Ixp33_ASAP7_75t_L g515 ( 
.A1(n_501),
.A2(n_490),
.B(n_467),
.C(n_397),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_515),
.A2(n_498),
.B(n_505),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_493),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_338),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g523 ( 
.A(n_517),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_518),
.A2(n_521),
.B(n_513),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_519),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_520),
.A2(n_510),
.B(n_513),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_511),
.A2(n_423),
.B(n_427),
.Y(n_521)
);

BUFx24_ASAP7_75t_SL g525 ( 
.A(n_522),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_525),
.A2(n_526),
.B(n_528),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_527),
.A2(n_508),
.B(n_524),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_530),
.B(n_519),
.C(n_427),
.Y(n_532)
);

OAI22xp33_ASAP7_75t_L g531 ( 
.A1(n_529),
.A2(n_509),
.B1(n_514),
.B2(n_523),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_531),
.B(n_532),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_427),
.Y(n_534)
);


endmodule