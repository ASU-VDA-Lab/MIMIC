module fake_jpeg_5944_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx24_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_17),
.B(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_14),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_12),
.B1(n_11),
.B2(n_14),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_18),
.B(n_20),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_21),
.B(n_16),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_16),
.C(n_19),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_34),
.C(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_22),
.A2(n_13),
.B(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_39),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_15),
.B(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_23),
.B(n_28),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_42),
.B(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_2),
.Y(n_44)
);

AOI31xp33_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_46),
.A3(n_3),
.B(n_4),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_37),
.B1(n_24),
.B2(n_6),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g48 ( 
.A(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_45),
.Y(n_49)
);

BUFx24_ASAP7_75t_SL g50 ( 
.A(n_49),
.Y(n_50)
);


endmodule