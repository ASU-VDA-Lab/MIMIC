module fake_netlist_1_605_n_24 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_24);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_24;
wire n_20;
wire n_23;
wire n_22;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
wire n_21;
OR2x6_ASAP7_75t_L g12 ( .A(n_1), .B(n_10), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_5), .B(n_11), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
OR2x2_ASAP7_75t_L g15 ( .A(n_4), .B(n_2), .Y(n_15) );
OAI22xp33_ASAP7_75t_L g16 ( .A1(n_7), .A2(n_1), .B1(n_6), .B2(n_3), .Y(n_16) );
NOR2xp33_ASAP7_75t_R g17 ( .A(n_13), .B(n_8), .Y(n_17) );
NAND3xp33_ASAP7_75t_SL g18 ( .A(n_15), .B(n_0), .C(n_3), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
O2A1O1Ixp33_ASAP7_75t_SL g21 ( .A1(n_20), .A2(n_18), .B(n_14), .C(n_16), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
AOI21xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_12), .B(n_4), .Y(n_24) );
endmodule