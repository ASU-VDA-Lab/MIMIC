module real_jpeg_31464_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_0),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_0),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_0),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_1),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_1),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_1),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_1),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_1),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_1),
.B(n_63),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_2),
.B(n_449),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_2),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_3),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_3),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_3),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_3),
.B(n_56),
.Y(n_269)
);

AND2x2_ASAP7_75t_SL g331 ( 
.A(n_3),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_3),
.B(n_371),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_4),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_5),
.Y(n_130)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_6),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_7),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_7),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_7),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_7),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_7),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_7),
.B(n_247),
.Y(n_246)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_82),
.Y(n_81)
);

NAND2x1_ASAP7_75t_L g92 ( 
.A(n_8),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_8),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_8),
.B(n_29),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_8),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_9),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_9),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_9),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_9),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_9),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_SL g354 ( 
.A(n_9),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_9),
.B(n_369),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_10),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_11),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_11),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_13),
.Y(n_120)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_13),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_14),
.B(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_14),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_14),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_14),
.B(n_128),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_14),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_14),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_14),
.B(n_387),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_15),
.Y(n_141)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_15),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_16),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_16),
.B(n_108),
.Y(n_107)
);

AND2x4_ASAP7_75t_SL g172 ( 
.A(n_16),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_16),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_16),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_17),
.B(n_33),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_17),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_17),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g254 ( 
.A(n_17),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_17),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_17),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_17),
.B(n_335),
.Y(n_334)
);

OAI311xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_230),
.A3(n_448),
.B1(n_450),
.C1(n_453),
.Y(n_18)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_19),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_228),
.Y(n_19)
);

NOR2x1_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_183),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_L g229 ( 
.A(n_21),
.B(n_183),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_101),
.C(n_131),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_23),
.B(n_101),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_68),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_24),
.B(n_100),
.C(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.C(n_54),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_26),
.B(n_40),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_27),
.B(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_27),
.A2(n_28),
.B1(n_302),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_28),
.A2(n_103),
.B(n_110),
.Y(n_102)
);

OAI221xp5_ASAP7_75t_L g110 ( 
.A1(n_28),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.C(n_109),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_28),
.B(n_35),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_28),
.B(n_35),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_28),
.B(n_104),
.C(n_106),
.Y(n_194)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_29),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_31),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_34),
.Y(n_177)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_34),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_35),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_35),
.A2(n_38),
.B1(n_245),
.B2(n_246),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_36),
.Y(n_369)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_37),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

MAJx2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_46),
.C(n_50),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_41),
.B(n_46),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_45),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_45),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_48),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_49),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_49),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_50),
.A2(n_51),
.B1(n_223),
.B2(n_227),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_50),
.B(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_53),
.Y(n_257)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_54),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_62),
.C(n_66),
.Y(n_77)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_78),
.B1(n_99),
.B2(n_100),
.Y(n_68)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_77),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_71),
.B(n_75),
.C(n_77),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_72),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_72),
.A2(n_75),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_78),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_91),
.C(n_96),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_79),
.A2(n_80),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.C(n_88),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_88),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_85),
.B(n_107),
.Y(n_297)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_98),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_111),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_102),
.B(n_112),
.C(n_115),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_109),
.Y(n_103)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_106),
.A2(n_107),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_114),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_114),
.A2(n_278),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_171),
.C(n_175),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_116),
.B(n_218),
.C(n_219),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_116),
.A2(n_117),
.B1(n_175),
.B2(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_120),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_120),
.Y(n_383)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_132),
.B(n_438),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_157),
.C(n_179),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_134),
.B(n_426),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.C(n_143),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_135),
.B(n_137),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_137),
.A2(n_138),
.B(n_142),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_143),
.B(n_415),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_150),
.C(n_153),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_144),
.A2(n_145),
.B1(n_153),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_150),
.B(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_153),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_156),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_158),
.B(n_180),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_170),
.B(n_178),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_164),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_160),
.B(n_164),
.Y(n_410)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_169),
.Y(n_284)
);

XNOR2x2_ASAP7_75t_L g409 ( 
.A(n_170),
.B(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_171),
.B(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_173),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_174),
.Y(n_360)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_175),
.Y(n_290)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_203),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_202),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_213),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_251),
.C(n_254),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_208),
.B(n_251),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_209),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_220),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g220 ( 
.A(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_230),
.B(n_451),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_435),
.B(n_445),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_418),
.B(n_431),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_402),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_311),
.B(n_401),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_291),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_235),
.B(n_291),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_259),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_237),
.B(n_274),
.C(n_404),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_242),
.B2(n_258),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_238),
.B(n_243),
.C(n_250),
.Y(n_407)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_249),
.B2(n_250),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_253),
.B(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_274),
.Y(n_259)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_260),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.C(n_273),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_263),
.B(n_273),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_269),
.C(n_270),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_265),
.B(n_271),
.Y(n_344)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_269),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2x2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_288),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_276),
.B(n_288),
.C(n_417),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_277),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.C(n_285),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_280),
.B1(n_285),
.B2(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_296),
.B(n_305),
.C(n_308),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_292),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_293),
.A2(n_296),
.B1(n_309),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_293),
.Y(n_399)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.C(n_301),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_297),
.Y(n_349)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_301),
.B(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_305),
.A2(n_306),
.B1(n_397),
.B2(n_398),
.Y(n_396)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_393),
.B(n_400),
.Y(n_311)
);

OAI21xp33_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_350),
.B(n_392),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_340),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_314),
.B(n_340),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_330),
.C(n_337),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_315),
.A2(n_316),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_324),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_323),
.C(n_324),
.Y(n_342)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_330),
.A2(n_337),
.B1(n_338),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_330),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_334),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_334),
.Y(n_353)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx4f_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_347),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_345),
.B2(n_346),
.Y(n_341)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_342),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_343),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_343),
.B(n_345),
.C(n_395),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_347),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_365),
.B(n_391),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_361),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_361),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.C(n_357),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_354),
.A2(n_357),
.B1(n_358),
.B2(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_354),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_378),
.B(n_390),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_375),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_367),
.B(n_375),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_370),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_368),
.B(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_SL g371 ( 
.A(n_372),
.Y(n_371)
);

INVx8_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_385),
.B(n_389),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_384),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_384),
.Y(n_389)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_396),
.Y(n_400)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_405),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_405),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_413),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_414),
.C(n_416),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_409),
.C(n_411),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

AOI21x1_ASAP7_75t_L g432 ( 
.A1(n_419),
.A2(n_433),
.B(n_434),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_421),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_422),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_424),
.A2(n_425),
.B1(n_427),
.B2(n_428),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_428),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVxp33_ASAP7_75t_SL g435 ( 
.A(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_439),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_437),
.B(n_439),
.Y(n_447)
);

MAJx2_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_442),
.C(n_444),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_446),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_448),
.B(n_452),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_448),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);


endmodule