module fake_jpeg_9202_n_171 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_171);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_6),
.B(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_42),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_50),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_21),
.B1(n_32),
.B2(n_20),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_22),
.B1(n_33),
.B2(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_20),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_21),
.B1(n_24),
.B2(n_16),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_66),
.B1(n_23),
.B2(n_40),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_16),
.B1(n_15),
.B2(n_30),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_74),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_81),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_23),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_76),
.Y(n_103)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_80),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_90),
.B1(n_56),
.B2(n_51),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_43),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_43),
.B(n_41),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_52),
.B(n_49),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_88),
.Y(n_101)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_55),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_49),
.Y(n_91)
);

XNOR2x1_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_91),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_70),
.B1(n_86),
.B2(n_77),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_106),
.B(n_108),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_52),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_88),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_39),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_39),
.B(n_3),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_2),
.B(n_3),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_2),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_114),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_90),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_125),
.C(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_116),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_122),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_89),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_67),
.B1(n_64),
.B2(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_87),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_87),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_113),
.C(n_100),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_99),
.B(n_118),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_99),
.B(n_106),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_122),
.B(n_125),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_84),
.B1(n_75),
.B2(n_70),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_121),
.B1(n_96),
.B2(n_64),
.Y(n_143)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_141),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_135),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_146),
.B1(n_148),
.B2(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_138),
.B(n_137),
.C(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_109),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_147),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_121),
.B1(n_96),
.B2(n_73),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_105),
.C(n_73),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_152),
.B(n_140),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_131),
.B1(n_8),
.B2(n_10),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_154),
.Y(n_160)
);

OAI321xp33_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_14),
.C(n_3),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_144),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_155),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_4),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_161),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_147),
.C(n_150),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_158),
.A2(n_146),
.B1(n_152),
.B2(n_4),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_164),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_162),
.C(n_166),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_169),
.C(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_160),
.Y(n_171)
);


endmodule