module fake_jpeg_8181_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_SL g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_26),
.B1(n_14),
.B2(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_15),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_1),
.B1(n_9),
.B2(n_4),
.Y(n_26)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_26),
.B(n_22),
.C(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_24),
.C(n_27),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_45),
.C(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_48),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_17),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_18),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_12),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_34),
.C(n_11),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_12),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_30),
.C(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_55),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_51),
.C(n_52),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_30),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_45),
.C(n_39),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_17),
.C(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_SL g66 ( 
.A(n_63),
.B(n_17),
.C(n_4),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_61),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_17),
.B(n_20),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_66),
.B(n_60),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_58),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_70),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_67),
.C(n_68),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_69),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.B1(n_20),
.B2(n_27),
.Y(n_76)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_27),
.A3(n_13),
.B1(n_8),
.B2(n_2),
.C1(n_36),
.C2(n_31),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_36),
.Y(n_78)
);


endmodule