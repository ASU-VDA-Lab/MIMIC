module fake_jpeg_22481_n_101 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_32),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_29),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_18),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_24),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_25),
.A2(n_24),
.B1(n_15),
.B2(n_16),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_20),
.B1(n_16),
.B2(n_15),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_48),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_23),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_21),
.C(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_21),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_63),
.C(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_56),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_42),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_22),
.B1(n_17),
.B2(n_5),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_65),
.B1(n_2),
.B2(n_9),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_44),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_41),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_2),
.B1(n_3),
.B2(n_8),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_51),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_76),
.C(n_68),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_75),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_10),
.B1(n_42),
.B2(n_50),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_65),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_70),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_53),
.B1(n_64),
.B2(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_83),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_73),
.C(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_78),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_88),
.C(n_77),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_90),
.A2(n_93),
.B1(n_58),
.B2(n_72),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_62),
.C(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_89),
.B(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_81),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_79),
.B1(n_84),
.B2(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_96),
.B(n_90),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_98),
.B(n_95),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_10),
.Y(n_101)
);


endmodule