module fake_jpeg_25381_n_322 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_22),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_25),
.Y(n_48)
);

CKINVDCx9p33_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_19),
.B(n_8),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_43),
.B(n_26),
.C(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_17),
.B1(n_27),
.B2(n_33),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_69),
.B1(n_43),
.B2(n_36),
.Y(n_78)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_56),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_17),
.B1(n_27),
.B2(n_33),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_43),
.B1(n_26),
.B2(n_36),
.Y(n_74)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_17),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_43),
.B1(n_35),
.B2(n_38),
.Y(n_84)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_43),
.B1(n_35),
.B2(n_38),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_92),
.B1(n_36),
.B2(n_61),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_52),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_86),
.C(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_78),
.B1(n_40),
.B2(n_39),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_79),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_64),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_69),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_45),
.B(n_43),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_38),
.C(n_44),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_45),
.A2(n_35),
.B1(n_38),
.B2(n_36),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_19),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_70),
.B(n_76),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_67),
.B1(n_49),
.B2(n_35),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_113),
.B1(n_123),
.B2(n_109),
.Y(n_132)
);

OA22x2_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_38),
.B1(n_49),
.B2(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_114),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_35),
.B1(n_51),
.B2(n_36),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_102),
.A2(n_77),
.B1(n_89),
.B2(n_87),
.Y(n_141)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_70),
.B(n_36),
.CI(n_39),
.CON(n_105),
.SN(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_122),
.B(n_116),
.C(n_100),
.D(n_114),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_68),
.B1(n_58),
.B2(n_57),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_34),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_122),
.B1(n_96),
.B2(n_84),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_40),
.B(n_39),
.C(n_60),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_39),
.B(n_40),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_118),
.Y(n_140)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_124),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_86),
.B1(n_84),
.B2(n_96),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_145),
.B1(n_150),
.B2(n_99),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_29),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_26),
.B(n_19),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_134),
.B(n_146),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_132),
.A2(n_148),
.B1(n_34),
.B2(n_18),
.Y(n_175)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_136),
.B(n_144),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_40),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_112),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_103),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_139),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_103),
.A2(n_79),
.B1(n_21),
.B2(n_30),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_89),
.B1(n_87),
.B2(n_82),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_107),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_147),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_82),
.B1(n_95),
.B2(n_77),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_40),
.B1(n_39),
.B2(n_32),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_90),
.C(n_64),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_116),
.C(n_104),
.Y(n_159)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_24),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_107),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_154),
.B(n_21),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_106),
.A2(n_30),
.B(n_21),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_139),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_142),
.Y(n_189)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_99),
.A3(n_116),
.B1(n_108),
.B2(n_29),
.Y(n_157)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_166),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_132),
.B1(n_136),
.B2(n_133),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_99),
.C(n_112),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_164),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_124),
.B1(n_104),
.B2(n_111),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_163),
.A2(n_133),
.B1(n_135),
.B2(n_128),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_111),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_173),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_170),
.B(n_179),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_90),
.C(n_23),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_130),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_24),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_175),
.A2(n_140),
.B1(n_20),
.B2(n_22),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_23),
.C(n_20),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_125),
.B(n_20),
.Y(n_183)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_154),
.B(n_24),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_185),
.Y(n_190)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_126),
.B(n_146),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_204),
.B(n_169),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_201),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_149),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_191),
.B(n_197),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_199),
.B1(n_175),
.B2(n_156),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_194),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_160),
.B1(n_158),
.B2(n_182),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_195),
.A2(n_211),
.B1(n_28),
.B2(n_18),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_14),
.C(n_15),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_135),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_25),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_22),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_208),
.B(n_181),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_212),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_128),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_181),
.A2(n_140),
.B(n_24),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_164),
.C(n_161),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_218),
.C(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_174),
.C(n_159),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_209),
.B1(n_188),
.B2(n_212),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_220),
.A2(n_192),
.B1(n_202),
.B2(n_189),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_222),
.A2(n_208),
.B(n_204),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_239)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_230),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_156),
.B1(n_183),
.B2(n_165),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_226),
.A2(n_228),
.B1(n_28),
.B2(n_23),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_178),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_233),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_157),
.B1(n_168),
.B2(n_172),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_171),
.C(n_166),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_192),
.A2(n_170),
.B(n_172),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_SL g258 ( 
.A(n_232),
.B(n_23),
.C(n_1),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_168),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_28),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_235),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_18),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_23),
.C(n_22),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_203),
.C(n_20),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_257),
.B1(n_6),
.B2(n_14),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_210),
.B1(n_190),
.B2(n_202),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_244),
.A2(n_250),
.B1(n_23),
.B2(n_1),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_245),
.A2(n_254),
.B(n_258),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_203),
.B1(n_28),
.B2(n_18),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_251),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_215),
.B(n_227),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_248),
.B(n_8),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_213),
.A2(n_220),
.B1(n_234),
.B2(n_214),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_221),
.B(n_10),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_229),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_10),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_24),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_255),
.A2(n_228),
.B1(n_216),
.B2(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_259),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_218),
.C(n_231),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_270),
.C(n_6),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_266),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_232),
.B1(n_222),
.B2(n_224),
.Y(n_266)
);

O2A1O1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_217),
.B(n_237),
.C(n_2),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_267),
.A2(n_245),
.B(n_254),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_273),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_271),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_65),
.C(n_9),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_240),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_252),
.B(n_7),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_249),
.B1(n_241),
.B2(n_250),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_262),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_278),
.B(n_285),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_265),
.A2(n_257),
.B(n_240),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_256),
.B1(n_2),
.B2(n_3),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_284),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_6),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_269),
.Y(n_289)
);

AO22x1_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_287),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_12),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_263),
.C(n_271),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_13),
.C(n_15),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_260),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_296),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_270),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_272),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_284),
.C(n_283),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_277),
.A2(n_12),
.B(n_13),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_299),
.A2(n_297),
.B(n_280),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_301),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_279),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_303),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_286),
.C(n_282),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_288),
.B1(n_282),
.B2(n_285),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_308),
.C(n_291),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_2),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_305),
.B(n_308),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_313),
.B(n_4),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_312),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_292),
.C(n_289),
.Y(n_312)
);

A2O1A1O1Ixp25_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_299),
.B(n_4),
.C(n_5),
.D(n_3),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_317),
.C(n_309),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_316),
.B(n_4),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_319),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_5),
.C(n_310),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_5),
.Y(n_322)
);


endmodule