module fake_ariane_2449_n_879 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_879);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_879;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_670;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_761;
wire n_818;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_218;
wire n_839;
wire n_770;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_277;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_362;
wire n_260;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

BUFx3_ASAP7_75t_L g194 ( 
.A(n_7),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_43),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_175),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_136),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_151),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_7),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_67),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_14),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_50),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_72),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_39),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_74),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_68),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_107),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_128),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_10),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_46),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_146),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_71),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_75),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_102),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_64),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_123),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_36),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_178),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_99),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_63),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_167),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_91),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_0),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_85),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_162),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_188),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_122),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_18),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_15),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_84),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_70),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_133),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_160),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_154),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_176),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_164),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_88),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_150),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_112),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_33),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_32),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_156),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_105),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_10),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_81),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_83),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_25),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_22),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_193),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_187),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_3),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_87),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_127),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_179),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_97),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_158),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_58),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_114),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_89),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_42),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_5),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_54),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_110),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_L g274 ( 
.A(n_23),
.B(n_101),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_52),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_121),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_79),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_172),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_194),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_203),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_216),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_194),
.Y(n_282)
);

OA21x2_ASAP7_75t_L g283 ( 
.A1(n_200),
.A2(n_0),
.B(n_1),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_202),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_205),
.B(n_2),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_212),
.Y(n_286)
);

BUFx6f_ASAP7_75t_SL g287 ( 
.A(n_253),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_198),
.A2(n_232),
.B1(n_236),
.B2(n_201),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

BUFx8_ASAP7_75t_SL g290 ( 
.A(n_240),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_237),
.B(n_4),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_241),
.B(n_4),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_207),
.B(n_5),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_199),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_6),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_208),
.B(n_6),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_257),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_297)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_216),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_269),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_217),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_261),
.Y(n_304)
);

AOI22x1_ASAP7_75t_SL g305 ( 
.A1(n_220),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_224),
.B(n_12),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_216),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_13),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_197),
.B(n_13),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g310 ( 
.A(n_195),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_225),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_197),
.Y(n_312)
);

BUFx12f_ASAP7_75t_L g313 ( 
.A(n_196),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_216),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_262),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_233),
.Y(n_318)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_262),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_242),
.B(n_14),
.Y(n_320)
);

OA21x2_ASAP7_75t_L g321 ( 
.A1(n_247),
.A2(n_15),
.B(n_16),
.Y(n_321)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_215),
.B(n_17),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_249),
.B(n_19),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_250),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_251),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_259),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_263),
.B(n_192),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_276),
.B(n_20),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_204),
.Y(n_331)
);

BUFx12f_ASAP7_75t_L g332 ( 
.A(n_206),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_267),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_290),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_310),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_294),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_313),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_282),
.B(n_273),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_332),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_281),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_286),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_286),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_299),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_304),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_314),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_288),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_R g352 ( 
.A(n_301),
.B(n_209),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_288),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_333),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_R g355 ( 
.A(n_301),
.B(n_278),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_331),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_311),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_331),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_279),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_287),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_279),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_316),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_302),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_287),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_302),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_307),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_318),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g369 ( 
.A(n_295),
.B(n_226),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_307),
.Y(n_370)
);

NAND2xp33_ASAP7_75t_R g371 ( 
.A(n_321),
.B(n_210),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_285),
.Y(n_372)
);

AOI21x1_ASAP7_75t_L g373 ( 
.A1(n_324),
.A2(n_256),
.B(n_223),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_317),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_317),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_303),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_326),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_325),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_327),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_334),
.Y(n_380)
);

BUFx10_ASAP7_75t_L g381 ( 
.A(n_295),
.Y(n_381)
);

NAND2xp33_ASAP7_75t_R g382 ( 
.A(n_321),
.B(n_211),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_309),
.B(n_274),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_330),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_285),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_291),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_312),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_292),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_308),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_389),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_376),
.B(n_309),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_345),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_323),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_298),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_356),
.B(n_293),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_306),
.Y(n_398)
);

AND2x6_ASAP7_75t_L g399 ( 
.A(n_344),
.B(n_324),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_335),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_363),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_298),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_339),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_369),
.B(n_298),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_386),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_350),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_319),
.Y(n_409)
);

A2O1A1Ixp33_ASAP7_75t_L g410 ( 
.A1(n_387),
.A2(n_320),
.B(n_296),
.C(n_328),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_319),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_377),
.B(n_296),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_379),
.B(n_320),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_338),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_328),
.C(n_297),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_381),
.B(n_297),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_366),
.B(n_280),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_300),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_384),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_349),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_378),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g423 ( 
.A1(n_373),
.A2(n_283),
.B(n_319),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_368),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_381),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_385),
.B(n_322),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_360),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_390),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_L g429 ( 
.A(n_352),
.B(n_213),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_362),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_369),
.B(n_322),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_370),
.B(n_322),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_374),
.B(n_315),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_355),
.B(n_329),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_375),
.B(n_315),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_388),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_361),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_365),
.B(n_329),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_372),
.B(n_214),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_337),
.B(n_218),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_364),
.B(n_219),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_357),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_371),
.B(n_284),
.C(n_283),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_348),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_354),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_336),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_340),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_342),
.B(n_221),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_351),
.B(n_222),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_353),
.Y(n_452)
);

INVx8_ASAP7_75t_L g453 ( 
.A(n_383),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_376),
.B(n_284),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_376),
.B(n_227),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_383),
.B(n_228),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_335),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_389),
.B(n_230),
.Y(n_458)
);

INVx8_ASAP7_75t_L g459 ( 
.A(n_383),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_383),
.B(n_234),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_422),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_396),
.B(n_235),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_424),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_393),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_401),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_406),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_427),
.Y(n_468)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_418),
.B(n_239),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_398),
.B(n_458),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_391),
.B(n_243),
.Y(n_472)
);

OAI22xp33_ASAP7_75t_L g473 ( 
.A1(n_416),
.A2(n_305),
.B1(n_277),
.B2(n_275),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_399),
.A2(n_407),
.B1(n_444),
.B2(n_412),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_430),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_451),
.B(n_244),
.Y(n_476)
);

INVx8_ASAP7_75t_L g477 ( 
.A(n_453),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_425),
.B(n_245),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_400),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_454),
.A2(n_270),
.B1(n_268),
.B2(n_265),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_403),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_450),
.B(n_246),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_414),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_404),
.Y(n_484)
);

NOR2xp67_ASAP7_75t_L g485 ( 
.A(n_447),
.B(n_248),
.Y(n_485)
);

NAND3xp33_ASAP7_75t_L g486 ( 
.A(n_419),
.B(n_264),
.C(n_260),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_21),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_410),
.A2(n_413),
.B1(n_437),
.B2(n_428),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_421),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_415),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_399),
.B(n_252),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_457),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_446),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_459),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_459),
.A2(n_258),
.B1(n_255),
.B2(n_27),
.Y(n_495)
);

NAND2x1p5_ASAP7_75t_L g496 ( 
.A(n_438),
.B(n_24),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_406),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_443),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_406),
.Y(n_499)
);

AND2x4_ASAP7_75t_SL g500 ( 
.A(n_448),
.B(n_26),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_441),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_408),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_408),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_442),
.B(n_28),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_432),
.B(n_29),
.Y(n_505)
);

CKINVDCx8_ASAP7_75t_R g506 ( 
.A(n_399),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_408),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_420),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_440),
.Y(n_509)
);

NOR2x1_ASAP7_75t_L g510 ( 
.A(n_439),
.B(n_30),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_456),
.B(n_31),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_420),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_399),
.B(n_191),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_417),
.B(n_34),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_392),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_460),
.B(n_40),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_435),
.B(n_41),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_420),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_445),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_394),
.B(n_44),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_455),
.B(n_45),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_429),
.B(n_47),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_395),
.A2(n_402),
.B1(n_405),
.B2(n_411),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_449),
.B(n_190),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_423),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_452),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_434),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_436),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_433),
.B(n_409),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_475),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_501),
.B(n_452),
.Y(n_531)
);

NAND2x1p5_ASAP7_75t_L g532 ( 
.A(n_465),
.B(n_409),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_463),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_R g534 ( 
.A(n_477),
.B(n_431),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_471),
.A2(n_426),
.B1(n_49),
.B2(n_51),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_483),
.B(n_426),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_469),
.B(n_494),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_489),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_469),
.B(n_494),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_482),
.B(n_462),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_477),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_509),
.B(n_48),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_525),
.A2(n_53),
.B(n_55),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_478),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_464),
.Y(n_545)
);

NOR3xp33_ASAP7_75t_L g546 ( 
.A(n_519),
.B(n_56),
.C(n_57),
.Y(n_546)
);

O2A1O1Ixp33_ASAP7_75t_L g547 ( 
.A1(n_488),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_461),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_527),
.B(n_62),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_525),
.A2(n_65),
.B(n_66),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_528),
.B(n_498),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_466),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_505),
.B(n_69),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_505),
.B(n_73),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_469),
.B(n_76),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_484),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_472),
.A2(n_77),
.B(n_78),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_529),
.A2(n_80),
.B(n_82),
.Y(n_558)
);

A2O1A1Ixp33_ASAP7_75t_SL g559 ( 
.A1(n_524),
.A2(n_86),
.B(n_90),
.C(n_92),
.Y(n_559)
);

OAI21xp33_ASAP7_75t_L g560 ( 
.A1(n_480),
.A2(n_93),
.B(n_94),
.Y(n_560)
);

INVx6_ASAP7_75t_L g561 ( 
.A(n_478),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_514),
.B(n_95),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_474),
.B(n_96),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_R g564 ( 
.A(n_506),
.B(n_98),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_526),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_468),
.Y(n_566)
);

INVx3_ASAP7_75t_SL g567 ( 
.A(n_500),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_520),
.A2(n_100),
.B(n_103),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_491),
.A2(n_104),
.B(n_106),
.Y(n_569)
);

AO32x2_ASAP7_75t_L g570 ( 
.A1(n_493),
.A2(n_108),
.A3(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_494),
.Y(n_571)
);

NOR3xp33_ASAP7_75t_SL g572 ( 
.A(n_473),
.B(n_470),
.C(n_486),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_513),
.A2(n_115),
.B(n_116),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_490),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_468),
.B(n_117),
.Y(n_575)
);

CKINVDCx8_ASAP7_75t_R g576 ( 
.A(n_487),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_512),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_476),
.B(n_118),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_495),
.A2(n_120),
.B1(n_124),
.B2(n_125),
.Y(n_579)
);

O2A1O1Ixp33_ASAP7_75t_SL g580 ( 
.A1(n_521),
.A2(n_126),
.B(n_129),
.C(n_130),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_504),
.A2(n_511),
.B(n_516),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_496),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_479),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_497),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_485),
.B(n_131),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_499),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_522),
.A2(n_132),
.B(n_134),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_538),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_566),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_551),
.B(n_481),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_544),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_540),
.A2(n_517),
.B(n_512),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_537),
.Y(n_593)
);

NAND2x1p5_ASAP7_75t_L g594 ( 
.A(n_537),
.B(n_467),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_530),
.Y(n_595)
);

NAND2x1p5_ASAP7_75t_L g596 ( 
.A(n_539),
.B(n_467),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_577),
.Y(n_597)
);

BUFx2_ASAP7_75t_SL g598 ( 
.A(n_539),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_545),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_544),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_533),
.Y(n_601)
);

CKINVDCx6p67_ASAP7_75t_R g602 ( 
.A(n_567),
.Y(n_602)
);

BUFx12f_ASAP7_75t_L g603 ( 
.A(n_565),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_571),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_571),
.Y(n_605)
);

INVx8_ASAP7_75t_L g606 ( 
.A(n_541),
.Y(n_606)
);

AO21x2_ASAP7_75t_L g607 ( 
.A1(n_563),
.A2(n_507),
.B(n_503),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_556),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_552),
.Y(n_609)
);

OAI21x1_ASAP7_75t_L g610 ( 
.A1(n_581),
.A2(n_510),
.B(n_523),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_561),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_576),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_584),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_561),
.A2(n_515),
.B1(n_487),
.B2(n_518),
.Y(n_614)
);

OAI21x1_ASAP7_75t_L g615 ( 
.A1(n_573),
.A2(n_518),
.B(n_502),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_548),
.B(n_492),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_574),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_532),
.Y(n_618)
);

NAND2x1p5_ASAP7_75t_L g619 ( 
.A(n_582),
.B(n_502),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_575),
.A2(n_508),
.B(n_487),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_536),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_584),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_583),
.B(n_487),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_578),
.A2(n_135),
.B(n_137),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_586),
.B(n_138),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_586),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_562),
.A2(n_139),
.B(n_140),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_549),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_531),
.B(n_141),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_557),
.A2(n_142),
.B(n_143),
.Y(n_630)
);

BUFx2_ASAP7_75t_SL g631 ( 
.A(n_555),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_564),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_568),
.A2(n_144),
.B(n_145),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_534),
.Y(n_634)
);

BUFx12f_ASAP7_75t_L g635 ( 
.A(n_603),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_602),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_SL g637 ( 
.A1(n_590),
.A2(n_553),
.B1(n_554),
.B2(n_579),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_589),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_621),
.A2(n_560),
.B1(n_542),
.B2(n_546),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_589),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_599),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_603),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_609),
.A2(n_572),
.B1(n_547),
.B2(n_535),
.Y(n_643)
);

INVx6_ASAP7_75t_L g644 ( 
.A(n_593),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_595),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_595),
.B(n_585),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_601),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_601),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_616),
.A2(n_543),
.B1(n_550),
.B2(n_569),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_608),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_616),
.A2(n_587),
.B1(n_558),
.B2(n_570),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_608),
.Y(n_652)
);

AOI21x1_ASAP7_75t_L g653 ( 
.A1(n_620),
.A2(n_559),
.B(n_570),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_588),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_612),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_617),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_597),
.B(n_147),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_597),
.B(n_148),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_604),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_606),
.Y(n_660)
);

NAND2x1p5_ASAP7_75t_L g661 ( 
.A(n_612),
.B(n_593),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_611),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_617),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_606),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_632),
.B(n_570),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_606),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_612),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_SL g668 ( 
.A1(n_631),
.A2(n_580),
.B1(n_152),
.B2(n_153),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_628),
.B(n_626),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_614),
.A2(n_149),
.B1(n_155),
.B2(n_157),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_598),
.B(n_159),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_613),
.B(n_626),
.Y(n_672)
);

AO21x1_ASAP7_75t_L g673 ( 
.A1(n_623),
.A2(n_161),
.B(n_163),
.Y(n_673)
);

OA21x2_ASAP7_75t_L g674 ( 
.A1(n_615),
.A2(n_165),
.B(n_166),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_622),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_613),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_622),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_638),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_640),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_SL g680 ( 
.A1(n_670),
.A2(n_612),
.B1(n_629),
.B2(n_625),
.Y(n_680)
);

INVx6_ASAP7_75t_L g681 ( 
.A(n_667),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_641),
.Y(n_682)
);

CKINVDCx11_ASAP7_75t_R g683 ( 
.A(n_635),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_654),
.B(n_591),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_636),
.B(n_600),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_659),
.Y(n_686)
);

NOR2x1p5_ASAP7_75t_L g687 ( 
.A(n_642),
.B(n_602),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_645),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_647),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_655),
.B(n_604),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_654),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_663),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_R g693 ( 
.A(n_655),
.B(n_605),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_648),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_650),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_662),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_652),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_644),
.Y(n_698)
);

NOR3xp33_ASAP7_75t_SL g699 ( 
.A(n_643),
.B(n_592),
.C(n_625),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_662),
.B(n_605),
.Y(n_700)
);

NAND3xp33_ASAP7_75t_L g701 ( 
.A(n_637),
.B(n_618),
.C(n_619),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_656),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_661),
.B(n_594),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_669),
.B(n_594),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_669),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_672),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_667),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_657),
.B(n_596),
.Y(n_708)
);

AOI221xp5_ASAP7_75t_L g709 ( 
.A1(n_643),
.A2(n_634),
.B1(n_619),
.B2(n_596),
.C(n_607),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_661),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_637),
.A2(n_607),
.B1(n_610),
.B2(n_630),
.Y(n_711)
);

AO31x2_ASAP7_75t_L g712 ( 
.A1(n_673),
.A2(n_620),
.A3(n_615),
.B(n_610),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_646),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_644),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_644),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_658),
.B(n_665),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_676),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_660),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_675),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_646),
.Y(n_720)
);

AND2x2_ASAP7_75t_SL g721 ( 
.A(n_671),
.B(n_624),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_677),
.B(n_624),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_639),
.B(n_627),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_674),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_682),
.B(n_651),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_691),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_722),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_689),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_686),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_716),
.B(n_651),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_705),
.B(n_653),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_707),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_705),
.B(n_674),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_717),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_678),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_694),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_704),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_713),
.B(n_670),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_678),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_695),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_697),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_713),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_698),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_720),
.B(n_706),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_702),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_703),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_720),
.Y(n_747)
);

NOR2x1_ASAP7_75t_SL g748 ( 
.A(n_701),
.B(n_703),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_679),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_688),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_722),
.B(n_668),
.Y(n_751)
);

AND2x4_ASAP7_75t_SL g752 ( 
.A(n_690),
.B(n_666),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_724),
.B(n_630),
.Y(n_753)
);

OA21x2_ASAP7_75t_L g754 ( 
.A1(n_711),
.A2(n_633),
.B(n_649),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_699),
.B(n_721),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_719),
.B(n_668),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_692),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_719),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_712),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_708),
.B(n_649),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_684),
.B(n_633),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_712),
.B(n_690),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_700),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_741),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_734),
.B(n_696),
.Y(n_765)
);

AND2x4_ASAP7_75t_SL g766 ( 
.A(n_743),
.B(n_698),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_741),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_742),
.B(n_709),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_728),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_735),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_736),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_729),
.B(n_685),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_740),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_726),
.B(n_685),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_735),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_745),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_739),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_744),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_739),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_747),
.B(n_723),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_737),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_763),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_743),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_730),
.B(n_725),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_730),
.B(n_710),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_749),
.Y(n_786)
);

NOR2xp67_ASAP7_75t_L g787 ( 
.A(n_743),
.B(n_714),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_750),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_757),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_760),
.B(n_727),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_780),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_790),
.B(n_727),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_784),
.B(n_725),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_785),
.B(n_760),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_772),
.B(n_762),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_765),
.B(n_762),
.Y(n_796)
);

NOR2x1_ASAP7_75t_L g797 ( 
.A(n_774),
.B(n_732),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_767),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_780),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_769),
.B(n_755),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_771),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_773),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_776),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_781),
.B(n_755),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_782),
.B(n_751),
.Y(n_805)
);

XOR2xp5_ASAP7_75t_L g806 ( 
.A(n_794),
.B(n_718),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_791),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_793),
.B(n_791),
.Y(n_808)
);

O2A1O1Ixp5_ASAP7_75t_R g809 ( 
.A1(n_800),
.A2(n_768),
.B(n_732),
.C(n_783),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_800),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_797),
.B(n_761),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_796),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_799),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_798),
.Y(n_814)
);

AND2x2_ASAP7_75t_SL g815 ( 
.A(n_805),
.B(n_768),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_810),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_814),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_815),
.A2(n_804),
.B1(n_805),
.B2(n_756),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_812),
.B(n_792),
.Y(n_819)
);

OAI22xp33_ASAP7_75t_L g820 ( 
.A1(n_809),
.A2(n_751),
.B1(n_799),
.B2(n_756),
.Y(n_820)
);

NAND2x1_ASAP7_75t_SL g821 ( 
.A(n_818),
.B(n_811),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_819),
.B(n_811),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_817),
.B(n_813),
.C(n_807),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_820),
.B(n_813),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_816),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_817),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_824),
.B(n_807),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_826),
.B(n_803),
.Y(n_828)
);

AOI221xp5_ASAP7_75t_L g829 ( 
.A1(n_823),
.A2(n_802),
.B1(n_801),
.B2(n_778),
.C(n_806),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_822),
.B(n_683),
.Y(n_830)
);

NOR3xp33_ASAP7_75t_SL g831 ( 
.A(n_830),
.B(n_821),
.C(n_687),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_829),
.A2(n_825),
.B1(n_680),
.B2(n_786),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_827),
.B(n_714),
.C(n_715),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_832),
.A2(n_828),
.B(n_808),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_833),
.A2(n_787),
.B(n_758),
.Y(n_835)
);

AOI322xp5_ASAP7_75t_L g836 ( 
.A1(n_831),
.A2(n_795),
.A3(n_738),
.B1(n_761),
.B2(n_733),
.C1(n_731),
.C2(n_759),
.Y(n_836)
);

OAI221xp5_ASAP7_75t_SL g837 ( 
.A1(n_832),
.A2(n_738),
.B1(n_753),
.B2(n_759),
.C(n_731),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_836),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_835),
.B(n_664),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_834),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_837),
.B(n_766),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_834),
.B(n_752),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_834),
.A2(n_754),
.B1(n_788),
.B2(n_789),
.Y(n_843)
);

AOI221xp5_ASAP7_75t_L g844 ( 
.A1(n_834),
.A2(n_759),
.B1(n_733),
.B2(n_789),
.C(n_788),
.Y(n_844)
);

AOI221xp5_ASAP7_75t_L g845 ( 
.A1(n_840),
.A2(n_779),
.B1(n_752),
.B2(n_764),
.C(n_715),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_838),
.B(n_783),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_842),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_839),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_844),
.B(n_766),
.Y(n_849)
);

OR5x1_ASAP7_75t_L g850 ( 
.A(n_841),
.B(n_693),
.C(n_748),
.D(n_681),
.E(n_753),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_843),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_842),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_846),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_847),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_848),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_852),
.B(n_754),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_851),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_850),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_849),
.Y(n_859)
);

NAND5xp2_ASAP7_75t_L g860 ( 
.A(n_845),
.B(n_681),
.C(n_746),
.D(n_754),
.E(n_753),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_854),
.Y(n_861)
);

AND4x1_ASAP7_75t_L g862 ( 
.A(n_857),
.B(n_168),
.C(n_169),
.D(n_170),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_855),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_855),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_853),
.Y(n_865)
);

AO22x2_ASAP7_75t_L g866 ( 
.A1(n_859),
.A2(n_775),
.B1(n_777),
.B2(n_770),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_864),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_865),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_863),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_861),
.B(n_858),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_SL g871 ( 
.A1(n_862),
.A2(n_860),
.B1(n_856),
.B2(n_746),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_868),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_869),
.A2(n_866),
.B1(n_753),
.B2(n_746),
.Y(n_873)
);

OAI321xp33_ASAP7_75t_L g874 ( 
.A1(n_872),
.A2(n_870),
.A3(n_867),
.B1(n_871),
.B2(n_746),
.C(n_770),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_873),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_874),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_876),
.A2(n_875),
.B(n_870),
.Y(n_877)
);

OR2x6_ASAP7_75t_L g878 ( 
.A(n_877),
.B(n_171),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_878),
.A2(n_777),
.B1(n_173),
.B2(n_177),
.Y(n_879)
);


endmodule