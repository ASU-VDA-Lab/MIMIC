module fake_ibex_223_n_1382 (n_151, n_147, n_85, n_251, n_167, n_128, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_250, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1382);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_250;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1382;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_433;
wire n_262;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_1301;
wire n_257;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_870;
wire n_1298;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_252;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_256;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_258;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_291;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_266;
wire n_1339;
wire n_485;
wire n_1315;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_260;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_255;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_326;
wire n_270;
wire n_1340;
wire n_259;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_253;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_354;
wire n_1057;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1374;
wire n_792;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_478;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_254;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g252 ( 
.A(n_145),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_215),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_139),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_180),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_11),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_82),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_236),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_49),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_26),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_101),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_131),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_188),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_39),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_130),
.B(n_6),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_127),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_164),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_184),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_177),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_L g272 ( 
.A(n_192),
.B(n_162),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_172),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_193),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_167),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_3),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_147),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_93),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_85),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_52),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_156),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_37),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_152),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_174),
.B(n_217),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_227),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_15),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_74),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_166),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_121),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_123),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_98),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_83),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_56),
.B(n_62),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_4),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_74),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_129),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_56),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_201),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_39),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_114),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_191),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_2),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_171),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_47),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_126),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_36),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_211),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_213),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_212),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_207),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_222),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_117),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_221),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_118),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_239),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_105),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_175),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_203),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_51),
.Y(n_323)
);

BUFx8_ASAP7_75t_SL g324 ( 
.A(n_178),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_103),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_122),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_232),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_88),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_169),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_9),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_78),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_94),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_13),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_66),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_21),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_73),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_229),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_8),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_206),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_199),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_163),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_77),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_47),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_234),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_33),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_198),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_5),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_61),
.Y(n_348)
);

BUFx10_ASAP7_75t_L g349 ( 
.A(n_5),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_250),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_135),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_61),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_204),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_161),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_246),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_168),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_86),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_69),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_4),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_194),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_155),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_189),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_35),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_216),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_240),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_200),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_140),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_119),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_251),
.Y(n_369)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_233),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_176),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_243),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_108),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_53),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_148),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_132),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_219),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_97),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_110),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_84),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_159),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_170),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_19),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_113),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_21),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_72),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_42),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_73),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_81),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_49),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_134),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_214),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_51),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_197),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_53),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_183),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_165),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_143),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_31),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_208),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_158),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_72),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_60),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_66),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_146),
.B(n_151),
.Y(n_405)
);

BUFx10_ASAP7_75t_L g406 ( 
.A(n_45),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_27),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_6),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_181),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_87),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_196),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_112),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_19),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_149),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_179),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_120),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_142),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_136),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_144),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_79),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_60),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_157),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_182),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_195),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_185),
.Y(n_425)
);

BUFx10_ASAP7_75t_L g426 ( 
.A(n_230),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_128),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_80),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_54),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_133),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_68),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_65),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_1),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_96),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_210),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_218),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_242),
.Y(n_437)
);

INVx6_ASAP7_75t_L g438 ( 
.A(n_305),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_260),
.B(n_0),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_373),
.B(n_2),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_387),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_282),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_293),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_263),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_293),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_381),
.B(n_7),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_296),
.B(n_10),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_316),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_282),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_316),
.Y(n_450)
);

OA21x2_ASAP7_75t_L g451 ( 
.A1(n_257),
.A2(n_90),
.B(n_89),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_347),
.B(n_10),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_299),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_453)
);

OA21x2_ASAP7_75t_L g454 ( 
.A1(n_257),
.A2(n_92),
.B(n_91),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_419),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_301),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_347),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_386),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_282),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_346),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_386),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_433),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_301),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_266),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_293),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_315),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_271),
.B(n_16),
.Y(n_467)
);

NOR2x1_ASAP7_75t_L g468 ( 
.A(n_276),
.B(n_95),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_315),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_292),
.A2(n_100),
.B(n_99),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_305),
.Y(n_471)
);

AND2x2_ASAP7_75t_SL g472 ( 
.A(n_258),
.B(n_102),
.Y(n_472)
);

BUFx8_ASAP7_75t_SL g473 ( 
.A(n_299),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_307),
.A2(n_106),
.B(n_104),
.Y(n_474)
);

BUFx12f_ASAP7_75t_L g475 ( 
.A(n_305),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_280),
.Y(n_476)
);

BUFx12f_ASAP7_75t_L g477 ( 
.A(n_426),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_304),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_282),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_315),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_315),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_426),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_412),
.B(n_17),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_346),
.B(n_17),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_282),
.Y(n_486)
);

OAI22x1_ASAP7_75t_R g487 ( 
.A1(n_331),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_310),
.B(n_18),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_370),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_370),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_426),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_391),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_391),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_392),
.Y(n_495)
);

INVx5_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

AOI22x1_ASAP7_75t_SL g497 ( 
.A1(n_331),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_370),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_392),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_L g500 ( 
.A(n_370),
.B(n_107),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_370),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_281),
.B(n_23),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_370),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_307),
.A2(n_137),
.B(n_248),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_385),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_412),
.B(n_24),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_366),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_366),
.B(n_319),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_385),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_323),
.B(n_24),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_422),
.B(n_25),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_324),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_335),
.Y(n_513)
);

BUFx8_ASAP7_75t_L g514 ( 
.A(n_370),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_371),
.B(n_25),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_349),
.B(n_26),
.Y(n_516)
);

NOR2x1_ASAP7_75t_L g517 ( 
.A(n_336),
.B(n_109),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_385),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_385),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_402),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_402),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_320),
.B(n_341),
.Y(n_522)
);

INVx6_ASAP7_75t_L g523 ( 
.A(n_349),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_256),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_255),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_320),
.A2(n_141),
.B(n_247),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_341),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_402),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_402),
.Y(n_529)
);

BUFx12f_ASAP7_75t_L g530 ( 
.A(n_349),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_377),
.A2(n_138),
.B(n_244),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_377),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_397),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_338),
.Y(n_534)
);

AOI22x1_ASAP7_75t_SL g535 ( 
.A1(n_348),
.A2(n_388),
.B1(n_428),
.B2(n_283),
.Y(n_535)
);

CKINVDCx6p67_ASAP7_75t_R g536 ( 
.A(n_269),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_406),
.B(n_27),
.Y(n_537)
);

INVx6_ASAP7_75t_L g538 ( 
.A(n_406),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_400),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_343),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_400),
.B(n_28),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_401),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_348),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_492),
.B(n_259),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_514),
.B(n_401),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_452),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_452),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_514),
.B(n_414),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_514),
.B(n_414),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_452),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_534),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_512),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_471),
.B(n_430),
.Y(n_553)
);

BUFx6f_ASAP7_75t_SL g554 ( 
.A(n_472),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_442),
.Y(n_555)
);

INVx8_ASAP7_75t_L g556 ( 
.A(n_475),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_530),
.B(n_359),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_484),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_442),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_534),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_449),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_484),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_523),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_447),
.Y(n_564)
);

AOI21x1_ASAP7_75t_L g565 ( 
.A1(n_470),
.A2(n_504),
.B(n_474),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_459),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_459),
.Y(n_567)
);

AND3x2_ASAP7_75t_L g568 ( 
.A(n_456),
.B(n_324),
.C(n_363),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_508),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_530),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_527),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_471),
.B(n_374),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_479),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_527),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_441),
.A2(n_288),
.B1(n_297),
.B2(n_287),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_479),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_483),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_492),
.B(n_306),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_490),
.Y(n_581)
);

INVx8_ASAP7_75t_L g582 ( 
.A(n_475),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_490),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_491),
.Y(n_584)
);

AOI21x1_ASAP7_75t_L g585 ( 
.A1(n_470),
.A2(n_254),
.B(n_252),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_491),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_523),
.B(n_330),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_498),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_498),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_542),
.Y(n_591)
);

HAxp5_ASAP7_75t_SL g592 ( 
.A(n_535),
.B(n_388),
.CON(n_592),
.SN(n_592)
);

INVxp67_ASAP7_75t_R g593 ( 
.A(n_487),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_501),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_444),
.B(n_334),
.C(n_333),
.Y(n_595)
);

AO21x2_ASAP7_75t_L g596 ( 
.A1(n_474),
.A2(n_405),
.B(n_264),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_512),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_464),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_503),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_L g600 ( 
.A(n_471),
.B(n_265),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_532),
.B(n_533),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_503),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_482),
.B(n_438),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_476),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_482),
.B(n_342),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_532),
.B(n_262),
.Y(n_606)
);

INVx8_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_L g608 ( 
.A1(n_462),
.A2(n_428),
.B1(n_395),
.B2(n_399),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_522),
.B(n_270),
.Y(n_609)
);

BUFx6f_ASAP7_75t_SL g610 ( 
.A(n_472),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_478),
.Y(n_611)
);

NAND3xp33_ASAP7_75t_L g612 ( 
.A(n_455),
.B(n_352),
.C(n_345),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_445),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_523),
.B(n_358),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_438),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_532),
.B(n_268),
.Y(n_616)
);

NOR2x1p5_ASAP7_75t_L g617 ( 
.A(n_477),
.B(n_393),
.Y(n_617)
);

AND3x2_ASAP7_75t_L g618 ( 
.A(n_463),
.B(n_431),
.C(n_407),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_482),
.B(n_383),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_513),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_525),
.B(n_390),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_532),
.B(n_273),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_525),
.B(n_438),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_465),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_466),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_536),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_461),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_532),
.B(n_275),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_446),
.B(n_267),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_540),
.Y(n_630)
);

AOI21x1_ASAP7_75t_L g631 ( 
.A1(n_504),
.A2(n_531),
.B(n_526),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_525),
.B(n_278),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_466),
.Y(n_633)
);

AND3x2_ASAP7_75t_L g634 ( 
.A(n_511),
.B(n_290),
.C(n_279),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_538),
.B(n_403),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_466),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_461),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_466),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_SL g639 ( 
.A(n_506),
.B(n_269),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_469),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_469),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g642 ( 
.A(n_522),
.B(n_506),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_469),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_461),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_446),
.A2(n_410),
.B1(n_408),
.B2(n_404),
.Y(n_645)
);

INVx8_ASAP7_75t_L g646 ( 
.A(n_522),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_469),
.Y(n_647)
);

BUFx10_ASAP7_75t_L g648 ( 
.A(n_467),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_524),
.B(n_302),
.Y(n_649)
);

INVxp67_ASAP7_75t_R g650 ( 
.A(n_516),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_480),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_457),
.Y(n_652)
);

CKINVDCx6p67_ASAP7_75t_R g653 ( 
.A(n_536),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_448),
.Y(n_654)
);

AND2x6_ASAP7_75t_L g655 ( 
.A(n_516),
.B(n_303),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_481),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_448),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_533),
.B(n_309),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_481),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_485),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_539),
.B(n_450),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_485),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_539),
.B(n_314),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_485),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_450),
.B(n_317),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_458),
.Y(n_666)
);

AO22x2_ASAP7_75t_L g667 ( 
.A1(n_497),
.A2(n_326),
.B1(n_327),
.B2(n_318),
.Y(n_667)
);

AND2x2_ASAP7_75t_SL g668 ( 
.A(n_500),
.B(n_332),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_488),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_460),
.B(n_413),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_510),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_460),
.B(n_440),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_489),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_511),
.B(n_420),
.Y(n_674)
);

AND3x1_ASAP7_75t_L g675 ( 
.A(n_537),
.B(n_356),
.C(n_351),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_L g676 ( 
.A(n_453),
.B(n_295),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_539),
.B(n_357),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_539),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_522),
.Y(n_679)
);

AO21x2_ASAP7_75t_L g680 ( 
.A1(n_531),
.A2(n_362),
.B(n_360),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_522),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_537),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_494),
.Y(n_683)
);

NOR2x1p5_ASAP7_75t_L g684 ( 
.A(n_473),
.B(n_421),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_473),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_494),
.Y(n_686)
);

BUFx6f_ASAP7_75t_SL g687 ( 
.A(n_509),
.Y(n_687)
);

INVx8_ASAP7_75t_L g688 ( 
.A(n_507),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_541),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_669),
.B(n_671),
.Y(n_690)
);

INVxp67_ASAP7_75t_SL g691 ( 
.A(n_578),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_564),
.B(n_467),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_544),
.B(n_502),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_672),
.B(n_515),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_657),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_551),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_560),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_672),
.B(n_515),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_598),
.B(n_439),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_604),
.B(n_468),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_611),
.B(n_517),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_648),
.B(n_353),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_627),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_627),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_569),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_637),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_603),
.B(n_274),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_572),
.B(n_277),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_570),
.B(n_543),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_595),
.B(n_500),
.C(n_432),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_620),
.B(n_284),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_630),
.B(n_286),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_572),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_580),
.B(n_253),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_565),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_668),
.A2(n_410),
.B1(n_507),
.B2(n_454),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_682),
.B(n_429),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_637),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_615),
.B(n_311),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_605),
.B(n_329),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_632),
.B(n_289),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_632),
.B(n_291),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_631),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_689),
.B(n_298),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_556),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_621),
.B(n_300),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_668),
.B(n_308),
.Y(n_727)
);

BUFx6f_ASAP7_75t_SL g728 ( 
.A(n_557),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_674),
.B(n_294),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_644),
.Y(n_730)
);

BUFx5_ASAP7_75t_L g731 ( 
.A(n_679),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_571),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_619),
.B(n_337),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_655),
.B(n_312),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_574),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_639),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_563),
.B(n_313),
.Y(n_737)
);

NOR2x1p5_ASAP7_75t_L g738 ( 
.A(n_653),
.B(n_355),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_652),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_670),
.B(n_321),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_L g741 ( 
.A(n_655),
.B(n_322),
.Y(n_741)
);

NOR3xp33_ASAP7_75t_L g742 ( 
.A(n_575),
.B(n_365),
.C(n_364),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_649),
.B(n_325),
.Y(n_743)
);

NOR3xp33_ASAP7_75t_L g744 ( 
.A(n_608),
.B(n_384),
.C(n_376),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_639),
.Y(n_745)
);

NOR2xp67_ASAP7_75t_L g746 ( 
.A(n_612),
.B(n_507),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_562),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_623),
.B(n_328),
.Y(n_748)
);

CKINVDCx14_ASAP7_75t_R g749 ( 
.A(n_685),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_666),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_608),
.B(n_394),
.C(n_389),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_650),
.B(n_507),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_546),
.B(n_451),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_587),
.B(n_339),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_547),
.B(n_451),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_550),
.B(n_451),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_562),
.B(n_454),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_614),
.B(n_340),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_591),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_553),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_678),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_629),
.B(n_344),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_635),
.B(n_350),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_553),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_654),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_665),
.B(n_354),
.Y(n_766)
);

BUFx5_ASAP7_75t_L g767 ( 
.A(n_681),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_675),
.B(n_398),
.C(n_396),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_558),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_556),
.B(n_29),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_646),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_582),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_600),
.B(n_361),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_582),
.B(n_367),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_558),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_661),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_582),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_545),
.B(n_368),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_607),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_548),
.B(n_369),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_549),
.B(n_372),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_552),
.B(n_505),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_607),
.B(n_375),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_634),
.B(n_378),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_607),
.B(n_379),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_555),
.B(n_380),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_559),
.B(n_382),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_688),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_685),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_645),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_L g791 ( 
.A(n_626),
.B(n_597),
.C(n_642),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_661),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_561),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_554),
.B(n_610),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_610),
.A2(n_425),
.B1(n_437),
.B2(n_416),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_566),
.B(n_567),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_617),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_642),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_618),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_606),
.B(n_415),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_593),
.B(n_568),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_606),
.B(n_417),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_601),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_684),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_609),
.B(n_411),
.C(n_409),
.Y(n_805)
);

OAI221xp5_ASAP7_75t_L g806 ( 
.A1(n_676),
.A2(n_436),
.B1(n_435),
.B2(n_434),
.C(n_427),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_573),
.A2(n_261),
.B(n_272),
.C(n_285),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_616),
.B(n_418),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_576),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_577),
.B(n_423),
.Y(n_810)
);

BUFx5_ASAP7_75t_L g811 ( 
.A(n_687),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_616),
.B(n_424),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_SL g813 ( 
.A(n_579),
.B(n_443),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_585),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_581),
.B(n_583),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_680),
.B(n_30),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_583),
.B(n_505),
.Y(n_817)
);

NAND3xp33_ASAP7_75t_L g818 ( 
.A(n_609),
.B(n_443),
.C(n_493),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_584),
.B(n_505),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_690),
.B(n_584),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_690),
.B(n_622),
.Y(n_821)
);

INVx4_ASAP7_75t_L g822 ( 
.A(n_788),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_713),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_691),
.B(n_586),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_757),
.A2(n_596),
.B(n_680),
.Y(n_825)
);

BUFx8_ASAP7_75t_SL g826 ( 
.A(n_789),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_772),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_744),
.A2(n_667),
.B1(n_588),
.B2(n_599),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_779),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_777),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_753),
.A2(n_628),
.B(n_622),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_753),
.A2(n_756),
.B(n_755),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_699),
.B(n_589),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_699),
.B(n_692),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_692),
.B(n_589),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_693),
.A2(n_594),
.B(n_602),
.C(n_599),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_749),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_751),
.A2(n_663),
.B(n_658),
.C(n_677),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_809),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_779),
.B(n_601),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_694),
.B(n_667),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_SL g842 ( 
.A(n_811),
.B(n_443),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_698),
.B(n_528),
.Y(n_843)
);

NOR2xp67_ASAP7_75t_L g844 ( 
.A(n_725),
.B(n_804),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_760),
.A2(n_528),
.B(n_529),
.C(n_519),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_747),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_788),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_747),
.Y(n_848)
);

AND3x1_ASAP7_75t_SL g849 ( 
.A(n_738),
.B(n_592),
.C(n_31),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_739),
.B(n_32),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_750),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_715),
.A2(n_625),
.B(n_624),
.Y(n_852)
);

AOI21xp33_ASAP7_75t_L g853 ( 
.A1(n_816),
.A2(n_496),
.B(n_493),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_736),
.A2(n_683),
.B(n_625),
.C(n_633),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_729),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_764),
.B(n_33),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_715),
.A2(n_636),
.B(n_633),
.Y(n_857)
);

AND2x2_ASAP7_75t_SL g858 ( 
.A(n_770),
.B(n_34),
.Y(n_858)
);

NOR3xp33_ASAP7_75t_L g859 ( 
.A(n_768),
.B(n_638),
.C(n_636),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_745),
.A2(n_683),
.B(n_638),
.C(n_640),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_705),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_723),
.A2(n_641),
.B(n_640),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_702),
.B(n_35),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_728),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_717),
.B(n_36),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_720),
.B(n_38),
.Y(n_866)
);

AND2x2_ASAP7_75t_SL g867 ( 
.A(n_709),
.B(n_38),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_696),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_733),
.B(n_40),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_697),
.B(n_41),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_752),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_797),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_714),
.B(n_43),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_754),
.B(n_44),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_762),
.B(n_44),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_798),
.A2(n_518),
.B(n_521),
.C(n_520),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_795),
.A2(n_673),
.B(n_643),
.C(n_647),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_759),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_761),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_771),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_758),
.B(n_46),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_732),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_700),
.B(n_46),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_771),
.Y(n_884)
);

BUFx12f_ASAP7_75t_L g885 ( 
.A(n_799),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_735),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_700),
.B(n_48),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_815),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_701),
.B(n_48),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_723),
.A2(n_815),
.B(n_796),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_701),
.B(n_727),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_724),
.B(n_743),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_703),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_704),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_765),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_801),
.B(n_794),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_710),
.A2(n_520),
.B(n_509),
.C(n_518),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_728),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_721),
.B(n_722),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_711),
.B(n_50),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_716),
.A2(n_520),
.B(n_509),
.C(n_518),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_805),
.A2(n_651),
.B(n_664),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_718),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_774),
.B(n_50),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_SL g905 ( 
.A1(n_781),
.A2(n_656),
.B(n_662),
.C(n_660),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_695),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_712),
.B(n_52),
.Y(n_907)
);

AO21x1_ASAP7_75t_L g908 ( 
.A1(n_795),
.A2(n_659),
.B(n_499),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_763),
.B(n_55),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_810),
.A2(n_686),
.B(n_613),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_730),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_786),
.A2(n_686),
.B(n_613),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_787),
.A2(n_686),
.B(n_613),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_783),
.B(n_55),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_706),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_706),
.B(n_57),
.Y(n_916)
);

AO21x1_ASAP7_75t_L g917 ( 
.A1(n_776),
.A2(n_495),
.B(n_499),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_726),
.B(n_766),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_742),
.A2(n_58),
.B(n_59),
.C(n_62),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_793),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_817),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_737),
.Y(n_922)
);

INVx4_ASAP7_75t_L g923 ( 
.A(n_769),
.Y(n_923)
);

AOI21xp33_ASAP7_75t_L g924 ( 
.A1(n_734),
.A2(n_499),
.B(n_495),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_817),
.Y(n_925)
);

NAND2x1p5_ASAP7_75t_L g926 ( 
.A(n_708),
.B(n_495),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_741),
.A2(n_499),
.B1(n_590),
.B2(n_64),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_792),
.A2(n_59),
.B(n_63),
.C(n_64),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_778),
.B(n_63),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_780),
.B(n_65),
.Y(n_930)
);

AND2x6_ASAP7_75t_L g931 ( 
.A(n_803),
.B(n_111),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_740),
.B(n_67),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_818),
.A2(n_173),
.B(n_238),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_814),
.A2(n_748),
.B(n_707),
.Y(n_934)
);

AOI21xp33_ASAP7_75t_L g935 ( 
.A1(n_775),
.A2(n_160),
.B(n_237),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_785),
.B(n_68),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_791),
.A2(n_70),
.B1(n_71),
.B2(n_75),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_746),
.B(n_71),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_819),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_807),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_834),
.A2(n_899),
.B(n_892),
.C(n_918),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_SL g942 ( 
.A(n_842),
.B(n_813),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_880),
.Y(n_943)
);

INVxp67_ASAP7_75t_SL g944 ( 
.A(n_820),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_888),
.A2(n_782),
.B1(n_719),
.B2(n_773),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_934),
.A2(n_800),
.B(n_802),
.Y(n_946)
);

OAI21x1_ASAP7_75t_SL g947 ( 
.A1(n_833),
.A2(n_908),
.B(n_932),
.Y(n_947)
);

NOR2x1_ASAP7_75t_SL g948 ( 
.A(n_835),
.B(n_784),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_851),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_827),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_841),
.B(n_808),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_855),
.B(n_812),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_822),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_882),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_886),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_829),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_858),
.B(n_880),
.Y(n_957)
);

AO31x2_ASAP7_75t_L g958 ( 
.A1(n_917),
.A2(n_901),
.A3(n_876),
.B(n_845),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_920),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_878),
.Y(n_960)
);

NAND2xp33_ASAP7_75t_L g961 ( 
.A(n_884),
.B(n_731),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_940),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_962)
);

AOI21x1_ASAP7_75t_L g963 ( 
.A1(n_910),
.A2(n_767),
.B(n_731),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_830),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_831),
.A2(n_767),
.B(n_79),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_868),
.B(n_78),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_921),
.Y(n_967)
);

BUFx24_ASAP7_75t_L g968 ( 
.A(n_826),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_939),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_836),
.A2(n_80),
.B(n_115),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_870),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_852),
.A2(n_862),
.B(n_857),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_870),
.Y(n_973)
);

AO31x2_ASAP7_75t_L g974 ( 
.A1(n_897),
.A2(n_116),
.A3(n_124),
.B(n_125),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_919),
.A2(n_150),
.B(n_153),
.C(n_154),
.Y(n_975)
);

BUFx2_ASAP7_75t_SL g976 ( 
.A(n_864),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_823),
.B(n_828),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_SL g978 ( 
.A1(n_856),
.A2(n_186),
.B(n_187),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_912),
.A2(n_913),
.B(n_843),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_895),
.B(n_249),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_850),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_867),
.B(n_190),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_884),
.Y(n_983)
);

BUFx12f_ASAP7_75t_L g984 ( 
.A(n_837),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_922),
.B(n_205),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_853),
.A2(n_220),
.B(n_223),
.Y(n_986)
);

AOI21xp33_ASAP7_75t_L g987 ( 
.A1(n_838),
.A2(n_224),
.B(n_226),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_898),
.B(n_228),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_865),
.B(n_821),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_861),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_871),
.B(n_821),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_891),
.B(n_824),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_925),
.Y(n_993)
);

NOR3xp33_ASAP7_75t_L g994 ( 
.A(n_863),
.B(n_936),
.C(n_875),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_872),
.B(n_896),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_904),
.B(n_914),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_840),
.B(n_844),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_877),
.A2(n_900),
.B(n_907),
.C(n_873),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_883),
.A2(n_887),
.B(n_889),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_879),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_920),
.B(n_909),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_903),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_885),
.Y(n_1003)
);

OAI22x1_ASAP7_75t_L g1004 ( 
.A1(n_849),
.A2(n_926),
.B1(n_938),
.B2(n_869),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_911),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_929),
.A2(n_930),
.B(n_866),
.C(n_881),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_933),
.A2(n_902),
.B(n_860),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_933),
.A2(n_902),
.B(n_854),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_893),
.Y(n_1009)
);

AO21x1_ASAP7_75t_L g1010 ( 
.A1(n_935),
.A2(n_874),
.B(n_916),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_915),
.B(n_846),
.Y(n_1011)
);

AND2x6_ASAP7_75t_L g1012 ( 
.A(n_847),
.B(n_848),
.Y(n_1012)
);

NAND3xp33_ASAP7_75t_L g1013 ( 
.A(n_937),
.B(n_927),
.C(n_928),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_906),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_923),
.B(n_915),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_894),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_839),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_923),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_924),
.A2(n_935),
.B(n_859),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_905),
.A2(n_842),
.B(n_906),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_931),
.B(n_790),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_822),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_834),
.B(n_690),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_832),
.A2(n_825),
.B(n_890),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_832),
.A2(n_825),
.B(n_890),
.Y(n_1025)
);

OR2x6_ASAP7_75t_L g1026 ( 
.A(n_885),
.B(n_556),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_832),
.A2(n_825),
.B(n_834),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_834),
.B(n_690),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_834),
.B(n_690),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_832),
.A2(n_825),
.B(n_834),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_834),
.B(n_690),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_832),
.A2(n_825),
.B(n_834),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_832),
.A2(n_825),
.B(n_834),
.Y(n_1033)
);

AOI211x1_ASAP7_75t_L g1034 ( 
.A1(n_841),
.A2(n_834),
.B(n_892),
.C(n_768),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_SL g1035 ( 
.A(n_919),
.B(n_685),
.C(n_512),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_834),
.A2(n_820),
.B1(n_888),
.B2(n_833),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_888),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_888),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_832),
.A2(n_825),
.B(n_890),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_832),
.A2(n_825),
.B(n_834),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_834),
.B(n_779),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_832),
.A2(n_825),
.B(n_834),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_834),
.B(n_690),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_832),
.A2(n_825),
.B(n_834),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_834),
.A2(n_899),
.B(n_892),
.C(n_918),
.Y(n_1045)
);

AO31x2_ASAP7_75t_L g1046 ( 
.A1(n_825),
.A2(n_908),
.A3(n_917),
.B(n_901),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_829),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_SL g1048 ( 
.A(n_919),
.B(n_685),
.C(n_512),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_SL g1049 ( 
.A1(n_834),
.A2(n_820),
.B(n_833),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_834),
.A2(n_899),
.B(n_892),
.C(n_918),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_834),
.B(n_690),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_832),
.A2(n_825),
.B(n_834),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_834),
.B(n_690),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_832),
.A2(n_825),
.B(n_834),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_834),
.B(n_690),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_829),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_834),
.B(n_690),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_827),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_834),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_827),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_888),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_834),
.B(n_690),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_834),
.A2(n_820),
.B1(n_888),
.B2(n_833),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_822),
.Y(n_1064)
);

NOR3xp33_ASAP7_75t_L g1065 ( 
.A(n_855),
.B(n_806),
.C(n_834),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_822),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_829),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_822),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_834),
.B(n_690),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_822),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_941),
.A2(n_1050),
.B(n_1045),
.Y(n_1071)
);

OAI221xp5_ASAP7_75t_L g1072 ( 
.A1(n_1023),
.A2(n_1029),
.B1(n_1031),
.B2(n_1043),
.C(n_1057),
.Y(n_1072)
);

AO21x1_ASAP7_75t_L g1073 ( 
.A1(n_1036),
.A2(n_1063),
.B(n_970),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_1062),
.B(n_1069),
.Y(n_1074)
);

AO21x1_ASAP7_75t_L g1075 ( 
.A1(n_1036),
.A2(n_1063),
.B(n_970),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1055),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_959),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_1028),
.B(n_1051),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_959),
.B(n_953),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_SL g1080 ( 
.A1(n_1049),
.A2(n_986),
.B(n_965),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1053),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_953),
.B(n_1064),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1059),
.B(n_944),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_949),
.Y(n_1084)
);

AOI21xp33_ASAP7_75t_L g1085 ( 
.A1(n_1013),
.A2(n_975),
.B(n_947),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_954),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_993),
.B(n_1037),
.Y(n_1087)
);

NAND2x1p5_ASAP7_75t_L g1088 ( 
.A(n_1064),
.B(n_1066),
.Y(n_1088)
);

INVx5_ASAP7_75t_L g1089 ( 
.A(n_943),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_968),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1027),
.A2(n_1032),
.B(n_1030),
.Y(n_1091)
);

BUFx12f_ASAP7_75t_L g1092 ( 
.A(n_1003),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_1035),
.A2(n_1048),
.B1(n_1065),
.B2(n_994),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1038),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1061),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_1066),
.B(n_1070),
.Y(n_1096)
);

BUFx5_ASAP7_75t_L g1097 ( 
.A(n_1012),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1033),
.A2(n_1042),
.B(n_1040),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1044),
.A2(n_1054),
.B(n_1052),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_991),
.B(n_980),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_955),
.Y(n_1101)
);

OA21x2_ASAP7_75t_L g1102 ( 
.A1(n_1019),
.A2(n_1008),
.B(n_1007),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_SL g1103 ( 
.A(n_1026),
.Y(n_1103)
);

BUFx12f_ASAP7_75t_L g1104 ( 
.A(n_1026),
.Y(n_1104)
);

CKINVDCx11_ASAP7_75t_R g1105 ( 
.A(n_1026),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_965),
.A2(n_973),
.B(n_971),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_967),
.Y(n_1107)
);

AO21x2_ASAP7_75t_L g1108 ( 
.A1(n_1019),
.A2(n_1010),
.B(n_979),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_950),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_956),
.B(n_1056),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_1058),
.Y(n_1111)
);

BUFx4f_ASAP7_75t_SL g1112 ( 
.A(n_984),
.Y(n_1112)
);

AO21x2_ASAP7_75t_L g1113 ( 
.A1(n_986),
.A2(n_998),
.B(n_1006),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_1070),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1020),
.A2(n_972),
.B(n_963),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_990),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1002),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_992),
.B(n_977),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1005),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1000),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_969),
.B(n_981),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_991),
.B(n_980),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_987),
.A2(n_999),
.B(n_946),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1047),
.B(n_1067),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_SL g1125 ( 
.A1(n_948),
.A2(n_962),
.B(n_989),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_SL g1126 ( 
.A1(n_962),
.A2(n_1001),
.B(n_983),
.Y(n_1126)
);

BUFx2_ASAP7_75t_SL g1127 ( 
.A(n_1060),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_960),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1021),
.A2(n_951),
.B(n_1013),
.C(n_978),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_SL g1130 ( 
.A1(n_982),
.A2(n_996),
.B1(n_942),
.B2(n_997),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1012),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1012),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_966),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_976),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_1017),
.Y(n_1135)
);

NAND2x1_ASAP7_75t_L g1136 ( 
.A(n_1012),
.B(n_1068),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1017),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1009),
.Y(n_1138)
);

INVx8_ASAP7_75t_L g1139 ( 
.A(n_1011),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_957),
.Y(n_1140)
);

AO21x2_ASAP7_75t_L g1141 ( 
.A1(n_945),
.A2(n_1046),
.B(n_961),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1018),
.B(n_1011),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_952),
.B(n_1041),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_964),
.B(n_995),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1034),
.B(n_1016),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1022),
.A2(n_1015),
.B(n_1046),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_SL g1147 ( 
.A1(n_988),
.A2(n_978),
.B(n_1004),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_985),
.A2(n_1014),
.B(n_1046),
.C(n_974),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_958),
.B(n_974),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1062),
.B(n_1069),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1062),
.B(n_1069),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_941),
.A2(n_1050),
.B(n_1045),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_L g1153 ( 
.A(n_1035),
.B(n_1048),
.C(n_1045),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1049),
.Y(n_1154)
);

BUFx12f_ASAP7_75t_L g1155 ( 
.A(n_1003),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1049),
.Y(n_1156)
);

OA21x2_ASAP7_75t_L g1157 ( 
.A1(n_1024),
.A2(n_1039),
.B(n_1025),
.Y(n_1157)
);

NAND2x1p5_ASAP7_75t_L g1158 ( 
.A(n_1062),
.B(n_1069),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1049),
.A2(n_1063),
.B(n_1036),
.Y(n_1159)
);

BUFx2_ASAP7_75t_R g1160 ( 
.A(n_1003),
.Y(n_1160)
);

AO21x2_ASAP7_75t_L g1161 ( 
.A1(n_947),
.A2(n_1025),
.B(n_1024),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1062),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1062),
.Y(n_1163)
);

OA21x2_ASAP7_75t_L g1164 ( 
.A1(n_1024),
.A2(n_1039),
.B(n_1025),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1076),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1110),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_1154),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_1105),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1154),
.Y(n_1169)
);

INVx4_ASAP7_75t_R g1170 ( 
.A(n_1105),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1084),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1086),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1091),
.A2(n_1099),
.B(n_1098),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1072),
.A2(n_1078),
.B1(n_1150),
.B2(n_1074),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1156),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_1090),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1081),
.B(n_1072),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1101),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1116),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1117),
.Y(n_1180)
);

CKINVDCx20_ASAP7_75t_R g1181 ( 
.A(n_1090),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_1139),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1104),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1074),
.A2(n_1150),
.B1(n_1083),
.B2(n_1143),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1119),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_1134),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1094),
.B(n_1095),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1120),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1159),
.A2(n_1158),
.B1(n_1162),
.B2(n_1151),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1087),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_1124),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1139),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1153),
.A2(n_1159),
.B1(n_1075),
.B2(n_1073),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1134),
.Y(n_1194)
);

OAI222xp33_ASAP7_75t_L g1195 ( 
.A1(n_1130),
.A2(n_1151),
.B1(n_1093),
.B2(n_1140),
.C1(n_1100),
.C2(n_1122),
.Y(n_1195)
);

NOR2x1_ASAP7_75t_L g1196 ( 
.A(n_1114),
.B(n_1136),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1162),
.B(n_1121),
.Y(n_1197)
);

INVx6_ASAP7_75t_L g1198 ( 
.A(n_1139),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_1137),
.Y(n_1199)
);

INVxp33_ASAP7_75t_L g1200 ( 
.A(n_1082),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_1111),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1157),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1164),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1153),
.A2(n_1071),
.B1(n_1152),
.B2(n_1130),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1071),
.B(n_1152),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1089),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1137),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1164),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1133),
.A2(n_1125),
.B1(n_1163),
.B2(n_1106),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_1082),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1106),
.A2(n_1103),
.B1(n_1118),
.B2(n_1122),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1118),
.B(n_1144),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1107),
.Y(n_1213)
);

AOI222xp33_ASAP7_75t_L g1214 ( 
.A1(n_1103),
.A2(n_1109),
.B1(n_1112),
.B2(n_1144),
.C1(n_1111),
.C2(n_1145),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1128),
.B(n_1138),
.Y(n_1215)
);

BUFx12f_ASAP7_75t_L g1216 ( 
.A(n_1092),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1135),
.A2(n_1140),
.B1(n_1129),
.B2(n_1077),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1126),
.A2(n_1113),
.B1(n_1080),
.B2(n_1147),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1127),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1088),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1205),
.B(n_1161),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1169),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1205),
.B(n_1129),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1210),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1204),
.A2(n_1085),
.B1(n_1142),
.B2(n_1149),
.Y(n_1225)
);

NOR2x1_ASAP7_75t_L g1226 ( 
.A(n_1196),
.B(n_1206),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1187),
.B(n_1108),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1166),
.Y(n_1228)
);

NOR2x1_ASAP7_75t_L g1229 ( 
.A(n_1206),
.B(n_1114),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1197),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1206),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1204),
.A2(n_1142),
.B1(n_1149),
.B2(n_1141),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1215),
.B(n_1146),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1215),
.B(n_1102),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1190),
.B(n_1148),
.Y(n_1235)
);

INVx3_ASAP7_75t_SL g1236 ( 
.A(n_1182),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1177),
.B(n_1079),
.Y(n_1237)
);

OAI21xp33_ASAP7_75t_L g1238 ( 
.A1(n_1193),
.A2(n_1200),
.B(n_1218),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1212),
.B(n_1079),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1201),
.B(n_1186),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1184),
.A2(n_1088),
.B1(n_1096),
.B2(n_1097),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1210),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1199),
.B(n_1096),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1193),
.B(n_1123),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1167),
.B(n_1115),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1175),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1213),
.B(n_1123),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1173),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1220),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1211),
.A2(n_1131),
.B1(n_1132),
.B2(n_1097),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1207),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1221),
.B(n_1234),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1240),
.B(n_1194),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1221),
.B(n_1234),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1246),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_1242),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1222),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1236),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1227),
.B(n_1202),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1222),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1235),
.B(n_1203),
.Y(n_1261)
);

NAND3xp33_ASAP7_75t_L g1262 ( 
.A(n_1238),
.B(n_1214),
.C(n_1229),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1236),
.B(n_1200),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1247),
.B(n_1208),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1225),
.A2(n_1211),
.B1(n_1174),
.B2(n_1189),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_1228),
.Y(n_1266)
);

AND2x4_ASAP7_75t_SL g1267 ( 
.A(n_1241),
.B(n_1182),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1247),
.B(n_1173),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1231),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1235),
.B(n_1217),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1233),
.B(n_1218),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1230),
.B(n_1171),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1252),
.B(n_1244),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1258),
.B(n_1236),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1257),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1252),
.B(n_1254),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1270),
.B(n_1223),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1270),
.B(n_1223),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1252),
.B(n_1244),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1261),
.B(n_1257),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1260),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1268),
.B(n_1233),
.Y(n_1282)
);

INVxp67_ASAP7_75t_SL g1283 ( 
.A(n_1255),
.Y(n_1283)
);

INVx6_ASAP7_75t_L g1284 ( 
.A(n_1258),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1254),
.B(n_1259),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1268),
.B(n_1245),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1268),
.B(n_1248),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1264),
.B(n_1245),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1284),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1277),
.B(n_1266),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1275),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1283),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1277),
.B(n_1266),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1284),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1275),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1281),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1284),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1281),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_1280),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1283),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1278),
.B(n_1273),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1276),
.B(n_1271),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1284),
.Y(n_1303)
);

INVxp67_ASAP7_75t_L g1304 ( 
.A(n_1290),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1291),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1303),
.A2(n_1284),
.B1(n_1262),
.B2(n_1258),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1292),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1293),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1291),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1299),
.A2(n_1262),
.B1(n_1278),
.B2(n_1286),
.Y(n_1310)
);

OAI221xp5_ASAP7_75t_L g1311 ( 
.A1(n_1294),
.A2(n_1265),
.B1(n_1238),
.B2(n_1219),
.C(n_1274),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1301),
.B(n_1253),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1295),
.Y(n_1313)
);

OAI221xp5_ASAP7_75t_L g1314 ( 
.A1(n_1294),
.A2(n_1256),
.B1(n_1258),
.B2(n_1280),
.C(n_1241),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1300),
.B(n_1285),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1302),
.A2(n_1286),
.B1(n_1288),
.B2(n_1287),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1302),
.B(n_1273),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1295),
.Y(n_1318)
);

AOI21xp33_ASAP7_75t_L g1319 ( 
.A1(n_1289),
.A2(n_1256),
.B(n_1251),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1296),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1289),
.B(n_1286),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1310),
.A2(n_1286),
.B1(n_1282),
.B2(n_1279),
.Y(n_1322)
);

AOI21xp33_ASAP7_75t_L g1323 ( 
.A1(n_1311),
.A2(n_1272),
.B(n_1297),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1304),
.B(n_1273),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_SL g1325 ( 
.A(n_1306),
.B(n_1168),
.C(n_1297),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1308),
.B(n_1279),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1305),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1314),
.A2(n_1282),
.B1(n_1279),
.B2(n_1287),
.Y(n_1328)
);

AOI211xp5_ASAP7_75t_L g1329 ( 
.A1(n_1306),
.A2(n_1319),
.B(n_1303),
.C(n_1195),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1309),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1325),
.A2(n_1263),
.B(n_1321),
.Y(n_1331)
);

NOR3xp33_ASAP7_75t_L g1332 ( 
.A(n_1329),
.B(n_1183),
.C(n_1191),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1328),
.A2(n_1312),
.B1(n_1316),
.B2(n_1321),
.Y(n_1333)
);

AND4x1_ASAP7_75t_L g1334 ( 
.A(n_1322),
.B(n_1170),
.C(n_1216),
.D(n_1160),
.Y(n_1334)
);

OAI32xp33_ASAP7_75t_L g1335 ( 
.A1(n_1323),
.A2(n_1315),
.A3(n_1307),
.B1(n_1317),
.B2(n_1168),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1324),
.A2(n_1271),
.B1(n_1326),
.B2(n_1267),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1327),
.A2(n_1181),
.B(n_1176),
.Y(n_1337)
);

AOI221xp5_ASAP7_75t_L g1338 ( 
.A1(n_1330),
.A2(n_1320),
.B1(n_1313),
.B2(n_1318),
.C(n_1282),
.Y(n_1338)
);

NAND4xp25_ASAP7_75t_L g1339 ( 
.A(n_1325),
.B(n_1250),
.C(n_1232),
.D(n_1209),
.Y(n_1339)
);

O2A1O1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1325),
.A2(n_1181),
.B(n_1176),
.C(n_1243),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1336),
.B(n_1276),
.Y(n_1341)
);

NAND4xp25_ASAP7_75t_L g1342 ( 
.A(n_1340),
.B(n_1332),
.C(n_1337),
.D(n_1335),
.Y(n_1342)
);

AOI211xp5_ASAP7_75t_L g1343 ( 
.A1(n_1331),
.A2(n_1183),
.B(n_1272),
.C(n_1237),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1333),
.Y(n_1344)
);

NAND4xp75_ASAP7_75t_L g1345 ( 
.A(n_1338),
.B(n_1229),
.C(n_1226),
.D(n_1160),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1334),
.B(n_1282),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1339),
.B(n_1296),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1337),
.Y(n_1348)
);

NAND3xp33_ASAP7_75t_L g1349 ( 
.A(n_1344),
.B(n_1209),
.C(n_1178),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1347),
.B(n_1285),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1347),
.Y(n_1351)
);

OA22x2_ASAP7_75t_L g1352 ( 
.A1(n_1348),
.A2(n_1267),
.B1(n_1269),
.B2(n_1182),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_SL g1353 ( 
.A(n_1342),
.B(n_1216),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1341),
.B(n_1298),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1346),
.Y(n_1355)
);

NAND2xp33_ASAP7_75t_L g1356 ( 
.A(n_1355),
.B(n_1345),
.Y(n_1356)
);

NOR2x1_ASAP7_75t_L g1357 ( 
.A(n_1353),
.B(n_1112),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1351),
.B(n_1343),
.Y(n_1358)
);

NAND4xp25_ASAP7_75t_L g1359 ( 
.A(n_1349),
.B(n_1243),
.C(n_1249),
.D(n_1239),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1350),
.B(n_1287),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1354),
.Y(n_1361)
);

NOR2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1352),
.B(n_1155),
.Y(n_1362)
);

NOR3x1_ASAP7_75t_L g1363 ( 
.A(n_1355),
.B(n_1192),
.C(n_1224),
.Y(n_1363)
);

NOR2x1_ASAP7_75t_L g1364 ( 
.A(n_1357),
.B(n_1249),
.Y(n_1364)
);

NAND4xp75_ASAP7_75t_L g1365 ( 
.A(n_1363),
.B(n_1192),
.C(n_1226),
.D(n_1165),
.Y(n_1365)
);

NAND2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1362),
.B(n_1249),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1364),
.Y(n_1367)
);

AO22x1_ASAP7_75t_L g1368 ( 
.A1(n_1365),
.A2(n_1358),
.B1(n_1361),
.B2(n_1356),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1366),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1368),
.B(n_1359),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1369),
.A2(n_1360),
.B1(n_1198),
.B2(n_1267),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_1370),
.Y(n_1372)
);

XNOR2xp5_ASAP7_75t_L g1373 ( 
.A(n_1371),
.B(n_1367),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1370),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1373),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1372),
.Y(n_1376)
);

AOI21xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1374),
.A2(n_1224),
.B(n_1179),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1375),
.A2(n_1198),
.B1(n_1185),
.B2(n_1180),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_SL g1379 ( 
.A1(n_1378),
.A2(n_1377),
.B(n_1376),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1379),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1380),
.A2(n_1172),
.B(n_1188),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1381),
.A2(n_1380),
.B1(n_1198),
.B2(n_1231),
.Y(n_1382)
);


endmodule