module real_jpeg_25414_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_258;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_1),
.A2(n_67),
.B1(n_68),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_74),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_2),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_3),
.A2(n_27),
.B1(n_39),
.B2(n_42),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_3),
.A2(n_27),
.B1(n_51),
.B2(n_52),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_3),
.A2(n_27),
.B1(n_67),
.B2(n_68),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_5),
.A2(n_51),
.B1(n_52),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_5),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_5),
.A2(n_67),
.B1(n_68),
.B2(n_87),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_5),
.A2(n_39),
.B1(n_42),
.B2(n_87),
.Y(n_136)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_7),
.A2(n_67),
.B1(n_68),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_7),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_9),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_9),
.A2(n_51),
.B1(n_52),
.B2(n_66),
.Y(n_94)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_11),
.A2(n_31),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_11),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_11),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_11),
.A2(n_44),
.B1(n_67),
.B2(n_68),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_12),
.A2(n_39),
.B1(n_42),
.B2(n_58),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_12),
.A2(n_36),
.B1(n_58),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_12),
.A2(n_51),
.B1(n_52),
.B2(n_58),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_12),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_13),
.B(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_13),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_13),
.B(n_38),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_13),
.B(n_52),
.C(n_54),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_13),
.A2(n_39),
.B1(n_42),
.B2(n_161),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_13),
.B(n_110),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_13),
.A2(n_51),
.B1(n_52),
.B2(n_161),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_13),
.B(n_67),
.C(n_82),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_13),
.A2(n_69),
.B(n_221),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_15),
.A2(n_39),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_15),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_15),
.A2(n_49),
.B1(n_67),
.B2(n_68),
.Y(n_170)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_16),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_16),
.B(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_16),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_146),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_144),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_20),
.B(n_121),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_88),
.C(n_98),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_21),
.A2(n_22),
.B1(n_88),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_62),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_46),
.B2(n_47),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_25),
.B(n_46),
.C(n_62),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_38),
.B2(n_43),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_26),
.Y(n_100)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g112 ( 
.A1(n_31),
.A2(n_35),
.A3(n_42),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_31),
.A2(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_32),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_32),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_32),
.A2(n_141),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_42),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g115 ( 
.A(n_34),
.B(n_39),
.Y(n_115)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_37),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_37),
.B(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_42),
.B1(n_54),
.B2(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_39),
.B(n_187),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_43),
.Y(n_138)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B(n_56),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_48),
.A2(n_50),
.B1(n_60),
.B2(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_50),
.A2(n_56),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_52),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_52),
.B(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_57),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_59),
.A2(n_108),
.B1(n_110),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_60),
.A2(n_107),
.B(n_109),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_60),
.A2(n_109),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_78),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_63),
.B(n_78),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_73),
.B2(n_75),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_65),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_116)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_70),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_68),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_68),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_73),
.B1(n_75),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_90),
.B(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_69),
.A2(n_119),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_69),
.B(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_69),
.A2(n_220),
.B(n_221),
.Y(n_219)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_77),
.B(n_161),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_79),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_79),
.A2(n_209),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_80),
.A2(n_94),
.B1(n_95),
.B2(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_80),
.B(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_80),
.A2(n_95),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_84),
.A2(n_85),
.B(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_84),
.A2(n_157),
.B(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_84),
.B(n_161),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_88),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_95),
.B(n_158),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_98),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_106),
.C(n_111),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_99),
.B(n_106),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_111),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_112),
.B(n_116),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_117),
.A2(n_232),
.B1(n_234),
.B2(n_236),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_120),
.A2(n_189),
.B(n_190),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_143),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_131),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_142),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B(n_140),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_179),
.B(n_264),
.C(n_269),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_173),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_163),
.C(n_164),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_149),
.A2(n_150),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_159),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_155),
.C(n_159),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_154),
.Y(n_166)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_163),
.B(n_164),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_169),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_174),
.B(n_177),
.C(n_178),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_258),
.B(n_263),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_210),
.B(n_257),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_199),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_184),
.B(n_199),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.C(n_196),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_185),
.B(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_192),
.A2(n_196),
.B1(n_197),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_195),
.Y(n_208)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_200),
.B(n_206),
.C(n_207),
.Y(n_262)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_251),
.B(n_256),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_229),
.B(n_250),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_223),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_223),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_219),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_218),
.C(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_220),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_227),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_239),
.B(n_249),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_237),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_237),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_233),
.A2(n_235),
.B(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_244),
.B(n_248),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_242),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_255),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_262),
.Y(n_263)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);


endmodule