module fake_jpeg_18818_n_254 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_254);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_13;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_14),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_10),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_17),
.B1(n_19),
.B2(n_11),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_17),
.B1(n_30),
.B2(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_27),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_52),
.B1(n_57),
.B2(n_17),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_55),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_31),
.B(n_20),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_54),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_30),
.B(n_26),
.C(n_24),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_33),
.B1(n_42),
.B2(n_25),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_42),
.B1(n_38),
.B2(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_43),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_25),
.C(n_42),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_57),
.C(n_46),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_57),
.B1(n_53),
.B2(n_52),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_70),
.B1(n_65),
.B2(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_88),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_61),
.B1(n_59),
.B2(n_55),
.Y(n_94)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_49),
.C(n_57),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_90),
.B(n_75),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_104),
.B1(n_25),
.B2(n_46),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_108),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_99),
.A2(n_100),
.B(n_109),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_64),
.B(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_61),
.B1(n_70),
.B2(n_74),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_74),
.B(n_67),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_11),
.B(n_15),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_107),
.A2(n_85),
.B1(n_59),
.B2(n_46),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_90),
.B(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_31),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_88),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_20),
.C(n_16),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_81),
.C(n_86),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_120),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_126),
.B1(n_39),
.B2(n_41),
.Y(n_153)
);

CKINVDCx12_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_46),
.C(n_82),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_82),
.B1(n_68),
.B2(n_66),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_124),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_82),
.B1(n_66),
.B2(n_92),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_28),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_130),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_66),
.B1(n_59),
.B2(n_51),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_102),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_92),
.Y(n_129)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

OA21x2_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_23),
.B(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_73),
.Y(n_132)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_136),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_19),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_135),
.B(n_137),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_39),
.C(n_24),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_19),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_130),
.B(n_111),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_144),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_102),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_149),
.B(n_157),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_133),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_19),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_161),
.B1(n_124),
.B2(n_118),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_34),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_158),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_39),
.B1(n_17),
.B2(n_58),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_159),
.B1(n_136),
.B2(n_17),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_115),
.B(n_11),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_41),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_17),
.B1(n_58),
.B2(n_50),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_41),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_166),
.B1(n_172),
.B2(n_177),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_114),
.C(n_134),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_173),
.C(n_179),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_134),
.B1(n_138),
.B2(n_121),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_125),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_159),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_138),
.B(n_121),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_21),
.B(n_15),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_126),
.C(n_50),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_178),
.Y(n_193)
);

FAx1_ASAP7_75t_SL g175 ( 
.A(n_160),
.B(n_20),
.CI(n_21),
.CON(n_175),
.SN(n_175)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_154),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_15),
.B(n_21),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_147),
.A2(n_58),
.B1(n_41),
.B2(n_47),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_22),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_26),
.C(n_24),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_141),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_181),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_165),
.B(n_170),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_187),
.C(n_18),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_147),
.B1(n_162),
.B2(n_161),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_186),
.Y(n_200)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_164),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_156),
.C(n_153),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_180),
.A2(n_158),
.B1(n_155),
.B2(n_162),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_142),
.B1(n_26),
.B2(n_3),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_178),
.B1(n_169),
.B2(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_181),
.B(n_174),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_175),
.B(n_179),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_204),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_175),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_189),
.A2(n_0),
.B(n_1),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_185),
.B(n_193),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_207),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_185),
.C(n_182),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_196),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_190),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_213),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_193),
.C(n_23),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_221),
.C(n_210),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_208),
.B(n_21),
.Y(n_215)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_201),
.C(n_209),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_1),
.B(n_3),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_23),
.C(n_22),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_222)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_228),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_200),
.C(n_199),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_218),
.C(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_216),
.A2(n_13),
.B1(n_12),
.B2(n_22),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_1),
.B(n_3),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_13),
.B1(n_12),
.B2(n_6),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_236),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_22),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_235),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_16),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_4),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_227),
.B1(n_231),
.B2(n_13),
.Y(n_240)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_16),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_4),
.C2(n_9),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_244),
.C(n_12),
.Y(n_247)
);

AOI21x1_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_232),
.B(n_234),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_241),
.B(n_6),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_4),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_16),
.C2(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_249),
.B(n_7),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_4),
.B(n_7),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_8),
.B(n_9),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_253),
.A2(n_8),
.B(n_251),
.Y(n_254)
);


endmodule