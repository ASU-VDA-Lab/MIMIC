module fake_aes_12661_n_732 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_732);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_732;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g100 ( .A(n_84), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_20), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_98), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_8), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_16), .B(n_94), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_11), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_87), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_73), .Y(n_107) );
BUFx5_ASAP7_75t_L g108 ( .A(n_40), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_96), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_27), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_74), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_81), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_61), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_57), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_44), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_55), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_95), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_92), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_25), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_3), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_12), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_80), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_68), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_54), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_83), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_58), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_53), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_28), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_49), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_43), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_78), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_36), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_91), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_64), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_29), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_66), .Y(n_136) );
INVx1_ASAP7_75t_SL g137 ( .A(n_46), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_19), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_6), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_108), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_100), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_120), .B(n_111), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_100), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_122), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_110), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_112), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_122), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_112), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_120), .B(n_0), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_138), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_108), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_113), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_139), .Y(n_154) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_113), .A2(n_39), .B(n_97), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_111), .B(n_0), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_139), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_114), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_103), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_158), .B(n_116), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_158), .B(n_126), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_143), .A2(n_121), .B1(n_103), .B2(n_101), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_145), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_158), .B(n_102), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_145), .Y(n_165) );
AND3x2_ASAP7_75t_L g166 ( .A(n_142), .B(n_130), .C(n_106), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_154), .B(n_107), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_140), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_157), .Y(n_169) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_158), .B(n_104), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_152), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
INVx2_ASAP7_75t_SL g175 ( .A(n_143), .Y(n_175) );
INVxp67_ASAP7_75t_SL g176 ( .A(n_146), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_145), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_146), .B(n_109), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
NAND2x1_ASAP7_75t_L g180 ( .A(n_157), .B(n_115), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_147), .A2(n_138), .B1(n_105), .B2(n_127), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_147), .B(n_119), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_145), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_149), .B(n_114), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_145), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_148), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_148), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_176), .A2(n_153), .B1(n_149), .B2(n_156), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_176), .A2(n_153), .B1(n_150), .B2(n_117), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_184), .B(n_117), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_184), .A2(n_141), .B1(n_144), .B2(n_148), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_169), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_169), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_184), .B(n_118), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_182), .B(n_159), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_175), .B(n_118), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_169), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_160), .B(n_125), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_161), .B(n_125), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_170), .B(n_129), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_170), .A2(n_134), .B1(n_129), .B2(n_131), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_169), .Y(n_205) );
NAND2xp33_ASAP7_75t_SL g206 ( .A(n_180), .B(n_131), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_182), .A2(n_141), .B1(n_144), .B2(n_148), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_182), .A2(n_141), .B1(n_144), .B2(n_148), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_180), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_175), .B(n_134), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_179), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_179), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_179), .Y(n_213) );
NOR2x1p5_ASAP7_75t_L g214 ( .A(n_167), .B(n_136), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_175), .B(n_136), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_170), .B(n_159), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_182), .B(n_167), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_178), .B(n_155), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_164), .B(n_137), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_178), .B(n_123), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_166), .B(n_124), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_162), .A2(n_133), .B1(n_135), .B2(n_128), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_179), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_166), .B(n_162), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_181), .A2(n_132), .B1(n_144), .B2(n_141), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_189), .B(n_141), .Y(n_226) );
NOR2x2_ASAP7_75t_L g227 ( .A(n_174), .B(n_155), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_189), .B(n_141), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_189), .B(n_144), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_189), .A2(n_144), .B1(n_108), .B2(n_3), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_168), .A2(n_108), .B1(n_2), .B2(n_4), .Y(n_231) );
INVx3_ASAP7_75t_SL g232 ( .A(n_227), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_217), .B(n_168), .Y(n_233) );
CKINVDCx11_ASAP7_75t_R g234 ( .A(n_191), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_218), .A2(n_171), .B(n_172), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_193), .B(n_174), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_191), .B(n_171), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_218), .A2(n_172), .B(n_173), .C(n_177), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_192), .B(n_173), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_203), .A2(n_108), .B1(n_190), .B2(n_177), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_198), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_199), .B(n_108), .Y(n_242) );
INVxp67_ASAP7_75t_L g243 ( .A(n_197), .Y(n_243) );
NOR2x1_ASAP7_75t_L g244 ( .A(n_214), .B(n_183), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_195), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_192), .A2(n_190), .B1(n_183), .B2(n_186), .Y(n_246) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_228), .A2(n_188), .B(n_187), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_198), .B(n_108), .Y(n_248) );
NOR2xp33_ASAP7_75t_SL g249 ( .A(n_224), .B(n_108), .Y(n_249) );
AO32x2_ASAP7_75t_L g250 ( .A1(n_209), .A2(n_188), .A3(n_187), .B1(n_185), .B2(n_165), .Y(n_250) );
INVx4_ASAP7_75t_L g251 ( .A(n_195), .Y(n_251) );
INVx2_ASAP7_75t_SL g252 ( .A(n_214), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_204), .B(n_1), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_196), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_220), .A2(n_186), .B(n_187), .C(n_188), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_199), .A2(n_185), .B(n_165), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_216), .A2(n_185), .B(n_165), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_205), .A2(n_163), .B(n_41), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_SL g259 ( .A1(n_229), .A2(n_163), .B(n_42), .C(n_45), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_201), .A2(n_163), .B(n_2), .C(n_4), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_202), .A2(n_1), .B(n_5), .C(n_6), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_205), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_204), .B(n_5), .Y(n_263) );
NOR2x1_ASAP7_75t_L g264 ( .A(n_221), .B(n_7), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_212), .Y(n_265) );
BUFx2_ASAP7_75t_R g266 ( .A(n_232), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_235), .A2(n_230), .B(n_225), .C(n_231), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_262), .Y(n_268) );
AO31x2_ASAP7_75t_L g269 ( .A1(n_238), .A2(n_226), .A3(n_212), .B(n_196), .Y(n_269) );
CKINVDCx11_ASAP7_75t_R g270 ( .A(n_234), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_235), .A2(n_230), .B(n_225), .C(n_222), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_236), .A2(n_210), .B1(n_215), .B2(n_206), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_247), .A2(n_194), .B(n_223), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_256), .A2(n_223), .B(n_200), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_256), .A2(n_200), .B(n_213), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_241), .B(n_222), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_243), .B(n_219), .Y(n_277) );
AOI21x1_ASAP7_75t_L g278 ( .A1(n_258), .A2(n_213), .B(n_211), .Y(n_278) );
BUFx12f_ASAP7_75t_L g279 ( .A(n_252), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_239), .B(n_209), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_233), .A2(n_211), .B1(n_208), .B2(n_207), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_248), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_258), .A2(n_48), .B(n_93), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_253), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_254), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_257), .A2(n_50), .B(n_90), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_257), .A2(n_242), .B(n_237), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_263), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_276), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_288), .B(n_265), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_278), .A2(n_255), .B(n_264), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_277), .A2(n_244), .B1(n_246), .B2(n_251), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_268), .Y(n_293) );
AO31x2_ASAP7_75t_L g294 ( .A1(n_271), .A2(n_260), .A3(n_261), .B(n_251), .Y(n_294) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_287), .A2(n_259), .B(n_255), .Y(n_295) );
NOR3xp33_ASAP7_75t_L g296 ( .A(n_277), .B(n_245), .C(n_249), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_268), .B(n_254), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_274), .A2(n_275), .B(n_267), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_282), .Y(n_299) );
AO31x2_ASAP7_75t_L g300 ( .A1(n_271), .A2(n_250), .A3(n_240), .B(n_254), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_273), .Y(n_301) );
INVx2_ASAP7_75t_SL g302 ( .A(n_285), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_280), .B(n_250), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
AO31x2_ASAP7_75t_L g306 ( .A1(n_267), .A2(n_250), .A3(n_10), .B(n_11), .Y(n_306) );
AOI21xp33_ASAP7_75t_SL g307 ( .A1(n_284), .A2(n_9), .B(n_10), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_269), .Y(n_308) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_283), .A2(n_51), .B(n_89), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_269), .Y(n_310) );
NAND2x1p5_ASAP7_75t_L g311 ( .A(n_286), .B(n_47), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_293), .B(n_269), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_293), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_298), .A2(n_281), .B(n_272), .Y(n_314) );
OA21x2_ASAP7_75t_L g315 ( .A1(n_298), .A2(n_56), .B(n_99), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_293), .B(n_12), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_301), .Y(n_317) );
AO21x2_ASAP7_75t_L g318 ( .A1(n_301), .A2(n_13), .B(n_14), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_301), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_305), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_305), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_308), .B(n_13), .Y(n_322) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_291), .A2(n_59), .B(n_88), .Y(n_323) );
NAND3xp33_ASAP7_75t_L g324 ( .A(n_307), .B(n_270), .C(n_266), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_297), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_297), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_303), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_299), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_299), .B(n_279), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_306), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_306), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_300), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_308), .B(n_14), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_306), .Y(n_335) );
NOR2xp67_ASAP7_75t_SL g336 ( .A(n_309), .B(n_279), .Y(n_336) );
INVxp67_ASAP7_75t_L g337 ( .A(n_289), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_310), .B(n_15), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_310), .B(n_15), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_300), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_306), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_306), .B(n_16), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_306), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_300), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_327), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_312), .B(n_306), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_320), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_324), .A2(n_296), .B1(n_292), .B2(n_290), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_320), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_312), .B(n_300), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_312), .B(n_300), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_324), .A2(n_296), .B1(n_290), .B2(n_303), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_337), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_332), .B(n_300), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_333), .B(n_300), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_327), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_328), .B(n_304), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_333), .B(n_304), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_317), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_333), .B(n_294), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_328), .B(n_294), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_327), .Y(n_362) );
INVx3_ASAP7_75t_L g363 ( .A(n_317), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_333), .B(n_294), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_313), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_332), .B(n_294), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_313), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_317), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_319), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_326), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_333), .B(n_294), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_340), .B(n_294), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_319), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_321), .B(n_302), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_340), .B(n_291), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_340), .B(n_291), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_344), .B(n_295), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_316), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_344), .B(n_321), .Y(n_379) );
INVx4_ASAP7_75t_L g380 ( .A(n_316), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_321), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_344), .B(n_295), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_342), .A2(n_302), .B1(n_295), .B2(n_309), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_325), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_319), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_330), .Y(n_386) );
INVx4_ASAP7_75t_R g387 ( .A(n_322), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_326), .B(n_295), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_325), .B(n_302), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_330), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_331), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_326), .B(n_62), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_331), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_335), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_323), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_335), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_323), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_341), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_326), .B(n_307), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_358), .B(n_343), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_358), .B(n_343), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_358), .B(n_341), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_353), .B(n_339), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_365), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_350), .B(n_342), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_350), .B(n_351), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_365), .B(n_339), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_350), .B(n_342), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_366), .B(n_339), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_359), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_367), .Y(n_411) );
INVxp33_ASAP7_75t_L g412 ( .A(n_345), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_366), .B(n_338), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_359), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_351), .B(n_326), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_351), .B(n_338), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_357), .B(n_338), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_348), .B(n_329), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_367), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_360), .B(n_334), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_345), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_347), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_356), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_347), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_360), .B(n_322), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_349), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_360), .B(n_322), .Y(n_428) );
NOR2xp33_ASAP7_75t_R g429 ( .A(n_387), .B(n_329), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_364), .B(n_334), .Y(n_430) );
AND2x4_ASAP7_75t_SL g431 ( .A(n_380), .B(n_334), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_349), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_356), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_381), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_357), .B(n_316), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_359), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_364), .B(n_314), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_381), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_364), .B(n_314), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_346), .B(n_318), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_371), .B(n_314), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_371), .B(n_318), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_371), .B(n_318), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_346), .B(n_318), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g445 ( .A(n_392), .B(n_336), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_346), .B(n_323), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_379), .B(n_336), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_386), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_355), .B(n_323), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_380), .A2(n_323), .B1(n_315), .B2(n_309), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_355), .B(n_315), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_354), .B(n_315), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_379), .B(n_17), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_379), .B(n_17), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_386), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_352), .B(n_18), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_391), .Y(n_457) );
NAND2x1p5_ASAP7_75t_L g458 ( .A(n_392), .B(n_315), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_355), .B(n_315), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_372), .B(n_18), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_391), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_372), .B(n_309), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_372), .B(n_309), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_375), .B(n_19), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_394), .B(n_311), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_394), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_374), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_375), .B(n_311), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_396), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_362), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_396), .B(n_311), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_375), .B(n_311), .Y(n_472) );
INVx4_ASAP7_75t_L g473 ( .A(n_392), .Y(n_473) );
NOR2xp67_ASAP7_75t_SL g474 ( .A(n_380), .B(n_21), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_376), .B(n_22), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_368), .Y(n_476) );
NOR2xp67_ASAP7_75t_L g477 ( .A(n_362), .B(n_23), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_384), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_361), .B(n_24), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_406), .B(n_370), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_406), .B(n_370), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_409), .B(n_374), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_415), .B(n_370), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_400), .B(n_361), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_415), .B(n_384), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_416), .B(n_380), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_448), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_467), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_409), .B(n_378), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_404), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_413), .B(n_378), .Y(n_491) );
NAND2x1_ASAP7_75t_SL g492 ( .A(n_473), .B(n_392), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_413), .B(n_398), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_416), .B(n_398), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_473), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_400), .B(n_390), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_426), .B(n_390), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_467), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_401), .B(n_390), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_455), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_478), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_401), .B(n_393), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_457), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_402), .B(n_393), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_461), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_426), .B(n_428), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_466), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_478), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_424), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_402), .B(n_393), .Y(n_510) );
AOI31xp33_ASAP7_75t_L g511 ( .A1(n_445), .A2(n_387), .A3(n_383), .B(n_399), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_469), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_428), .B(n_376), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_430), .B(n_376), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_405), .B(n_377), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_419), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_430), .B(n_389), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_423), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_425), .Y(n_519) );
INVxp67_ASAP7_75t_L g520 ( .A(n_422), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_421), .B(n_389), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_407), .B(n_363), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_405), .B(n_382), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_408), .B(n_382), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_424), .B(n_473), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_431), .B(n_388), .Y(n_526) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_477), .B(n_392), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_427), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_408), .B(n_432), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_421), .B(n_431), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_445), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_434), .B(n_382), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_464), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_438), .Y(n_534) );
NAND4xp75_ASAP7_75t_L g535 ( .A(n_464), .B(n_399), .C(n_377), .D(n_385), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_444), .B(n_388), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_407), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_403), .B(n_373), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_443), .B(n_388), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_470), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_433), .Y(n_541) );
NAND2x1p5_ASAP7_75t_L g542 ( .A(n_474), .B(n_373), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_421), .B(n_388), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_437), .B(n_388), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_470), .Y(n_545) );
OAI33xp33_ASAP7_75t_L g546 ( .A1(n_460), .A2(n_385), .A3(n_369), .B1(n_368), .B2(n_395), .B3(n_397), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_411), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_417), .B(n_373), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_418), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_443), .B(n_385), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_412), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_420), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_437), .B(n_441), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_435), .B(n_373), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_439), .B(n_441), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_439), .B(n_363), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_453), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_440), .B(n_369), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_454), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_475), .B(n_363), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_442), .B(n_363), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_410), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_414), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_475), .B(n_369), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_412), .B(n_397), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_429), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_414), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_442), .B(n_397), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_490), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_487), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_540), .Y(n_571) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_516), .A2(n_456), .B(n_479), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_555), .B(n_442), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_551), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_556), .Y(n_575) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_520), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_533), .A2(n_566), .B1(n_511), .B2(n_535), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_500), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_566), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_501), .Y(n_580) );
AOI221xp5_ASAP7_75t_SL g581 ( .A1(n_511), .A2(n_447), .B1(n_446), .B2(n_451), .C(n_459), .Y(n_581) );
NOR2x1p5_ASAP7_75t_L g582 ( .A(n_531), .B(n_452), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_503), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_505), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_507), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_529), .B(n_452), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_512), .Y(n_587) );
INVx2_ASAP7_75t_SL g588 ( .A(n_509), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_537), .B(n_459), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_529), .B(n_436), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_553), .B(n_472), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_506), .B(n_472), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_508), .Y(n_593) );
AOI21xp33_ASAP7_75t_L g594 ( .A1(n_557), .A2(n_479), .B(n_465), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_525), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_513), .B(n_468), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_518), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_541), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_519), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_545), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_515), .B(n_476), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_528), .Y(n_602) );
NOR3xp33_ASAP7_75t_L g603 ( .A(n_559), .B(n_471), .C(n_395), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_514), .B(n_468), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_534), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_484), .B(n_451), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_547), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_515), .B(n_476), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_523), .B(n_436), .Y(n_609) );
INVxp67_ASAP7_75t_L g610 ( .A(n_488), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_549), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_562), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_563), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_484), .B(n_449), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_485), .B(n_462), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_498), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_525), .B(n_458), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_552), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_493), .Y(n_619) );
NAND2x1_ASAP7_75t_L g620 ( .A(n_495), .B(n_450), .Y(n_620) );
INVx2_ASAP7_75t_SL g621 ( .A(n_530), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_567), .Y(n_622) );
NAND2x1p5_ASAP7_75t_L g623 ( .A(n_527), .B(n_531), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_489), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_496), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_494), .B(n_449), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_491), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_523), .B(n_446), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_524), .B(n_463), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_542), .A2(n_458), .B(n_397), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_522), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_499), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_502), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_521), .B(n_463), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_524), .B(n_462), .Y(n_635) );
INVx2_ASAP7_75t_SL g636 ( .A(n_482), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_502), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_581), .A2(n_568), .B1(n_495), .B2(n_542), .C(n_492), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_581), .A2(n_486), .B1(n_543), .B2(n_561), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_570), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_578), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_579), .B(n_504), .Y(n_642) );
XNOR2xp5_ASAP7_75t_L g643 ( .A(n_588), .B(n_480), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_625), .B(n_517), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_579), .B(n_504), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_582), .A2(n_526), .B1(n_561), .B2(n_568), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g647 ( .A1(n_577), .A2(n_526), .B(n_481), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_583), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_586), .B(n_536), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_571), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_576), .Y(n_651) );
OA22x2_ASAP7_75t_L g652 ( .A1(n_595), .A2(n_510), .B1(n_497), .B2(n_483), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_584), .Y(n_653) );
OAI332xp33_ASAP7_75t_L g654 ( .A1(n_577), .A2(n_550), .A3(n_539), .B1(n_538), .B2(n_532), .B3(n_558), .C1(n_548), .C2(n_554), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_585), .Y(n_655) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_574), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_617), .A2(n_546), .B(n_558), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_587), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_597), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_623), .B(n_564), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_569), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_599), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_602), .Y(n_663) );
AOI21xp33_ASAP7_75t_L g664 ( .A1(n_620), .A2(n_565), .B(n_532), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_623), .A2(n_560), .B(n_544), .Y(n_665) );
NOR2xp67_ASAP7_75t_L g666 ( .A(n_621), .B(n_630), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_630), .B(n_550), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_605), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_612), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_632), .B(n_395), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_600), .Y(n_671) );
INVx1_ASAP7_75t_SL g672 ( .A(n_636), .Y(n_672) );
OAI321xp33_ASAP7_75t_L g673 ( .A1(n_610), .A2(n_395), .A3(n_30), .B1(n_31), .B2(n_32), .C(n_33), .Y(n_673) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_598), .A2(n_26), .B(n_34), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g675 ( .A1(n_572), .A2(n_35), .B(n_37), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_633), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_603), .A2(n_38), .B(n_52), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_647), .A2(n_572), .B(n_616), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_657), .B(n_600), .Y(n_679) );
OAI31xp33_ASAP7_75t_L g680 ( .A1(n_647), .A2(n_627), .A3(n_624), .B(n_619), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_652), .A2(n_637), .B1(n_626), .B2(n_589), .Y(n_681) );
INVxp67_ASAP7_75t_L g682 ( .A(n_656), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_654), .B(n_606), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_654), .B(n_606), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_664), .A2(n_594), .B1(n_607), .B2(n_611), .C(n_618), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_671), .B(n_614), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_666), .B(n_592), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_652), .A2(n_573), .B1(n_628), .B2(n_635), .Y(n_688) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_665), .A2(n_628), .B1(n_629), .B2(n_614), .Y(n_689) );
NAND3xp33_ASAP7_75t_SL g690 ( .A(n_665), .B(n_590), .C(n_629), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_660), .A2(n_594), .B(n_589), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_646), .A2(n_591), .B1(n_609), .B2(n_608), .Y(n_692) );
OAI21xp5_ASAP7_75t_L g693 ( .A1(n_651), .A2(n_580), .B(n_593), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_638), .A2(n_622), .B(n_613), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_639), .B(n_634), .Y(n_695) );
OAI222xp33_ASAP7_75t_L g696 ( .A1(n_672), .A2(n_601), .B1(n_575), .B2(n_631), .C1(n_604), .C2(n_596), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_676), .Y(n_697) );
INVxp67_ASAP7_75t_L g698 ( .A(n_642), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g699 ( .A1(n_661), .A2(n_615), .B(n_63), .C(n_65), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_645), .A2(n_60), .B1(n_67), .B2(n_69), .C(n_70), .Y(n_700) );
AOI22x1_ASAP7_75t_L g701 ( .A1(n_643), .A2(n_71), .B1(n_72), .B2(n_75), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_649), .A2(n_76), .B1(n_77), .B2(n_79), .Y(n_702) );
OAI21xp5_ASAP7_75t_SL g703 ( .A1(n_675), .A2(n_82), .B(n_85), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_L g704 ( .A1(n_640), .A2(n_86), .B(n_641), .C(n_668), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g705 ( .A1(n_667), .A2(n_677), .B(n_673), .C(n_674), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_648), .Y(n_706) );
AOI211xp5_ASAP7_75t_L g707 ( .A1(n_667), .A2(n_670), .B(n_659), .C(n_653), .Y(n_707) );
AND3x4_ASAP7_75t_L g708 ( .A(n_650), .B(n_669), .C(n_644), .Y(n_708) );
OAI21xp5_ASAP7_75t_SL g709 ( .A1(n_655), .A2(n_658), .B(n_662), .Y(n_709) );
NAND4xp25_ASAP7_75t_L g710 ( .A(n_663), .B(n_647), .C(n_577), .D(n_581), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_697), .Y(n_711) );
NOR2x1_ASAP7_75t_L g712 ( .A(n_708), .B(n_710), .Y(n_712) );
OAI211xp5_ASAP7_75t_L g713 ( .A1(n_680), .A2(n_678), .B(n_705), .C(n_679), .Y(n_713) );
AOI322xp5_ASAP7_75t_L g714 ( .A1(n_684), .A2(n_683), .A3(n_689), .B1(n_690), .B2(n_695), .C1(n_698), .C2(n_682), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_706), .Y(n_715) );
AND4x1_ASAP7_75t_L g716 ( .A(n_678), .B(n_694), .C(n_704), .D(n_685), .Y(n_716) );
NOR2x1_ASAP7_75t_L g717 ( .A(n_712), .B(n_703), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g718 ( .A(n_713), .B(n_700), .C(n_699), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_716), .B(n_709), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_714), .B(n_691), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_717), .B(n_702), .C(n_688), .Y(n_721) );
AND3x4_ASAP7_75t_L g722 ( .A(n_718), .B(n_687), .C(n_696), .Y(n_722) );
NAND3xp33_ASAP7_75t_SL g723 ( .A(n_720), .B(n_681), .C(n_707), .Y(n_723) );
XNOR2xp5_ASAP7_75t_L g724 ( .A(n_722), .B(n_701), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_723), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_725), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_724), .B(n_719), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_727), .A2(n_721), .B1(n_715), .B2(n_711), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_728), .Y(n_729) );
OA21x2_ASAP7_75t_L g730 ( .A1(n_729), .A2(n_726), .B(n_711), .Y(n_730) );
XOR2xp5_ASAP7_75t_L g731 ( .A(n_730), .B(n_692), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_731), .A2(n_687), .B1(n_686), .B2(n_693), .Y(n_732) );
endmodule