module real_jpeg_29454_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_312, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_312;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_0),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_66),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_0),
.A2(n_48),
.B1(n_51),
.B2(n_66),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_66),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_1),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_1),
.A2(n_48),
.B1(n_51),
.B2(n_160),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_160),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_160),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_2),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_28),
.B1(n_63),
.B2(n_64),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_2),
.A2(n_28),
.B1(n_48),
.B2(n_51),
.Y(n_236)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_4),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_4),
.A2(n_48),
.B1(n_51),
.B2(n_134),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_134),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_134),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_5),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_5),
.A2(n_11),
.B(n_29),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_7),
.A2(n_40),
.B1(n_48),
.B2(n_51),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_8),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_97),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_8),
.A2(n_48),
.B1(n_51),
.B2(n_97),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_97),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_69),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_9),
.A2(n_48),
.B1(n_51),
.B2(n_69),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_11),
.B(n_35),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_11),
.A2(n_35),
.B(n_43),
.C(n_148),
.D(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_11),
.B(n_32),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_11),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_11),
.A2(n_82),
.B(n_165),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_L g195 ( 
.A1(n_11),
.A2(n_30),
.B(n_31),
.C(n_196),
.D(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_11),
.B(n_30),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_180),
.Y(n_243)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_13),
.A2(n_48),
.B1(n_51),
.B2(n_54),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_54),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_16),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_113),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_112),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_98),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_21),
.B(n_98),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_71),
.C(n_79),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_22),
.A2(n_23),
.B1(n_71),
.B2(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_57),
.B2(n_70),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_41),
.B1(n_55),
.B2(n_56),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_26),
.B(n_56),
.C(n_57),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_27),
.A2(n_31),
.B1(n_32),
.B2(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

AOI32xp33_ASAP7_75t_L g206 ( 
.A1(n_29),
.A2(n_35),
.A3(n_196),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_31),
.B(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_31),
.A2(n_32),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g147 ( 
.A1(n_34),
.A2(n_45),
.A3(n_51),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_SL g208 ( 
.A(n_34),
.B(n_38),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_44),
.B(n_46),
.C(n_47),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_44),
.Y(n_46)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_38),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_39),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_41),
.A2(n_56),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_52),
.B(n_53),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_42),
.A2(n_52),
.B1(n_92),
.B2(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_42),
.A2(n_225),
.B(n_226),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_42),
.A2(n_52),
.B1(n_128),
.B2(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_47),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_43),
.A2(n_47),
.B1(n_74),
.B2(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_43),
.B(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_43),
.A2(n_47),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_51),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_44),
.B(n_48),
.Y(n_149)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_83),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_51),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_52),
.B(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_52),
.A2(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_52),
.B(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_52),
.A2(n_161),
.B(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_70),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_67),
.B1(n_68),
.B2(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_58),
.A2(n_132),
.B(n_135),
.Y(n_131)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_59),
.B(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_59),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_59),
.A2(n_60),
.B1(n_133),
.B2(n_266),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_60),
.B(n_96),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_61),
.A2(n_63),
.B(n_180),
.C(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_63),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_67),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_67),
.B(n_180),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_67),
.A2(n_95),
.B(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_73),
.B(n_76),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_78),
.A2(n_107),
.B1(n_109),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_79),
.A2(n_80),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_88),
.B(n_93),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_93),
.B1(n_94),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_81),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_81),
.A2(n_89),
.B1(n_90),
.B2(n_119),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_87),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_82),
.A2(n_86),
.B1(n_87),
.B2(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_82),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_82),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_82),
.B(n_167),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_82),
.A2(n_84),
.B1(n_205),
.B2(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_82),
.A2(n_84),
.B1(n_126),
.B2(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_84),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_84),
.A2(n_172),
.B(n_182),
.Y(n_181)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_85),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_85),
.A2(n_173),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_86),
.B(n_180),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_118),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_111),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_107),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_109),
.B(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_109),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_109),
.A2(n_130),
.B(n_216),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_139),
.B(n_310),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_136),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_115),
.B(n_136),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_298)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_122),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.C(n_131),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_123),
.A2(n_124),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_125),
.B(n_127),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_129),
.B(n_131),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_135),
.Y(n_244)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI321xp33_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_290),
.A3(n_299),
.B1(n_304),
.B2(n_309),
.C(n_312),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_254),
.C(n_286),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_228),
.B(n_253),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_210),
.B(n_227),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_191),
.B(n_209),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_168),
.B(n_190),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_153),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_146),
.B(n_153),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_150),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_163),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_158),
.C(n_163),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_159),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_164),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_177),
.B(n_189),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_170),
.B(n_176),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_183),
.B(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_184),
.B(n_188),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_179),
.B(n_181),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_193),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_202),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_199),
.C(n_202),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_197),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_206),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_212),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_222),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_223),
.C(n_224),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_219),
.C(n_220),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_215),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_221),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_229),
.B(n_230),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_241),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_232),
.B(n_233),
.C(n_241),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.Y(n_233)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_234),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_236),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_240),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_247),
.C(n_250),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_249),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_255),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_273),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_256),
.B(n_273),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_268),
.C(n_272),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_260),
.C(n_267),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_267),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_264),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_272),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_271),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_273)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_282),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_282),
.C(n_285),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_279),
.C(n_280),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_288),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_297),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_297),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.C(n_296),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_295),
.Y(n_303)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_300),
.A2(n_305),
.B(n_308),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_302),
.Y(n_308)
);


endmodule