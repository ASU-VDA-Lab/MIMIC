module fake_jpeg_10677_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_21),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_16),
.B1(n_25),
.B2(n_21),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_44),
.B1(n_37),
.B2(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_16),
.B1(n_25),
.B2(n_28),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_53),
.B1(n_29),
.B2(n_23),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_16),
.B1(n_21),
.B2(n_20),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_40),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_0),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_21),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_19),
.B1(n_28),
.B2(n_29),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_19),
.C(n_22),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_22),
.C(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_65),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_62),
.B(n_87),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_76),
.B1(n_79),
.B2(n_31),
.Y(n_103)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_32),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_71),
.C(n_77),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_78),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_39),
.C(n_30),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_37),
.B1(n_30),
.B2(n_24),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_1),
.B(n_4),
.Y(n_110)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_73),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_81),
.B1(n_88),
.B2(n_52),
.Y(n_91)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_23),
.B1(n_32),
.B2(n_26),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_47),
.C(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_38),
.B1(n_26),
.B2(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_26),
.B1(n_38),
.B2(n_17),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_52),
.B1(n_26),
.B2(n_31),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_17),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_0),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_26),
.C(n_31),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_96),
.B(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_100),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_31),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_104),
.B1(n_82),
.B2(n_68),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_69),
.Y(n_124)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_101),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_31),
.B1(n_14),
.B2(n_11),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_1),
.B(n_3),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_5),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_79),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_84),
.B(n_5),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_85),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_126),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_71),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_113),
.C(n_90),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_117),
.B1(n_99),
.B2(n_14),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_108),
.A2(n_63),
.B1(n_87),
.B2(n_64),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_79),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_122),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_127),
.B(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_76),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_129),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_1),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_92),
.B(n_5),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_135),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_6),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_136),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_6),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_6),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_148),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_135),
.A2(n_100),
.B1(n_103),
.B2(n_102),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_152),
.B1(n_158),
.B2(n_131),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_109),
.B(n_102),
.C(n_92),
.D(n_69),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_144),
.B(n_7),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_101),
.B(n_105),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_113),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_146),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_130),
.A2(n_90),
.B1(n_105),
.B2(n_99),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_120),
.B1(n_137),
.B2(n_125),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_155),
.B(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_7),
.Y(n_156)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_10),
.Y(n_160)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

BUFx4f_ASAP7_75t_SL g161 ( 
.A(n_138),
.Y(n_161)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_166),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_119),
.B1(n_117),
.B2(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_171),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_159),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_116),
.B1(n_133),
.B2(n_129),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_173),
.A2(n_176),
.B(n_177),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_150),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_9),
.B1(n_139),
.B2(n_158),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_145),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_188),
.C(n_192),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_181),
.B(n_147),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_150),
.C(n_142),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_184),
.A2(n_185),
.B(n_189),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_148),
.B(n_149),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_146),
.C(n_160),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_178),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_140),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_165),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_140),
.C(n_149),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_179),
.C(n_175),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_144),
.B(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_181),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_162),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_202),
.B(n_203),
.Y(n_210)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_204),
.A2(n_187),
.B1(n_147),
.B2(n_192),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_211),
.Y(n_215)
);

FAx1_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_190),
.CI(n_186),
.CON(n_206),
.SN(n_206)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_180),
.B(n_196),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_155),
.Y(n_218)
);

NOR2x1_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_175),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_199),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_196),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_218),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_143),
.C(n_156),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_143),
.C(n_208),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_221),
.B(n_222),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_210),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_170),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_206),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_220),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_170),
.B1(n_205),
.B2(n_206),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_217),
.C(n_207),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_228),
.A2(n_229),
.B(n_226),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_216),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_224),
.Y(n_232)
);


endmodule