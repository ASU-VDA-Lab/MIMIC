module fake_jpeg_23897_n_177 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_13),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_1),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_42),
.B1(n_15),
.B2(n_26),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_2),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_20),
.B(n_2),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_3),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_4),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_30),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_61),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_53),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_22),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_57),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_33),
.A2(n_27),
.B1(n_15),
.B2(n_18),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_16),
.B1(n_17),
.B2(n_23),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_85)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_34),
.A2(n_28),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_8),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_42),
.B1(n_30),
.B2(n_25),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_78),
.B1(n_81),
.B2(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_83),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_16),
.B1(n_17),
.B2(n_23),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_23),
.B1(n_45),
.B2(n_21),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_93),
.B(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_47),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_59),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_88),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_94),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_11),
.C(n_12),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_14),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_53),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_86),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_96),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_103),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_110),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_55),
.B1(n_59),
.B2(n_77),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_78),
.B1(n_75),
.B2(n_76),
.Y(n_115)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_88),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_75),
.B(n_90),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_75),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_121),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_100),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_74),
.B1(n_79),
.B2(n_93),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_126),
.B(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_107),
.B1(n_99),
.B2(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_109),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_94),
.B(n_111),
.C(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_97),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_119),
.B(n_126),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_121),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_143),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_122),
.B(n_119),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_97),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_140),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_127),
.C(n_131),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_131),
.B(n_117),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_149),
.B(n_144),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_152),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_116),
.Y(n_152)
);

AOI21x1_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_146),
.B(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_158),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_136),
.B1(n_141),
.B2(n_133),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_160),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_141),
.B1(n_138),
.B2(n_143),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_152),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_166),
.B(n_161),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_170),
.C(n_164),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_162),
.B(n_155),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_128),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_156),
.B(n_129),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

INVxp33_ASAP7_75t_SL g174 ( 
.A(n_172),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_173),
.B(n_170),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_174),
.Y(n_177)
);


endmodule