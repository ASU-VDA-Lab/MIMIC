module fake_jpeg_1941_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_41),
.Y(n_71)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_38),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_50),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_38),
.B1(n_39),
.B2(n_45),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_39),
.B1(n_40),
.B2(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_73),
.Y(n_88)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_44),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_36),
.B1(n_1),
.B2(n_2),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_74),
.B(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_75),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_1),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_64),
.B1(n_58),
.B2(n_54),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_36),
.B1(n_4),
.B2(n_5),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_7),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_73),
.C(n_65),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_100),
.C(n_21),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_6),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_101),
.C(n_4),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_2),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_109),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_87),
.B1(n_82),
.B2(n_7),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_108),
.C(n_112),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_5),
.B(n_6),
.Y(n_109)
);

OAI321xp33_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_22),
.A3(n_33),
.B1(n_32),
.B2(n_31),
.C(n_30),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_111),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_18),
.C(n_28),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_113),
.B(n_8),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_8),
.B(n_9),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_111),
.C(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_118),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_10),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_121),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_107),
.B1(n_97),
.B2(n_12),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_23),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_124),
.B(n_126),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_19),
.C(n_27),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_119),
.B(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_127),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_123),
.B(n_124),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_131),
.A3(n_34),
.B1(n_13),
.B2(n_17),
.C1(n_25),
.C2(n_26),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_10),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_133),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_11),
.Y(n_135)
);


endmodule