module fake_jpeg_7283_n_286 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_19;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_0),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_22),
.C(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_23),
.CON(n_46),
.SN(n_46)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_37),
.B1(n_33),
.B2(n_22),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_61),
.B(n_63),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_27),
.B1(n_28),
.B2(n_23),
.Y(n_61)
);

NAND2x1p5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_31),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_39),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_20),
.C(n_21),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_52),
.B1(n_44),
.B2(n_15),
.Y(n_92)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_71),
.Y(n_93)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_37),
.B1(n_39),
.B2(n_30),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_77),
.Y(n_89)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_37),
.B1(n_18),
.B2(n_22),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_26),
.B1(n_15),
.B2(n_18),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_20),
.B1(n_21),
.B2(n_47),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_38),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_94),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_92),
.B1(n_100),
.B2(n_73),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_71),
.B1(n_73),
.B2(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_32),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_14),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_15),
.B1(n_14),
.B2(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_62),
.B(n_10),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_62),
.B(n_15),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_108),
.B1(n_115),
.B2(n_84),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_95),
.B(n_85),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_110),
.B(n_127),
.Y(n_129)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_84),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_72),
.B1(n_81),
.B2(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_109),
.B(n_124),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_78),
.B(n_66),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_94),
.C(n_103),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_90),
.C(n_93),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_78),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_113),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_119),
.B1(n_110),
.B2(n_122),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_73),
.B1(n_65),
.B2(n_76),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_0),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_13),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_89),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_84),
.B1(n_82),
.B2(n_97),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_12),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_126),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_65),
.B(n_16),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_134),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_129),
.C(n_107),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_0),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_148),
.Y(n_153)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_142),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_91),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

CKINVDCx10_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_82),
.Y(n_139)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_146),
.B1(n_150),
.B2(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_89),
.Y(n_144)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_119),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_76),
.B1(n_64),
.B2(n_75),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_151),
.A2(n_140),
.B1(n_141),
.B2(n_135),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_112),
.B(n_121),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_154),
.B(n_164),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_129),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_156),
.B(n_157),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_167),
.B1(n_145),
.B2(n_137),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_132),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_166),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_122),
.B1(n_89),
.B2(n_64),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_121),
.B1(n_106),
.B2(n_107),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_171),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_152),
.C(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_180),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_142),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_194),
.B(n_153),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_187),
.B1(n_190),
.B2(n_192),
.Y(n_201)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_133),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_191),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_173),
.A2(n_134),
.B1(n_133),
.B2(n_130),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_131),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_195),
.B1(n_191),
.B2(n_184),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_130),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_116),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_196),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_16),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_167),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_154),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_159),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_216),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_209),
.C(n_211),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_213),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_207),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_182),
.C(n_162),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_180),
.A2(n_173),
.B1(n_163),
.B2(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_162),
.C(n_169),
.Y(n_211)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_153),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_153),
.C(n_163),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_36),
.C(n_24),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_185),
.A2(n_174),
.B1(n_116),
.B2(n_77),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_215),
.A2(n_194),
.B1(n_181),
.B2(n_189),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_174),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_186),
.B1(n_194),
.B2(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_16),
.B(n_11),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_203),
.B(n_9),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_77),
.B1(n_64),
.B2(n_11),
.Y(n_224)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_38),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_228),
.C(n_229),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_216),
.C(n_214),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_36),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_24),
.C(n_75),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_206),
.B(n_13),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_233),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_204),
.B(n_24),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_241),
.Y(n_258)
);

A2O1A1O1Ixp25_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_200),
.B(n_206),
.C(n_199),
.D(n_207),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_243),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_246),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_1),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_245),
.Y(n_255)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_1),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_247),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_220),
.C(n_231),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_231),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_237),
.B(n_226),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_252),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_247),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_253),
.B(n_255),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_220),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_256),
.C(n_257),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_227),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_229),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_262),
.B(n_264),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_238),
.C(n_239),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_259),
.A2(n_240),
.B1(n_243),
.B2(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_219),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_249),
.A2(n_219),
.B1(n_2),
.B2(n_3),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_265),
.A2(n_266),
.B1(n_256),
.B2(n_4),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_1),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_2),
.C(n_3),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_248),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_268),
.A2(n_250),
.B(n_257),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_274),
.B(n_3),
.Y(n_277)
);

AOI322xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_272),
.A3(n_265),
.B1(n_261),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_275)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_24),
.A3(n_19),
.B1(n_16),
.B2(n_5),
.C1(n_6),
.C2(n_2),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_277),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_L g278 ( 
.A1(n_273),
.A2(n_24),
.A3(n_19),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_5),
.Y(n_278)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_278),
.A3(n_19),
.B1(n_7),
.B2(n_8),
.C1(n_5),
.C2(n_4),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_279),
.C(n_7),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_4),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_19),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_19),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_19),
.Y(n_286)
);


endmodule