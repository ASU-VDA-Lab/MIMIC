module fake_netlist_1_2272_n_34 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_25;
wire n_26;
wire n_13;
wire n_33;
wire n_16;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_0), .Y(n_8) );
NOR2xp33_ASAP7_75t_R g9 ( .A(n_7), .B(n_0), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
CKINVDCx16_ASAP7_75t_R g11 ( .A(n_4), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx2_ASAP7_75t_SL g15 ( .A(n_10), .Y(n_15) );
BUFx8_ASAP7_75t_SL g16 ( .A(n_8), .Y(n_16) );
O2A1O1Ixp33_ASAP7_75t_L g17 ( .A1(n_12), .A2(n_1), .B(n_2), .C(n_3), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_11), .B(n_1), .Y(n_18) );
O2A1O1Ixp33_ASAP7_75t_L g19 ( .A1(n_12), .A2(n_3), .B(n_4), .C(n_14), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_11), .B(n_10), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_18), .B(n_14), .Y(n_21) );
AND2x6_ASAP7_75t_L g22 ( .A(n_18), .B(n_9), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_15), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_21), .B(n_20), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
INVx1_ASAP7_75t_SL g26 ( .A(n_22), .Y(n_26) );
NAND3xp33_ASAP7_75t_L g27 ( .A(n_24), .B(n_19), .C(n_17), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_24), .B(n_22), .Y(n_28) );
AO22x2_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_26), .B1(n_28), .B2(n_17), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_30), .B(n_26), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
OAI22xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_29), .B1(n_13), .B2(n_25), .Y(n_33) );
AOI22xp5_ASAP7_75t_SL g34 ( .A1(n_33), .A2(n_16), .B1(n_31), .B2(n_25), .Y(n_34) );
endmodule