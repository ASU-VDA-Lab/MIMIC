module fake_jpeg_5258_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_1),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_21),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_20),
.Y(n_49)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_21),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_28),
.B(n_22),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_27),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_60),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_15),
.B1(n_26),
.B2(n_25),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_63),
.B1(n_25),
.B2(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_18),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_27),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_15),
.B1(n_20),
.B2(n_28),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_62),
.B1(n_17),
.B2(n_24),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_15),
.B1(n_21),
.B2(n_28),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_29),
.B1(n_22),
.B2(n_26),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_63),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_32),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_73),
.Y(n_83)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_77),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_37),
.B1(n_35),
.B2(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_41),
.B1(n_40),
.B2(n_37),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_82),
.B1(n_76),
.B2(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_81),
.B(n_54),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_89),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_60),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_100),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_60),
.A3(n_52),
.B1(n_49),
.B2(n_54),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_44),
.B1(n_47),
.B2(n_58),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_52),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_90),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_52),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_95),
.B1(n_97),
.B2(n_99),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_64),
.B1(n_70),
.B2(n_59),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_40),
.B1(n_64),
.B2(n_35),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_59),
.B1(n_45),
.B2(n_55),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_57),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_78),
.B(n_36),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_74),
.B(n_19),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_103),
.B(n_19),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_105),
.Y(n_142)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_79),
.B(n_75),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_115),
.B(n_117),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_108),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_90),
.B1(n_85),
.B2(n_98),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_58),
.B1(n_72),
.B2(n_44),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_83),
.B(n_88),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_122),
.B1(n_123),
.B2(n_95),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_45),
.B1(n_58),
.B2(n_34),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_45),
.B1(n_34),
.B2(n_72),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_125),
.B1(n_140),
.B2(n_27),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_136),
.B1(n_112),
.B2(n_116),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_131),
.B(n_133),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_100),
.C(n_88),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_135),
.C(n_137),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_85),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_114),
.B(n_107),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_89),
.C(n_84),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_102),
.B(n_103),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_99),
.C(n_46),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_36),
.C(n_48),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_2),
.C(n_3),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_48),
.B1(n_31),
.B2(n_30),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_0),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_109),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_14),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_146),
.Y(n_172)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_123),
.B(n_108),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_106),
.B1(n_31),
.B2(n_78),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_151),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_153),
.A2(n_154),
.B1(n_142),
.B2(n_141),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_31),
.B1(n_30),
.B2(n_5),
.Y(n_154)
);

OAI22x1_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_30),
.B1(n_3),
.B2(n_5),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_163),
.B1(n_139),
.B2(n_144),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_157),
.C(n_158),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_14),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_2),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_2),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_130),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_167),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_129),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_153),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_169),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_128),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_171),
.B1(n_178),
.B2(n_124),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_125),
.C(n_135),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_154),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_137),
.B1(n_144),
.B2(n_126),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_161),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_184),
.B(n_185),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_157),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_187),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_139),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_192),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_138),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

XOR2x2_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_163),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_6),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_160),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_6),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_166),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_164),
.C(n_165),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_195),
.C(n_199),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_164),
.C(n_172),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_151),
.B1(n_126),
.B2(n_173),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_200),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_186),
.A2(n_147),
.B1(n_158),
.B2(n_156),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_SL g200 ( 
.A(n_192),
.B(n_3),
.C(n_5),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_6),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_181),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_207),
.B(n_197),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_7),
.Y(n_208)
);

AO22x1_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_203),
.B1(n_11),
.B2(n_14),
.Y(n_216)
);

AOI31xp67_ASAP7_75t_SL g210 ( 
.A1(n_200),
.A2(n_10),
.A3(n_11),
.B(n_13),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_211),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_193),
.C(n_194),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_216),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_208),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_217),
.B(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_214),
.Y(n_222)
);

AOI21x1_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_202),
.B(n_205),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_220),
.B(n_194),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_223),
.B(n_218),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_212),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_10),
.B(n_225),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_10),
.Y(n_228)
);


endmodule