module real_aes_5607_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_894, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_893, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_894;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_893;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_254;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_537;
wire n_320;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_889;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_869;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_0), .A2(n_21), .B1(n_418), .B2(n_419), .Y(n_417) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_1), .Y(n_650) );
AND2x4_ASAP7_75t_L g655 ( .A(n_1), .B(n_228), .Y(n_655) );
AND2x4_ASAP7_75t_L g665 ( .A(n_1), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g413 ( .A(n_2), .Y(n_413) );
AO22x1_ASAP7_75t_L g673 ( .A1(n_3), .A2(n_5), .B1(n_674), .B2(n_675), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_4), .A2(n_86), .B1(n_364), .B2(n_365), .Y(n_637) );
XOR2x2_ASAP7_75t_L g496 ( .A(n_5), .B(n_497), .Y(n_496) );
XNOR2xp5_ASAP7_75t_L g551 ( .A(n_5), .B(n_497), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_6), .A2(n_172), .B1(n_662), .B2(n_680), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_7), .A2(n_124), .B1(n_319), .B2(n_439), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_8), .A2(n_144), .B1(n_361), .B2(n_362), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_9), .B(n_521), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_10), .A2(n_178), .B1(n_244), .B2(n_429), .Y(n_595) );
AOI21xp33_ASAP7_75t_SL g420 ( .A1(n_11), .A2(n_421), .B(n_422), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_12), .A2(n_217), .B1(n_355), .B2(n_357), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_13), .A2(n_189), .B1(n_324), .B2(n_393), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_14), .A2(n_866), .B(n_867), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_15), .A2(n_203), .B1(n_352), .B2(n_358), .Y(n_606) );
INVx1_ASAP7_75t_L g506 ( .A(n_16), .Y(n_506) );
INVx1_ASAP7_75t_L g345 ( .A(n_17), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_17), .A2(n_103), .B1(n_670), .B2(n_707), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_18), .A2(n_29), .B1(n_547), .B2(n_548), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_19), .A2(n_102), .B1(n_305), .B2(n_403), .Y(n_573) );
AO22x1_ASAP7_75t_L g616 ( .A1(n_20), .A2(n_131), .B1(n_368), .B2(n_369), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_22), .A2(n_207), .B1(n_303), .B2(n_597), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_23), .A2(n_167), .B1(n_312), .B2(n_319), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_24), .A2(n_180), .B1(n_336), .B2(n_338), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_25), .A2(n_95), .B1(n_479), .B2(n_480), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_26), .A2(n_134), .B1(n_324), .B2(n_542), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_27), .A2(n_56), .B1(n_357), .B2(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g584 ( .A(n_28), .Y(n_584) );
INVx1_ASAP7_75t_L g517 ( .A(n_30), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_31), .A2(n_374), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g264 ( .A(n_32), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_32), .B(n_184), .Y(n_281) );
INVxp67_ASAP7_75t_L g300 ( .A(n_32), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_33), .A2(n_187), .B1(n_396), .B2(n_397), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_34), .A2(n_106), .B1(n_319), .B2(n_547), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_35), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_36), .A2(n_78), .B1(n_489), .B2(n_491), .Y(n_488) );
AOI21xp33_ASAP7_75t_SL g529 ( .A1(n_37), .A2(n_508), .B(n_530), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_38), .A2(n_128), .B1(n_312), .B2(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_39), .B(n_425), .Y(n_424) );
AO22x1_ASAP7_75t_L g614 ( .A1(n_40), .A2(n_125), .B1(n_364), .B2(n_365), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_41), .A2(n_62), .B1(n_350), .B2(n_374), .C(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_42), .B(n_249), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_43), .A2(n_224), .B1(n_290), .B2(n_292), .Y(n_289) );
OAI21x1_ASAP7_75t_L g621 ( .A1(n_44), .A2(n_622), .B(n_638), .Y(n_621) );
NAND4xp25_ASAP7_75t_L g638 ( .A(n_44), .B(n_623), .C(n_627), .D(n_635), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g243 ( .A1(n_45), .A2(n_65), .B1(n_244), .B2(n_267), .C(n_273), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_46), .A2(n_213), .B1(n_303), .B2(n_305), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_47), .A2(n_164), .B1(n_393), .B2(n_455), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_48), .A2(n_182), .B1(n_401), .B2(n_429), .Y(n_428) );
NAND2xp33_ASAP7_75t_L g348 ( .A(n_49), .B(n_349), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_50), .A2(n_148), .B1(n_669), .B2(n_675), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_51), .A2(n_140), .B1(n_501), .B2(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_52), .A2(n_92), .B1(n_303), .B2(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_53), .B(n_350), .Y(n_605) );
INVx2_ASAP7_75t_L g648 ( .A(n_54), .Y(n_648) );
XNOR2x1_ASAP7_75t_L g556 ( .A(n_55), .B(n_557), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_57), .A2(n_155), .B1(n_435), .B2(n_437), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_58), .A2(n_188), .B1(n_290), .B2(n_292), .Y(n_535) );
AND2x4_ASAP7_75t_L g656 ( .A(n_59), .B(n_648), .Y(n_656) );
INVx1_ASAP7_75t_L g664 ( .A(n_59), .Y(n_664) );
INVx1_ASAP7_75t_SL g705 ( .A(n_59), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_60), .A2(n_61), .B1(n_324), .B2(n_326), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_63), .A2(n_166), .B1(n_654), .B2(n_674), .Y(n_742) );
XNOR2x1_ASAP7_75t_L g862 ( .A(n_63), .B(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_63), .A2(n_883), .B1(n_885), .B2(n_889), .Y(n_882) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_64), .A2(n_581), .B(n_583), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_66), .A2(n_137), .B1(n_432), .B2(n_439), .Y(n_636) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_67), .Y(n_249) );
INVx1_ASAP7_75t_L g376 ( .A(n_68), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_69), .A2(n_165), .B1(n_355), .B2(n_357), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_70), .A2(n_173), .B1(n_352), .B2(n_353), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_71), .A2(n_159), .B1(n_352), .B2(n_358), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_72), .A2(n_221), .B1(n_361), .B2(n_626), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_73), .A2(n_205), .B1(n_390), .B2(n_391), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_74), .A2(n_139), .B1(n_662), .B2(n_667), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_75), .A2(n_119), .B1(n_332), .B2(n_464), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_76), .A2(n_108), .B1(n_575), .B2(n_576), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_77), .A2(n_152), .B1(n_674), .B2(n_675), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_79), .A2(n_171), .B1(n_669), .B2(n_675), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_80), .A2(n_191), .B1(n_432), .B2(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g253 ( .A(n_81), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_81), .B(n_183), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_82), .A2(n_142), .B1(n_433), .B2(n_550), .Y(n_873) );
INVx1_ASAP7_75t_L g630 ( .A(n_83), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_84), .A2(n_87), .B1(n_336), .B2(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_85), .A2(n_138), .B1(n_439), .B2(n_440), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_88), .A2(n_146), .B1(n_662), .B2(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_89), .A2(n_96), .B1(n_662), .B2(n_680), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_90), .A2(n_170), .B1(n_324), .B2(n_326), .Y(n_502) );
INVx1_ASAP7_75t_L g610 ( .A(n_91), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_93), .A2(n_199), .B1(n_390), .B2(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_94), .B(n_572), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_97), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_98), .A2(n_174), .B1(n_336), .B2(n_387), .Y(n_503) );
INVx1_ASAP7_75t_L g423 ( .A(n_99), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_100), .A2(n_186), .B1(n_695), .B2(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g408 ( .A(n_101), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_104), .A2(n_112), .B1(n_471), .B2(n_472), .Y(n_470) );
XNOR2x1_ASAP7_75t_L g382 ( .A(n_105), .B(n_383), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_107), .A2(n_160), .B1(n_324), .B2(n_393), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_109), .A2(n_220), .B1(n_662), .B2(n_680), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_110), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_111), .A2(n_227), .B1(n_336), .B2(n_564), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_113), .A2(n_122), .B1(n_541), .B2(n_542), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_114), .A2(n_163), .B1(n_326), .B2(n_541), .Y(n_588) );
AO22x1_ASAP7_75t_L g615 ( .A1(n_115), .A2(n_226), .B1(n_371), .B2(n_372), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_116), .A2(n_129), .B1(n_455), .B2(n_457), .Y(n_454) );
INVx1_ASAP7_75t_L g515 ( .A(n_117), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_118), .A2(n_181), .B1(n_364), .B2(n_365), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_120), .A2(n_196), .B1(n_312), .B2(n_319), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_121), .A2(n_200), .B1(n_329), .B2(n_332), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_123), .A2(n_204), .B1(n_336), .B2(n_564), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_126), .A2(n_229), .B1(n_485), .B2(n_487), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_127), .A2(n_130), .B1(n_537), .B2(n_538), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_132), .A2(n_218), .B1(n_680), .B2(n_704), .Y(n_703) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_133), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_135), .A2(n_147), .B1(n_361), .B2(n_362), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_136), .B(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_141), .A2(n_211), .B1(n_550), .B2(n_561), .Y(n_560) );
XNOR2x2_ASAP7_75t_L g602 ( .A(n_143), .B(n_603), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_145), .A2(n_192), .B1(n_669), .B2(n_670), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_149), .A2(n_209), .B1(n_336), .B2(n_387), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_150), .A2(n_190), .B1(n_403), .B2(n_405), .C(n_407), .Y(n_402) );
AO221x2_ASAP7_75t_L g672 ( .A1(n_151), .A2(n_198), .B1(n_662), .B2(n_667), .C(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_153), .A2(n_206), .B1(n_479), .B2(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g569 ( .A(n_154), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_156), .B(n_521), .Y(n_869) );
OA22x2_ASAP7_75t_L g247 ( .A1(n_157), .A2(n_184), .B1(n_248), .B2(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g288 ( .A(n_157), .Y(n_288) );
INVx1_ASAP7_75t_L g513 ( .A(n_158), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_161), .A2(n_214), .B1(n_387), .B2(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_162), .A2(n_233), .B1(n_312), .B2(n_464), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_168), .A2(n_225), .B1(n_324), .B2(n_326), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_169), .A2(n_223), .B1(n_654), .B2(n_669), .Y(n_697) );
INVx1_ASAP7_75t_L g531 ( .A(n_175), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_176), .A2(n_201), .B1(n_501), .B2(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_177), .A2(n_216), .B1(n_429), .B2(n_575), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_179), .A2(n_193), .B1(n_368), .B2(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g266 ( .A(n_183), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_183), .B(n_285), .Y(n_284) );
OAI21xp33_ASAP7_75t_L g309 ( .A1(n_184), .A2(n_195), .B(n_301), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_185), .Y(n_240) );
INVx1_ASAP7_75t_L g524 ( .A(n_192), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_194), .A2(n_231), .B1(n_371), .B2(n_372), .Y(n_370) );
INVx1_ASAP7_75t_L g255 ( .A(n_195), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_195), .B(n_222), .Y(n_282) );
CKINVDCx16_ASAP7_75t_R g868 ( .A(n_197), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_202), .A2(n_210), .B1(n_399), .B2(n_401), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_208), .A2(n_567), .B(n_568), .Y(n_566) );
OAI22xp33_ASAP7_75t_R g885 ( .A1(n_212), .A2(n_886), .B1(n_887), .B2(n_888), .Y(n_885) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_212), .Y(n_886) );
AOI21xp33_ASAP7_75t_SL g373 ( .A1(n_215), .A2(n_374), .B(n_375), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_219), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_222), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g666 ( .A(n_228), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_230), .Y(n_274) );
INVx1_ASAP7_75t_L g510 ( .A(n_232), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_448), .B(n_642), .C(n_651), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_235), .A2(n_448), .B(n_643), .Y(n_642) );
XOR2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_379), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_341), .B1(n_377), .B2(n_378), .Y(n_236) );
INVx2_ASAP7_75t_L g377 ( .A(n_237), .Y(n_377) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
XNOR2x1_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_310), .Y(n_241) );
NAND3xp33_ASAP7_75t_L g242 ( .A(n_243), .B(n_289), .C(n_302), .Y(n_242) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
BUFx3_ASAP7_75t_L g396 ( .A(n_245), .Y(n_396) );
BUFx3_ASAP7_75t_L g418 ( .A(n_245), .Y(n_418) );
INVx1_ASAP7_75t_L g509 ( .A(n_245), .Y(n_509) );
AND2x4_ASAP7_75t_L g245 ( .A(n_246), .B(n_256), .Y(n_245) );
AND2x4_ASAP7_75t_L g304 ( .A(n_246), .B(n_271), .Y(n_304) );
AND2x4_ASAP7_75t_L g357 ( .A(n_246), .B(n_256), .Y(n_357) );
AND2x2_ASAP7_75t_L g374 ( .A(n_246), .B(n_271), .Y(n_374) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_250), .Y(n_246) );
AND2x2_ASAP7_75t_L g270 ( .A(n_247), .B(n_251), .Y(n_270) );
AND2x2_ASAP7_75t_L g298 ( .A(n_247), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g315 ( .A(n_247), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_248), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp33_ASAP7_75t_L g252 ( .A(n_249), .B(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g259 ( .A(n_249), .Y(n_259) );
NAND2xp33_ASAP7_75t_L g265 ( .A(n_249), .B(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_249), .Y(n_279) );
INVx1_ASAP7_75t_L g301 ( .A(n_249), .Y(n_301) );
AND2x4_ASAP7_75t_L g314 ( .A(n_250), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_253), .B(n_288), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g299 ( .A1(n_255), .A2(n_300), .B(n_301), .Y(n_299) );
AND2x2_ASAP7_75t_L g291 ( .A(n_256), .B(n_270), .Y(n_291) );
AND2x4_ASAP7_75t_L g325 ( .A(n_256), .B(n_314), .Y(n_325) );
AND2x4_ASAP7_75t_L g352 ( .A(n_256), .B(n_270), .Y(n_352) );
AND2x4_ASAP7_75t_L g368 ( .A(n_256), .B(n_314), .Y(n_368) );
AND2x4_ASAP7_75t_L g256 ( .A(n_257), .B(n_261), .Y(n_256) );
INVx2_ASAP7_75t_L g272 ( .A(n_257), .Y(n_272) );
AND2x2_ASAP7_75t_L g295 ( .A(n_257), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g316 ( .A(n_257), .B(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g322 ( .A(n_257), .B(n_318), .Y(n_322) );
AND2x4_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_259), .B(n_264), .Y(n_263) );
INVxp67_ASAP7_75t_L g285 ( .A(n_259), .Y(n_285) );
NAND3xp33_ASAP7_75t_L g283 ( .A(n_260), .B(n_284), .C(n_286), .Y(n_283) );
AND2x4_ASAP7_75t_L g271 ( .A(n_261), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g318 ( .A(n_262), .Y(n_318) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
INVx2_ASAP7_75t_L g582 ( .A(n_267), .Y(n_582) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g519 ( .A(n_268), .Y(n_519) );
INVx2_ASAP7_75t_L g567 ( .A(n_268), .Y(n_567) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g427 ( .A(n_269), .Y(n_427) );
BUFx3_ASAP7_75t_L g477 ( .A(n_269), .Y(n_477) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
AND2x4_ASAP7_75t_L g330 ( .A(n_270), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g337 ( .A(n_270), .B(n_316), .Y(n_337) );
AND2x2_ASAP7_75t_L g350 ( .A(n_270), .B(n_271), .Y(n_350) );
AND2x4_ASAP7_75t_L g361 ( .A(n_270), .B(n_321), .Y(n_361) );
AND2x4_ASAP7_75t_L g364 ( .A(n_270), .B(n_316), .Y(n_364) );
AND2x2_ASAP7_75t_L g436 ( .A(n_270), .B(n_316), .Y(n_436) );
AND2x4_ASAP7_75t_L g307 ( .A(n_271), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g327 ( .A(n_271), .B(n_314), .Y(n_327) );
AND2x4_ASAP7_75t_L g355 ( .A(n_271), .B(n_308), .Y(n_355) );
AND2x4_ASAP7_75t_L g369 ( .A(n_271), .B(n_314), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_275), .B(n_376), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_275), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g572 ( .A(n_275), .Y(n_572) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_SL g410 ( .A(n_276), .Y(n_410) );
INVx2_ASAP7_75t_L g533 ( .A(n_276), .Y(n_533) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx3_ASAP7_75t_L g482 ( .A(n_277), .Y(n_482) );
AO21x2_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_280), .B(n_283), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_279), .B(n_297), .Y(n_296) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_280), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_285), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g308 ( .A(n_286), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g511 ( .A(n_290), .Y(n_511) );
BUFx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g400 ( .A(n_291), .Y(n_400) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_291), .Y(n_429) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx4_ASAP7_75t_L g397 ( .A(n_293), .Y(n_397) );
INVx5_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_L g419 ( .A(n_294), .Y(n_419) );
BUFx4f_ASAP7_75t_L g479 ( .A(n_294), .Y(n_479) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
AND2x4_ASAP7_75t_L g358 ( .A(n_295), .B(n_298), .Y(n_358) );
INVx2_ASAP7_75t_L g514 ( .A(n_303), .Y(n_514) );
BUFx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g404 ( .A(n_304), .Y(n_404) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_304), .Y(n_421) );
INVx2_ASAP7_75t_L g490 ( .A(n_304), .Y(n_490) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g491 ( .A(n_306), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_306), .A2(n_513), .B1(n_514), .B2(n_515), .Y(n_512) );
INVx3_ASAP7_75t_L g597 ( .A(n_306), .Y(n_597) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_307), .Y(n_401) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_307), .Y(n_538) );
AND2x4_ASAP7_75t_L g334 ( .A(n_308), .B(n_321), .Y(n_334) );
AND2x4_ASAP7_75t_L g340 ( .A(n_308), .B(n_316), .Y(n_340) );
AND2x4_ASAP7_75t_L g362 ( .A(n_308), .B(n_321), .Y(n_362) );
AND2x4_ASAP7_75t_L g365 ( .A(n_308), .B(n_316), .Y(n_365) );
NAND4xp25_ASAP7_75t_SL g310 ( .A(n_311), .B(n_323), .C(n_328), .D(n_335), .Y(n_310) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx12f_ASAP7_75t_L g439 ( .A(n_313), .Y(n_439) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_313), .Y(n_547) );
AND2x4_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
AND2x4_ASAP7_75t_L g320 ( .A(n_314), .B(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g371 ( .A(n_314), .B(n_316), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_314), .B(n_331), .Y(n_372) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_320), .Y(n_432) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_320), .Y(n_464) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_320), .Y(n_548) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g331 ( .A(n_322), .Y(n_331) );
BUFx12f_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx3_ASAP7_75t_L g456 ( .A(n_325), .Y(n_456) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_325), .Y(n_541) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx3_ASAP7_75t_L g393 ( .A(n_327), .Y(n_393) );
BUFx5_ASAP7_75t_L g542 ( .A(n_327), .Y(n_542) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_330), .Y(n_390) );
BUFx12f_ASAP7_75t_L g437 ( .A(n_330), .Y(n_437) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_330), .Y(n_550) );
BUFx3_ASAP7_75t_L g593 ( .A(n_330), .Y(n_593) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g391 ( .A(n_333), .Y(n_391) );
INVx5_ASAP7_75t_L g433 ( .A(n_333), .Y(n_433) );
INVx3_ASAP7_75t_L g626 ( .A(n_333), .Y(n_626) );
INVx6_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx12f_ASAP7_75t_L g501 ( .A(n_334), .Y(n_501) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx8_ASAP7_75t_L g459 ( .A(n_337), .Y(n_459) );
INVx4_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx4_ASAP7_75t_L g387 ( .A(n_339), .Y(n_387) );
INVx1_ASAP7_75t_L g440 ( .A(n_339), .Y(n_440) );
INVx2_ASAP7_75t_L g544 ( .A(n_339), .Y(n_544) );
INVx4_ASAP7_75t_L g564 ( .A(n_339), .Y(n_564) );
INVx8_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g378 ( .A(n_341), .Y(n_378) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx3_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
XNOR2x1_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
NOR2x1_ASAP7_75t_L g346 ( .A(n_347), .B(n_359), .Y(n_346) );
NAND3xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .C(n_356), .Y(n_347) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g406 ( .A(n_350), .Y(n_406) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx4_ASAP7_75t_L g570 ( .A(n_358), .Y(n_570) );
NAND4xp25_ASAP7_75t_SL g359 ( .A(n_360), .B(n_363), .C(n_366), .D(n_373), .Y(n_359) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_370), .Y(n_366) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
XNOR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_411), .Y(n_381) );
NAND4xp75_ASAP7_75t_L g383 ( .A(n_384), .B(n_388), .C(n_394), .D(n_402), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
BUFx3_ASAP7_75t_L g471 ( .A(n_390), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_391), .Y(n_472) );
BUFx2_ASAP7_75t_L g457 ( .A(n_393), .Y(n_457) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_398), .Y(n_394) );
INVx2_ASAP7_75t_L g486 ( .A(n_396), .Y(n_486) );
INVx2_ASAP7_75t_L g585 ( .A(n_397), .Y(n_585) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g576 ( .A(n_400), .Y(n_576) );
INVx2_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_SL g537 ( .A(n_404), .Y(n_537) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
OAI21x1_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B(n_442), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_412), .B(n_428), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_413), .Y(n_412) );
NOR2xp67_ASAP7_75t_L g414 ( .A(n_415), .B(n_430), .Y(n_414) );
NAND3xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_424), .C(n_428), .Y(n_415) );
INVx1_ASAP7_75t_L g446 ( .A(n_416), .Y(n_446) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .Y(n_416) );
INVxp67_ASAP7_75t_L g444 ( .A(n_424), .Y(n_444) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g528 ( .A(n_426), .Y(n_528) );
INVx2_ASAP7_75t_L g866 ( .A(n_426), .Y(n_866) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx3_ASAP7_75t_L g487 ( .A(n_429), .Y(n_487) );
INVx1_ASAP7_75t_L g447 ( .A(n_430), .Y(n_447) );
NAND4xp25_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .C(n_438), .D(n_441), .Y(n_430) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx4f_ASAP7_75t_L g561 ( .A(n_436), .Y(n_561) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_439), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_447), .Y(n_442) );
NOR3xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .C(n_446), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B1(n_552), .B2(n_641), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
XNOR2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_495), .Y(n_450) );
AO211x2_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_468), .B(n_493), .C(n_494), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_460), .Y(n_452) );
AO22x2_ASAP7_75t_L g494 ( .A1(n_453), .A2(n_469), .B1(n_492), .B2(n_894), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_454), .B(n_458), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AO22x1_ASAP7_75t_L g493 ( .A1(n_460), .A2(n_483), .B1(n_492), .B2(n_893), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B1(n_465), .B2(n_466), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_483), .C(n_492), .Y(n_468) );
NAND2x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_478), .Y(n_473) );
INVx1_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
BUFx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx4_ASAP7_75t_L g521 ( .A(n_481), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_481), .B(n_610), .Y(n_609) );
INVx4_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g631 ( .A(n_482), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_488), .Y(n_483) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AOI22x1_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_522), .B1(n_523), .B2(n_551), .Y(n_495) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .Y(n_497) );
AND4x1_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .C(n_502), .D(n_503), .Y(n_498) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_512), .C(n_516), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B1(n_510), .B2(n_511), .Y(n_505) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g575 ( .A(n_509), .Y(n_575) );
OAI21xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_520), .Y(n_516) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
XNOR2x1_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
NOR4xp75_ASAP7_75t_L g525 ( .A(n_526), .B(n_534), .C(n_539), .D(n_545), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_540), .B(n_543), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_546), .B(n_549), .Y(n_545) );
INVx1_ASAP7_75t_L g641 ( .A(n_552), .Y(n_641) );
XNOR2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_600), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B1(n_577), .B2(n_599), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_565), .Y(n_557) );
NAND4xp25_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .C(n_562), .D(n_563), .Y(n_558) );
NAND3xp33_ASAP7_75t_SL g565 ( .A(n_566), .B(n_573), .C(n_574), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B(n_571), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g867 ( .A1(n_570), .A2(n_868), .B(n_869), .Y(n_867) );
INVx2_ASAP7_75t_SL g599 ( .A(n_577), .Y(n_599) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
XNOR2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_598), .Y(n_578) );
NAND4xp75_ASAP7_75t_L g579 ( .A(n_580), .B(n_587), .C(n_590), .D(n_594), .Y(n_579) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B(n_586), .Y(n_583) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AO22x2_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_617), .B1(n_639), .B2(n_640), .Y(n_600) );
INVx2_ASAP7_75t_L g639 ( .A(n_601), .Y(n_639) );
BUFx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_611), .Y(n_603) );
AND4x1_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .C(n_607), .D(n_608), .Y(n_604) );
NOR4xp25_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .C(n_615), .D(n_616), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g640 ( .A(n_619), .Y(n_640) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND3x1_ASAP7_75t_L g622 ( .A(n_623), .B(n_627), .C(n_635), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_632), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
BUFx10_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_649), .C(n_650), .Y(n_645) );
AND2x2_ASAP7_75t_L g879 ( .A(n_646), .B(n_880), .Y(n_879) );
AND2x2_ASAP7_75t_L g884 ( .A(n_646), .B(n_881), .Y(n_884) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OA21x2_ASAP7_75t_L g890 ( .A1(n_647), .A2(n_705), .B(n_891), .Y(n_890) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g663 ( .A(n_648), .B(n_664), .Y(n_663) );
AND3x4_ASAP7_75t_L g704 ( .A(n_648), .B(n_665), .C(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g880 ( .A(n_649), .B(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_650), .Y(n_881) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_657), .B1(n_860), .B2(n_877), .C(n_882), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_653), .Y(n_652) );
BUFx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x4_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
AND2x2_ASAP7_75t_L g669 ( .A(n_655), .B(n_663), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_655), .B(n_656), .Y(n_670) );
AND2x4_ASAP7_75t_L g674 ( .A(n_655), .B(n_663), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_655), .B(n_656), .Y(n_675) );
AND2x2_ASAP7_75t_L g707 ( .A(n_655), .B(n_663), .Y(n_707) );
CKINVDCx5p33_ASAP7_75t_R g891 ( .A(n_655), .Y(n_891) );
AND2x4_ASAP7_75t_L g667 ( .A(n_656), .B(n_665), .Y(n_667) );
AND2x4_ASAP7_75t_L g680 ( .A(n_656), .B(n_665), .Y(n_680) );
AOI221x1_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_737), .B1(n_738), .B2(n_743), .C(n_782), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_676), .B(n_689), .C(n_732), .Y(n_658) );
INVx1_ASAP7_75t_L g754 ( .A(n_659), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_671), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_660), .B(n_701), .Y(n_721) );
CKINVDCx6p67_ASAP7_75t_R g724 ( .A(n_660), .Y(n_724) );
AND2x2_ASAP7_75t_L g731 ( .A(n_660), .B(n_727), .Y(n_731) );
AND2x2_ASAP7_75t_L g746 ( .A(n_660), .B(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_L g776 ( .A(n_660), .B(n_767), .Y(n_776) );
AND2x2_ASAP7_75t_L g804 ( .A(n_660), .B(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g810 ( .A(n_660), .B(n_725), .Y(n_810) );
AND2x2_ASAP7_75t_L g828 ( .A(n_660), .B(n_734), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_660), .B(n_672), .Y(n_842) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_668), .Y(n_660) );
INVx3_ASAP7_75t_L g741 ( .A(n_662), .Y(n_741) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
AND2x2_ASAP7_75t_L g767 ( .A(n_671), .B(n_702), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_671), .B(n_724), .Y(n_837) );
NOR3xp33_ASAP7_75t_L g858 ( .A(n_671), .B(n_677), .C(n_738), .Y(n_858) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g725 ( .A(n_672), .B(n_702), .Y(n_725) );
AND2x2_ASAP7_75t_L g727 ( .A(n_672), .B(n_701), .Y(n_727) );
OR2x2_ASAP7_75t_L g735 ( .A(n_672), .B(n_702), .Y(n_735) );
AND2x2_ASAP7_75t_L g774 ( .A(n_672), .B(n_724), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g787 ( .A1(n_672), .A2(n_676), .B1(n_788), .B2(n_790), .C(n_791), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_681), .Y(n_676) );
INVx2_ASAP7_75t_L g709 ( .A(n_677), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_677), .B(n_686), .Y(n_712) );
INVx3_ASAP7_75t_L g726 ( .A(n_677), .Y(n_726) );
INVx2_ASAP7_75t_L g750 ( .A(n_677), .Y(n_750) );
AND2x2_ASAP7_75t_L g761 ( .A(n_677), .B(n_724), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_677), .B(n_768), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_677), .B(n_692), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_677), .B(n_842), .Y(n_841) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx2_ASAP7_75t_SL g696 ( .A(n_680), .Y(n_696) );
A2O1A1Ixp33_ASAP7_75t_L g732 ( .A1(n_681), .A2(n_731), .B(n_733), .C(n_736), .Y(n_732) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_686), .Y(n_681) );
INVx2_ASAP7_75t_L g698 ( .A(n_682), .Y(n_698) );
AND2x2_ASAP7_75t_L g719 ( .A(n_682), .B(n_692), .Y(n_719) );
OR2x2_ASAP7_75t_L g764 ( .A(n_682), .B(n_718), .Y(n_764) );
INVxp67_ASAP7_75t_L g794 ( .A(n_682), .Y(n_794) );
OR2x2_ASAP7_75t_L g796 ( .A(n_682), .B(n_686), .Y(n_796) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g751 ( .A(n_683), .B(n_686), .Y(n_751) );
AND2x2_ASAP7_75t_L g813 ( .A(n_683), .B(n_693), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_686), .B(n_709), .Y(n_708) );
INVx4_ASAP7_75t_L g718 ( .A(n_686), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_686), .B(n_709), .Y(n_770) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_699), .B(n_710), .C(n_728), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g775 ( .A1(n_690), .A2(n_776), .B(n_777), .C(n_778), .Y(n_775) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_691), .B(n_786), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_698), .Y(n_691) );
INVx2_ASAP7_75t_L g753 ( .A(n_692), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_692), .B(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g771 ( .A(n_692), .B(n_730), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_692), .B(n_751), .Y(n_781) );
OR2x2_ASAP7_75t_L g819 ( .A(n_692), .B(n_794), .Y(n_819) );
INVx4_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g736 ( .A(n_693), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_693), .B(n_757), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_693), .B(n_764), .Y(n_763) );
NOR3xp33_ASAP7_75t_SL g769 ( .A(n_693), .B(n_766), .C(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g829 ( .A(n_693), .B(n_830), .Y(n_829) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx3_ASAP7_75t_SL g744 ( .A(n_698), .Y(n_744) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_708), .Y(n_700) );
AOI211xp5_ASAP7_75t_L g791 ( .A1(n_701), .A2(n_712), .B(n_792), .C(n_798), .Y(n_791) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_706), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_709), .B(n_720), .Y(n_777) );
AND2x2_ASAP7_75t_L g844 ( .A(n_709), .B(n_774), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_709), .B(n_716), .Y(n_857) );
A2O1A1Ixp33_ASAP7_75t_SL g710 ( .A1(n_711), .A2(n_713), .B(n_720), .C(n_722), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_711), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI32xp33_ASAP7_75t_L g722 ( .A1(n_712), .A2(n_719), .A3(n_723), .B1(n_726), .B2(n_727), .Y(n_722) );
INVx1_ASAP7_75t_L g824 ( .A(n_713), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_719), .Y(n_713) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_714), .Y(n_785) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g820 ( .A(n_715), .Y(n_820) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_716), .Y(n_812) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g757 ( .A(n_717), .Y(n_757) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g730 ( .A(n_718), .Y(n_730) );
INVx1_ASAP7_75t_L g808 ( .A(n_719), .Y(n_808) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_721), .B(n_726), .Y(n_795) );
INVx1_ASAP7_75t_L g779 ( .A(n_723), .Y(n_779) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
AND2x2_ASAP7_75t_L g733 ( .A(n_724), .B(n_734), .Y(n_733) );
AOI322xp5_ASAP7_75t_L g762 ( .A1(n_724), .A2(n_744), .A3(n_763), .B1(n_765), .B2(n_769), .C1(n_771), .C2(n_772), .Y(n_762) );
AND2x2_ASAP7_75t_L g789 ( .A(n_724), .B(n_727), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_724), .B(n_767), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_724), .B(n_747), .Y(n_826) );
AND2x2_ASAP7_75t_L g747 ( .A(n_725), .B(n_726), .Y(n_747) );
INVx1_ASAP7_75t_L g797 ( .A(n_725), .Y(n_797) );
INVx3_ASAP7_75t_L g805 ( .A(n_726), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_726), .B(n_789), .Y(n_832) );
AND2x2_ASAP7_75t_L g760 ( .A(n_727), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g768 ( .A(n_727), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_727), .B(n_804), .Y(n_818) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g758 ( .A(n_731), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_731), .B(n_807), .Y(n_806) );
AND2x2_ASAP7_75t_L g803 ( .A(n_734), .B(n_804), .Y(n_803) );
AND2x2_ASAP7_75t_L g834 ( .A(n_734), .B(n_761), .Y(n_834) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_737), .B(n_753), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g737 ( .A(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_742), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI211xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B(n_748), .C(n_775), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_744), .A2(n_790), .B1(n_840), .B2(n_843), .Y(n_839) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
O2A1O1Ixp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B(n_754), .C(n_755), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_750), .B(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_750), .B(n_776), .Y(n_786) );
AND2x2_ASAP7_75t_L g847 ( .A(n_750), .B(n_830), .Y(n_847) );
OAI21xp33_ASAP7_75t_L g825 ( .A1(n_751), .A2(n_826), .B(n_827), .Y(n_825) );
INVx1_ASAP7_75t_L g859 ( .A(n_751), .Y(n_859) );
AOI221xp5_ASAP7_75t_SL g835 ( .A1(n_753), .A2(n_830), .B1(n_836), .B2(n_839), .C(n_845), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_754), .B(n_847), .Y(n_846) );
OAI211xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_758), .B(n_759), .C(n_762), .Y(n_755) );
INVx2_ASAP7_75t_L g790 ( .A(n_757), .Y(n_790) );
A2O1A1Ixp33_ASAP7_75t_SL g836 ( .A1(n_758), .A2(n_833), .B(n_837), .C(n_838), .Y(n_836) );
INVx1_ASAP7_75t_L g830 ( .A(n_764), .Y(n_830) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_768), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g807 ( .A(n_770), .Y(n_807) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g852 ( .A(n_776), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND5xp2_ASAP7_75t_L g782 ( .A(n_783), .B(n_821), .C(n_835), .D(n_848), .E(n_850), .Y(n_782) );
O2A1O1Ixp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_787), .B(n_799), .C(n_801), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_788), .B(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
AOI222xp33_ASAP7_75t_L g850 ( .A1(n_789), .A2(n_851), .B1(n_853), .B2(n_855), .C1(n_858), .C2(n_859), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_790), .B(n_803), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_795), .B1(n_796), .B2(n_797), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g816 ( .A(n_796), .Y(n_816) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_806), .B(n_808), .C(n_809), .Y(n_801) );
NOR2x1_ASAP7_75t_L g814 ( .A(n_805), .B(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g822 ( .A(n_805), .B(n_823), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_805), .B(n_816), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_808), .B(n_856), .Y(n_855) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B1(n_814), .B2(n_816), .C(n_817), .Y(n_809) );
AND2x2_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g823 ( .A(n_815), .Y(n_823) );
NOR3xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .C(n_820), .Y(n_817) );
AOI21xp33_ASAP7_75t_L g831 ( .A1(n_819), .A2(n_832), .B(n_833), .Y(n_831) );
AOI211xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_824), .B(n_825), .C(n_831), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVxp33_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_863), .Y(n_887) );
OR2x2_ASAP7_75t_L g863 ( .A(n_864), .B(n_872), .Y(n_863) );
NAND3xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_870), .C(n_871), .Y(n_864) );
NAND4xp25_ASAP7_75t_SL g872 ( .A(n_873), .B(n_874), .C(n_875), .D(n_876), .Y(n_872) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
BUFx3_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g888 ( .A(n_887), .Y(n_888) );
BUFx2_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
endmodule