module fake_jpeg_2481_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

INVx4_ASAP7_75t_SL g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g12 ( 
.A(n_4),
.B(n_0),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_1),
.C(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_15),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_10),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_32),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_16),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_27)
);

AO21x2_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_13),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_17),
.B(n_24),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

OAI21x1_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_13),
.B(n_28),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_39),
.B(n_29),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_26),
.B(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_43),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_35),
.B2(n_44),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_37),
.C(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_45),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_48),
.B(n_47),
.C(n_35),
.Y(n_50)
);


endmodule