module fake_jpeg_19964_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_8),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_30),
.B1(n_23),
.B2(n_27),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_45),
.B1(n_47),
.B2(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_49),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_30),
.B1(n_31),
.B2(n_19),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_30),
.B1(n_35),
.B2(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_39),
.B1(n_25),
.B2(n_22),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_16),
.B(n_26),
.Y(n_51)
);

FAx1_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_37),
.CI(n_38),
.CON(n_72),
.SN(n_72)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_16),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_56),
.B(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_59),
.B(n_67),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_47),
.Y(n_65)
);

INVxp67_ASAP7_75t_SL g92 ( 
.A(n_65),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_18),
.B1(n_20),
.B2(n_32),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_29),
.Y(n_67)
);

OR2x4_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_46),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_70),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_37),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_42),
.B1(n_53),
.B2(n_32),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_54),
.B1(n_53),
.B2(n_44),
.Y(n_88)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_80),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_31),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_41),
.A2(n_23),
.B(n_32),
.C(n_27),
.Y(n_81)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_22),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_21),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_93),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_52),
.B1(n_55),
.B2(n_27),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_70),
.B1(n_66),
.B2(n_73),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_53),
.B1(n_52),
.B2(n_38),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_89),
.A2(n_101),
.B1(n_61),
.B2(n_60),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_96),
.Y(n_115)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_52),
.B1(n_38),
.B2(n_40),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_58),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_120),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_58),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_113),
.C(n_118),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_76),
.C(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_132),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_116),
.B(n_123),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_72),
.C(n_64),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_126),
.B1(n_20),
.B2(n_18),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_90),
.B(n_57),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_68),
.A3(n_59),
.B1(n_80),
.B2(n_75),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_37),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_70),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_124),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_67),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_92),
.A2(n_60),
.B1(n_67),
.B2(n_82),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_131),
.B1(n_107),
.B2(n_101),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_85),
.A2(n_94),
.B1(n_103),
.B2(n_89),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_107),
.B1(n_102),
.B2(n_97),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_85),
.B1(n_94),
.B2(n_88),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_83),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_81),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_143),
.B1(n_144),
.B2(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_81),
.B1(n_106),
.B2(n_95),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_156),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_26),
.B(n_24),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_149),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_84),
.B1(n_106),
.B2(n_96),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_148),
.A2(n_158),
.B1(n_162),
.B2(n_133),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_155),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_93),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_120),
.B(n_25),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_84),
.C(n_37),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_161),
.C(n_129),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_38),
.B1(n_79),
.B2(n_62),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_110),
.A2(n_79),
.B1(n_20),
.B2(n_62),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_123),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_40),
.C(n_36),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_117),
.A2(n_40),
.B1(n_36),
.B2(n_26),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_144),
.B1(n_143),
.B2(n_152),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_154),
.C(n_140),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_135),
.B(n_153),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_183),
.B(n_185),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_124),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_121),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_179),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_150),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_111),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_176),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_122),
.B1(n_128),
.B2(n_112),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_177),
.B1(n_181),
.B2(n_24),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_40),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_153),
.B1(n_158),
.B2(n_148),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_36),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_184),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_SL g183 ( 
.A1(n_162),
.A2(n_36),
.B(n_1),
.C(n_2),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_26),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_9),
.B(n_15),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_0),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_191),
.B1(n_201),
.B2(n_183),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_172),
.B1(n_168),
.B2(n_180),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_138),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_186),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_197),
.C(n_182),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_149),
.B1(n_140),
.B2(n_160),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_199),
.B1(n_0),
.B2(n_1),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_139),
.C(n_159),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_24),
.B1(n_16),
.B2(n_9),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_170),
.B1(n_178),
.B2(n_174),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

AO21x1_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_24),
.B(n_9),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_185),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_208),
.B1(n_209),
.B2(n_217),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_192),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_206),
.B(n_214),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_210),
.C(n_197),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_191),
.A2(n_183),
.B1(n_179),
.B2(n_2),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_183),
.C(n_10),
.Y(n_210)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_198),
.B(n_196),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_215),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_10),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_188),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_10),
.B1(n_3),
.B2(n_5),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_224),
.C(n_194),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_186),
.C(n_190),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_190),
.C(n_194),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_205),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_232),
.C(n_223),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_226),
.A2(n_187),
.B1(n_216),
.B2(n_203),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_219),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_213),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_237),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_219),
.A2(n_211),
.B1(n_204),
.B2(n_209),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_0),
.B1(n_11),
.B2(n_13),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_217),
.B(n_201),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_236),
.B(n_218),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_222),
.A2(n_6),
.B(n_7),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_15),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_238),
.B(n_239),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_243),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_224),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_242),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_6),
.C(n_7),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_244),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_234),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_241),
.B(n_11),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_245),
.C(n_248),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_252),
.C(n_249),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_242),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_11),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_253),
.A2(n_254),
.B(n_14),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_14),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_14),
.Y(n_257)
);


endmodule