module fake_jpeg_13927_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_49),
.Y(n_69)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_43),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_47),
.B(n_51),
.C(n_29),
.Y(n_71)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_72),
.Y(n_82)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_3),
.C(n_4),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_69),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_55),
.B1(n_50),
.B2(n_39),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_79),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_87),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_56),
.B1(n_39),
.B2(n_51),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_44),
.B(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_4),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_86),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_100),
.B1(n_7),
.B2(n_11),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_75),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_96),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_5),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_44),
.C(n_77),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_44),
.C(n_8),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_6),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_6),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_107),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_108),
.B1(n_96),
.B2(n_88),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_17),
.B1(n_19),
.B2(n_23),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_110),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_92),
.B1(n_91),
.B2(n_101),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_103),
.C(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_103),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_111),
.B(n_113),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_104),
.B(n_95),
.Y(n_116)
);

OAI321xp33_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_90),
.A3(n_27),
.B1(n_31),
.B2(n_33),
.C(n_25),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_35),
.Y(n_118)
);


endmodule