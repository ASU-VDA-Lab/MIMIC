module fake_ariane_2041_n_1653 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1653);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1653;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1498;
wire n_1188;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_10),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_91),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_56),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_107),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_30),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_2),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_39),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_34),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_89),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_63),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_133),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_122),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_50),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_23),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_128),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_20),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_10),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_6),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_28),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_67),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_70),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_55),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_100),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_112),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_49),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_55),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_109),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_126),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_30),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_129),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_143),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_64),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_25),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_3),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_127),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_123),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g209 ( 
.A(n_23),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_72),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_94),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_137),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_20),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_35),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_7),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_33),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_69),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_21),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_61),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_51),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_42),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_2),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_49),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_106),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_145),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_118),
.Y(n_228)
);

BUFx2_ASAP7_75t_SL g229 ( 
.A(n_87),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_114),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_19),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_27),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_3),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_113),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_84),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_43),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_152),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_86),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_79),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_97),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_46),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_115),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_116),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_58),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_26),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_53),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_48),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_154),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_140),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_46),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_101),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_7),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_71),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_21),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_78),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_43),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_103),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_146),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_74),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_153),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_148),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_99),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_144),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_59),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_92),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_44),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_95),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_85),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_42),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_9),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_135),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_41),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_34),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_8),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_88),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_121),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_36),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_5),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_52),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_37),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_40),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_77),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_53),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_117),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_51),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_156),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_0),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_26),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_56),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_0),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_9),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_39),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_105),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_47),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_24),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_96),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_125),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_25),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_18),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_36),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_37),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_18),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_29),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_52),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_47),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_8),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_19),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_24),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_54),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_157),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_17),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_124),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_120),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_139),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_13),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_98),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_41),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_22),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_54),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_50),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_48),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_104),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_134),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_14),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_57),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_32),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_60),
.Y(n_327)
);

BUFx8_ASAP7_75t_SL g328 ( 
.A(n_33),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_269),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_328),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_301),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_R g334 ( 
.A(n_211),
.B(n_68),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_309),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_164),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_269),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_207),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_213),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_269),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_310),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_286),
.B(n_1),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_269),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_269),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_269),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_273),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_273),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_164),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_314),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_273),
.Y(n_350)
);

INVxp33_ASAP7_75t_SL g351 ( 
.A(n_161),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_195),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_199),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_273),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_273),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_214),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_215),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_273),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_196),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_216),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_273),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_266),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_219),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_193),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_182),
.B(n_1),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_273),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_221),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_285),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_285),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_163),
.B(n_4),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_232),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_285),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_285),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_208),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_285),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_222),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_161),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_168),
.B(n_4),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_167),
.B(n_5),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_288),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_288),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_236),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_241),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_247),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_250),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_252),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

NAND2xp33_ASAP7_75t_R g389 ( 
.A(n_162),
.B(n_75),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_194),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_194),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

INVxp33_ASAP7_75t_L g393 ( 
.A(n_166),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_266),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_256),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_287),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_245),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_298),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_245),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_305),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_168),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_306),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_270),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_254),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_168),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_254),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_274),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_194),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_311),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_270),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_169),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_320),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_248),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_348),
.B(n_274),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_346),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_333),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_339),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_R g421 ( 
.A(n_338),
.B(n_197),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_341),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_329),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_330),
.B(n_174),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_330),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_336),
.B(n_182),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_332),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_349),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_332),
.Y(n_431)
);

CKINVDCx8_ASAP7_75t_R g432 ( 
.A(n_364),
.Y(n_432)
);

BUFx8_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_359),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_342),
.B(n_183),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_372),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_R g440 ( 
.A(n_334),
.B(n_201),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_R g441 ( 
.A(n_352),
.B(n_203),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_331),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_374),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_319),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_353),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_367),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_335),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_362),
.B(n_319),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_412),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_343),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_R g451 ( 
.A(n_356),
.B(n_220),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_365),
.B(n_183),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_357),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_343),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_344),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_344),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_372),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_345),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_360),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_R g460 ( 
.A(n_363),
.B(n_226),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_395),
.B(n_248),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_378),
.A2(n_307),
.B1(n_169),
.B2(n_324),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_345),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_347),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_376),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_347),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_350),
.Y(n_467)
);

OA21x2_ASAP7_75t_L g468 ( 
.A1(n_350),
.A2(n_202),
.B(n_200),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_383),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_384),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_385),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_354),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_354),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_355),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_355),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_386),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_361),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_371),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_404),
.B(n_248),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_361),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_366),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_387),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_390),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_396),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_391),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_366),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_411),
.B(n_398),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_368),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_368),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_419),
.B(n_402),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_461),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_415),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_440),
.B(n_397),
.Y(n_493)
);

CKINVDCx6p67_ASAP7_75t_R g494 ( 
.A(n_435),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_417),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_428),
.B(n_351),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_419),
.B(n_406),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_452),
.A2(n_378),
.B1(n_370),
.B2(n_379),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_418),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_461),
.A2(n_377),
.B1(n_389),
.B2(n_410),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_448),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_434),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_444),
.B(n_413),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_415),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_428),
.B(n_399),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_440),
.B(n_401),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_487),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_417),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_422),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_427),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_461),
.B(n_182),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_422),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_483),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_434),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_429),
.Y(n_516)
);

NOR3xp33_ASAP7_75t_L g517 ( 
.A(n_419),
.B(n_272),
.C(n_209),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_483),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

AND3x2_ASAP7_75t_L g520 ( 
.A(n_447),
.B(n_289),
.C(n_380),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_427),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

BUFx10_ASAP7_75t_L g523 ( 
.A(n_459),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_427),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_447),
.B(n_403),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_479),
.A2(n_180),
.B1(n_283),
.B2(n_281),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_448),
.B(n_294),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_434),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_441),
.B(n_218),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_212),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_479),
.B(n_212),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_447),
.B(n_381),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_441),
.B(n_224),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_452),
.A2(n_438),
.B1(n_468),
.B2(n_448),
.Y(n_534)
);

INVxp33_ASAP7_75t_SL g535 ( 
.A(n_445),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_415),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_454),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_438),
.A2(n_185),
.B1(n_279),
.B2(n_326),
.Y(n_538)
);

NAND2x1p5_ASAP7_75t_L g539 ( 
.A(n_444),
.B(n_416),
.Y(n_539)
);

NOR3xp33_ASAP7_75t_L g540 ( 
.A(n_445),
.B(n_294),
.C(n_180),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_418),
.Y(n_541)
);

BUFx4f_ASAP7_75t_L g542 ( 
.A(n_444),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_434),
.B(n_398),
.Y(n_543)
);

INVx6_ASAP7_75t_L g544 ( 
.A(n_433),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_424),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_453),
.B(n_409),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_439),
.B(n_369),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_439),
.B(n_400),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_462),
.B(n_171),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_453),
.B(n_414),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_439),
.B(n_373),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_415),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_427),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_439),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_435),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_457),
.B(n_400),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_457),
.B(n_375),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_451),
.B(n_235),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_465),
.B(n_405),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_424),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_451),
.B(n_237),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_457),
.B(n_436),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_469),
.Y(n_564)
);

AND2x2_ASAP7_75t_SL g565 ( 
.A(n_462),
.B(n_257),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_446),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_468),
.A2(n_292),
.B1(n_295),
.B2(n_291),
.Y(n_567)
);

BUFx8_ASAP7_75t_SL g568 ( 
.A(n_442),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_456),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_457),
.B(n_405),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_460),
.B(n_239),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_463),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_457),
.B(n_375),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_463),
.Y(n_574)
);

BUFx4f_ASAP7_75t_L g575 ( 
.A(n_468),
.Y(n_575)
);

OR2x6_ASAP7_75t_L g576 ( 
.A(n_465),
.B(n_407),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_463),
.Y(n_577)
);

AND2x6_ASAP7_75t_L g578 ( 
.A(n_464),
.B(n_257),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_470),
.A2(n_281),
.B1(n_223),
.B2(n_185),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_460),
.B(n_240),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_437),
.B(n_382),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_415),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_416),
.B(n_408),
.Y(n_583)
);

BUFx8_ASAP7_75t_SL g584 ( 
.A(n_446),
.Y(n_584)
);

INVx4_ASAP7_75t_SL g585 ( 
.A(n_431),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_476),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_464),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_437),
.B(n_382),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_431),
.Y(n_589)
);

INVxp67_ASAP7_75t_SL g590 ( 
.A(n_431),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_416),
.B(n_171),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_450),
.B(n_388),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_468),
.A2(n_217),
.B1(n_321),
.B2(n_318),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_464),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_467),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_L g596 ( 
.A(n_431),
.B(n_172),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_455),
.B(n_388),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_455),
.B(n_253),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_426),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_466),
.B(n_392),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_466),
.B(n_261),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_467),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_472),
.B(n_392),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_472),
.B(n_408),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_431),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_SL g606 ( 
.A1(n_484),
.A2(n_280),
.B1(n_184),
.B2(n_278),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_471),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_468),
.A2(n_302),
.B1(n_179),
.B2(n_186),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_473),
.B(n_394),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_473),
.B(n_170),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_426),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_477),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_481),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_481),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_481),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_475),
.B(n_316),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_475),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_480),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_499),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_499),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_500),
.B(n_482),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_541),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_541),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_496),
.B(n_482),
.Y(n_625)
);

O2A1O1Ixp5_ASAP7_75t_L g626 ( 
.A1(n_528),
.A2(n_486),
.B(n_425),
.C(n_426),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_496),
.B(n_449),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_530),
.B(n_531),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_505),
.B(n_449),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_491),
.B(n_432),
.Y(n_630)
);

AND2x6_ASAP7_75t_SL g631 ( 
.A(n_546),
.B(n_187),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_512),
.A2(n_420),
.B1(n_423),
.B2(n_425),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_530),
.B(n_426),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_530),
.B(n_426),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_514),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_503),
.B(n_432),
.Y(n_636)
);

OAI22xp33_ASAP7_75t_L g637 ( 
.A1(n_526),
.A2(n_576),
.B1(n_542),
.B2(n_549),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_495),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_542),
.B(n_432),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_532),
.B(n_433),
.C(n_223),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_493),
.B(n_433),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_511),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_608),
.B(n_421),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_506),
.B(n_539),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_545),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_501),
.B(n_430),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_518),
.B(n_443),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_502),
.B(n_458),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_568),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_611),
.A2(n_489),
.B(n_488),
.C(n_191),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_560),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_SL g652 ( 
.A(n_544),
.B(n_535),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_560),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_562),
.A2(n_474),
.B(n_458),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_501),
.B(n_443),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_565),
.A2(n_489),
.B1(n_488),
.B2(n_205),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_565),
.A2(n_290),
.B1(n_206),
.B2(n_225),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_506),
.B(n_458),
.Y(n_658)
);

AO221x1_ASAP7_75t_L g659 ( 
.A1(n_507),
.A2(n_303),
.B1(n_304),
.B2(n_231),
.C(n_233),
.Y(n_659)
);

INVxp33_ASAP7_75t_L g660 ( 
.A(n_584),
.Y(n_660)
);

BUFx6f_ASAP7_75t_SL g661 ( 
.A(n_523),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_512),
.B(n_543),
.Y(n_662)
);

NOR3x1_ASAP7_75t_L g663 ( 
.A(n_525),
.B(n_299),
.C(n_300),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_512),
.B(n_474),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_501),
.B(n_162),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_555),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_544),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_543),
.B(n_474),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_498),
.A2(n_177),
.B1(n_258),
.B2(n_238),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_548),
.B(n_474),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_508),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_539),
.B(n_474),
.Y(n_672)
);

NOR2x1_ASAP7_75t_L g673 ( 
.A(n_576),
.B(n_192),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_618),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_523),
.B(n_165),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_564),
.B(n_173),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_618),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_556),
.B(n_570),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_544),
.Y(n_679)
);

NOR3xp33_ASAP7_75t_L g680 ( 
.A(n_490),
.B(n_308),
.C(n_246),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_570),
.B(n_204),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_564),
.B(n_173),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_611),
.B(n_175),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_502),
.B(n_175),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_576),
.B(n_478),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_617),
.B(n_176),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_566),
.Y(n_687)
);

O2A1O1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_619),
.A2(n_277),
.B(n_317),
.C(n_177),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_502),
.B(n_176),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_492),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_515),
.B(n_178),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_559),
.B(n_485),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_515),
.B(n_178),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_567),
.A2(n_282),
.B1(n_249),
.B2(n_320),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_509),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_586),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_550),
.B(n_478),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_515),
.B(n_181),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_509),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_617),
.B(n_189),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_510),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_504),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_504),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_554),
.B(n_189),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_536),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_510),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_536),
.Y(n_707)
);

BUFx6f_ASAP7_75t_SL g708 ( 
.A(n_586),
.Y(n_708)
);

OAI22xp33_ASAP7_75t_L g709 ( 
.A1(n_579),
.A2(n_324),
.B1(n_326),
.B2(n_325),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_497),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_552),
.Y(n_711)
);

BUFx6f_ASAP7_75t_SL g712 ( 
.A(n_586),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_585),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_567),
.A2(n_249),
.B1(n_282),
.B2(n_320),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_534),
.B(n_190),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_534),
.B(n_238),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_535),
.B(n_268),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_529),
.B(n_268),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_554),
.B(n_271),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_584),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_593),
.A2(n_282),
.B1(n_249),
.B2(n_258),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_513),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_582),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_583),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_554),
.B(n_276),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_599),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_575),
.B(n_511),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_516),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_612),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_533),
.A2(n_323),
.B1(n_322),
.B2(n_325),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_516),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_583),
.B(n_485),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_604),
.B(n_228),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_604),
.B(n_230),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_533),
.B(n_327),
.Y(n_735)
);

NAND2x1p5_ASAP7_75t_L g736 ( 
.A(n_575),
.B(n_188),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_591),
.B(n_6),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_511),
.B(n_275),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_519),
.Y(n_739)
);

HB1xp67_ASAP7_75t_SL g740 ( 
.A(n_568),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_527),
.B(n_11),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_558),
.B(n_284),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_527),
.B(n_234),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_581),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_527),
.B(n_242),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_561),
.B(n_243),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_561),
.B(n_251),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_571),
.B(n_255),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_571),
.B(n_259),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_580),
.B(n_262),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_580),
.B(n_229),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_494),
.B(n_11),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_538),
.B(n_264),
.C(n_313),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_589),
.B(n_12),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_588),
.Y(n_755)
);

AOI21x1_ASAP7_75t_L g756 ( 
.A1(n_727),
.A2(n_557),
.B(n_573),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_687),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_629),
.A2(n_569),
.B(n_616),
.C(n_563),
.Y(n_758)
);

NAND3xp33_ASAP7_75t_SL g759 ( 
.A(n_625),
.B(n_540),
.C(n_517),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_627),
.B(n_606),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_678),
.A2(n_590),
.B(n_551),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_662),
.B(n_511),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_713),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_713),
.Y(n_764)
);

OAI21xp33_ASAP7_75t_L g765 ( 
.A1(n_629),
.A2(n_598),
.B(n_601),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_655),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_670),
.A2(n_547),
.B(n_589),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_731),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_652),
.B(n_521),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_731),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_681),
.B(n_593),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_709),
.A2(n_686),
.B(n_700),
.C(n_683),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_638),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_637),
.B(n_598),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_657),
.B(n_609),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_657),
.B(n_609),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_648),
.A2(n_537),
.B(n_613),
.Y(n_777)
);

AOI21xp33_ASAP7_75t_L g778 ( 
.A1(n_718),
.A2(n_607),
.B(n_601),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_684),
.A2(n_553),
.B(n_522),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_744),
.B(n_572),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_755),
.B(n_572),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_647),
.B(n_520),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_654),
.A2(n_615),
.B(n_614),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_684),
.A2(n_522),
.B(n_521),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_644),
.B(n_521),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_667),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_656),
.B(n_574),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_689),
.A2(n_522),
.B(n_521),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_656),
.B(n_718),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_689),
.A2(n_553),
.B(n_522),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_735),
.B(n_742),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_672),
.A2(n_614),
.B(n_594),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_691),
.A2(n_553),
.B(n_605),
.Y(n_793)
);

AOI21x1_ASAP7_75t_L g794 ( 
.A1(n_727),
.A2(n_594),
.B(n_574),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_655),
.B(n_577),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_735),
.B(n_577),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_742),
.B(n_587),
.Y(n_797)
);

NOR2x1_ASAP7_75t_L g798 ( 
.A(n_639),
.B(n_592),
.Y(n_798)
);

AO21x1_ASAP7_75t_L g799 ( 
.A1(n_658),
.A2(n_610),
.B(n_603),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_692),
.B(n_587),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_644),
.B(n_595),
.Y(n_801)
);

NOR2x1_ASAP7_75t_L g802 ( 
.A(n_639),
.B(n_597),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_693),
.A2(n_605),
.B(n_553),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_698),
.A2(n_605),
.B(n_602),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_630),
.A2(n_578),
.B1(n_605),
.B2(n_585),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_704),
.A2(n_725),
.B(n_719),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_646),
.B(n_600),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_667),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_SL g809 ( 
.A1(n_754),
.A2(n_260),
.B(n_265),
.C(n_267),
.Y(n_809)
);

AOI21xp33_ASAP7_75t_L g810 ( 
.A1(n_721),
.A2(n_596),
.B(n_188),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_SL g811 ( 
.A1(n_754),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_636),
.B(n_524),
.Y(n_812)
);

OAI321xp33_ASAP7_75t_L g813 ( 
.A1(n_669),
.A2(n_172),
.A3(n_227),
.B1(n_297),
.B2(n_578),
.C(n_27),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_646),
.B(n_578),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_732),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_635),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_733),
.A2(n_293),
.B1(n_198),
.B2(n_210),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_710),
.B(n_578),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_664),
.A2(n_596),
.B(n_578),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_641),
.B(n_312),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_641),
.A2(n_244),
.B(n_198),
.C(n_293),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_630),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_690),
.A2(n_263),
.B(n_296),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_702),
.A2(n_297),
.B(n_227),
.Y(n_824)
);

O2A1O1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_650),
.A2(n_210),
.B(n_244),
.C(n_17),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_694),
.B(n_15),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_703),
.A2(n_297),
.B(n_227),
.Y(n_827)
);

AO21x1_ASAP7_75t_L g828 ( 
.A1(n_658),
.A2(n_172),
.B(n_227),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_737),
.A2(n_632),
.B(n_694),
.C(n_714),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_714),
.B(n_15),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_679),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_740),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_734),
.A2(n_172),
.B1(n_22),
.B2(n_28),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_705),
.A2(n_172),
.B(n_90),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_620),
.B(n_16),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_621),
.B(n_16),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_707),
.A2(n_93),
.B(n_155),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_623),
.B(n_31),
.Y(n_838)
);

O2A1O1Ixp5_ASAP7_75t_L g839 ( 
.A1(n_738),
.A2(n_32),
.B(n_35),
.C(n_38),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_685),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_711),
.A2(n_119),
.B(n_151),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_624),
.B(n_38),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_645),
.B(n_651),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_723),
.A2(n_83),
.B(n_138),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_642),
.B(n_44),
.Y(n_845)
);

CKINVDCx10_ASAP7_75t_R g846 ( 
.A(n_661),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_679),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_653),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_680),
.B(n_45),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_SL g850 ( 
.A1(n_685),
.A2(n_45),
.B1(n_62),
.B2(n_65),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_696),
.B(n_66),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_726),
.A2(n_73),
.B(n_76),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_696),
.B(n_80),
.Y(n_853)
);

BUFx8_ASAP7_75t_L g854 ( 
.A(n_661),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_642),
.B(n_82),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_649),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_674),
.A2(n_130),
.B1(n_136),
.B2(n_158),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_677),
.B(n_741),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_666),
.B(n_685),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_751),
.B(n_729),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_642),
.Y(n_861)
);

AOI21xp33_ASAP7_75t_L g862 ( 
.A1(n_751),
.A2(n_716),
.B(n_715),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_751),
.B(n_622),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_628),
.A2(n_753),
.B1(n_642),
.B2(n_634),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_743),
.B(n_745),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_708),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_747),
.B(n_750),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_633),
.A2(n_728),
.B(n_739),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_697),
.B(n_720),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_697),
.B(n_673),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_671),
.A2(n_695),
.B(n_722),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_699),
.A2(n_701),
.B(n_706),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_697),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_749),
.B(n_730),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_665),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_701),
.B(n_746),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_643),
.B(n_663),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_688),
.A2(n_640),
.B(n_748),
.C(n_682),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_736),
.A2(n_676),
.B(n_675),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_717),
.A2(n_659),
.B(n_752),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_708),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_660),
.A2(n_629),
.B(n_496),
.C(n_625),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_712),
.A2(n_626),
.B(n_678),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_631),
.B(n_712),
.Y(n_884)
);

OAI321xp33_ASAP7_75t_L g885 ( 
.A1(n_625),
.A2(n_627),
.A3(n_669),
.B1(n_657),
.B2(n_714),
.C(n_694),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_678),
.A2(n_670),
.B(n_668),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_626),
.A2(n_678),
.B(n_575),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_678),
.A2(n_670),
.B(n_668),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_678),
.A2(n_670),
.B(n_668),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_678),
.A2(n_670),
.B(n_668),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_649),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_655),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_629),
.B(n_625),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_629),
.B(n_625),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_724),
.B(n_696),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_629),
.A2(n_625),
.B1(n_496),
.B2(n_627),
.Y(n_896)
);

BUFx12f_ASAP7_75t_L g897 ( 
.A(n_685),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_678),
.A2(n_670),
.B(n_668),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_626),
.A2(n_678),
.B(n_575),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_886),
.A2(n_889),
.B(n_888),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_896),
.A2(n_774),
.B1(n_894),
.B2(n_893),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_794),
.A2(n_868),
.B(n_783),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_774),
.A2(n_822),
.B1(n_760),
.B2(n_759),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_786),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_890),
.A2(n_898),
.B(n_887),
.Y(n_905)
);

NOR2xp67_ASAP7_75t_L g906 ( 
.A(n_816),
.B(n_822),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_899),
.A2(n_761),
.B(n_767),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_786),
.Y(n_908)
);

NOR2x1_ASAP7_75t_SL g909 ( 
.A(n_763),
.B(n_764),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_800),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_791),
.B(n_789),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_815),
.B(n_766),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_775),
.B(n_776),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_872),
.A2(n_784),
.B(n_779),
.Y(n_914)
);

AOI21xp33_ASAP7_75t_L g915 ( 
.A1(n_885),
.A2(n_772),
.B(n_760),
.Y(n_915)
);

BUFx10_ASAP7_75t_L g916 ( 
.A(n_832),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_SL g917 ( 
.A(n_829),
.B(n_850),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_763),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_882),
.B(n_865),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_788),
.A2(n_793),
.B(n_790),
.Y(n_920)
);

NOR2x1_ASAP7_75t_L g921 ( 
.A(n_856),
.B(n_866),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_786),
.Y(n_922)
);

BUFx10_ASAP7_75t_L g923 ( 
.A(n_851),
.Y(n_923)
);

OAI21x1_ASAP7_75t_L g924 ( 
.A1(n_803),
.A2(n_804),
.B(n_792),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_871),
.A2(n_756),
.B(n_762),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_777),
.A2(n_758),
.B(n_762),
.Y(n_926)
);

OR2x6_ASAP7_75t_L g927 ( 
.A(n_869),
.B(n_892),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_882),
.B(n_795),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_757),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_L g930 ( 
.A1(n_765),
.A2(n_759),
.B(n_830),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_801),
.B(n_771),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_786),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_757),
.B(n_859),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_847),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_874),
.A2(n_826),
.B(n_801),
.C(n_812),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_780),
.B(n_781),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_858),
.A2(n_878),
.B1(n_787),
.B2(n_875),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_878),
.A2(n_875),
.B1(n_842),
.B2(n_835),
.Y(n_938)
);

OAI21x1_ASAP7_75t_L g939 ( 
.A1(n_785),
.A2(n_864),
.B(n_819),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_847),
.Y(n_940)
);

OAI22xp33_ASAP7_75t_L g941 ( 
.A1(n_869),
.A2(n_813),
.B1(n_873),
.B2(n_849),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_847),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_836),
.A2(n_838),
.B1(n_820),
.B2(n_851),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_867),
.B(n_812),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_895),
.B(n_853),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_843),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_796),
.B(n_797),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_895),
.B(n_853),
.Y(n_948)
);

NOR2xp67_ASAP7_75t_L g949 ( 
.A(n_816),
.B(n_881),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_825),
.A2(n_778),
.B(n_880),
.C(n_879),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_891),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_807),
.B(n_863),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_839),
.A2(n_827),
.B(n_824),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_834),
.A2(n_855),
.B(n_852),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_845),
.A2(n_860),
.B1(n_833),
.B2(n_821),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_798),
.A2(n_802),
.B(n_855),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_845),
.A2(n_805),
.B1(n_848),
.B2(n_876),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_831),
.B(n_808),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_768),
.A2(n_770),
.B1(n_769),
.B2(n_873),
.Y(n_959)
);

OAI21x1_ASAP7_75t_SL g960 ( 
.A1(n_837),
.A2(n_844),
.B(n_841),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_861),
.A2(n_823),
.B(n_809),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_861),
.A2(n_828),
.B(n_857),
.Y(n_962)
);

AOI221xp5_ASAP7_75t_L g963 ( 
.A1(n_877),
.A2(n_811),
.B1(n_782),
.B2(n_817),
.C(n_810),
.Y(n_963)
);

AO21x1_ASAP7_75t_L g964 ( 
.A1(n_809),
.A2(n_818),
.B(n_831),
.Y(n_964)
);

OA22x2_ASAP7_75t_L g965 ( 
.A1(n_869),
.A2(n_840),
.B1(n_870),
.B2(n_884),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_847),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_897),
.B(n_866),
.Y(n_967)
);

AO22x1_ASAP7_75t_L g968 ( 
.A1(n_854),
.A2(n_763),
.B1(n_764),
.B2(n_846),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_854),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_786),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_886),
.A2(n_678),
.B(n_888),
.Y(n_971)
);

OAI21x1_ASAP7_75t_SL g972 ( 
.A1(n_883),
.A2(n_879),
.B(n_806),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_893),
.B(n_894),
.Y(n_973)
);

AOI21x1_ASAP7_75t_L g974 ( 
.A1(n_794),
.A2(n_868),
.B(n_762),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_886),
.A2(n_678),
.B(n_888),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_886),
.A2(n_678),
.B(n_888),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_893),
.B(n_894),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_896),
.B(n_503),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_886),
.A2(n_678),
.B(n_888),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_814),
.B(n_795),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_886),
.A2(n_678),
.B(n_888),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_896),
.B(n_503),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_822),
.B(n_652),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_886),
.A2(n_678),
.B(n_888),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_896),
.B(n_503),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_763),
.Y(n_986)
);

AND2x2_ASAP7_75t_SL g987 ( 
.A(n_774),
.B(n_641),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_886),
.A2(n_678),
.B(n_888),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_L g989 ( 
.A(n_816),
.B(n_635),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_893),
.B(n_894),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_763),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_757),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_893),
.B(n_894),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_896),
.A2(n_894),
.B1(n_893),
.B2(n_789),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_886),
.A2(n_678),
.B(n_888),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_893),
.B(n_894),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_773),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_886),
.A2(n_678),
.B(n_888),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_773),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_800),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_822),
.B(n_652),
.Y(n_1001)
);

AO21x2_ASAP7_75t_L g1002 ( 
.A1(n_862),
.A2(n_799),
.B(n_828),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_773),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_832),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_763),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_869),
.B(n_685),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_896),
.A2(n_894),
.B1(n_893),
.B2(n_789),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_893),
.B(n_894),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_794),
.A2(n_868),
.B(n_783),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_887),
.A2(n_899),
.B(n_888),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_854),
.Y(n_1011)
);

OAI22x1_ASAP7_75t_L g1012 ( 
.A1(n_896),
.A2(n_774),
.B1(n_873),
.B2(n_462),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_794),
.A2(n_868),
.B(n_783),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_794),
.A2(n_868),
.B(n_783),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_854),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_786),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_896),
.A2(n_535),
.B1(n_774),
.B2(n_629),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_893),
.B(n_894),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_L g1019 ( 
.A1(n_794),
.A2(n_868),
.B(n_762),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_910),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_971),
.A2(n_976),
.B(n_975),
.Y(n_1021)
);

BUFx2_ASAP7_75t_SL g1022 ( 
.A(n_951),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_901),
.B(n_994),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_979),
.A2(n_984),
.B(n_981),
.Y(n_1024)
);

AOI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_987),
.A2(n_917),
.B(n_915),
.Y(n_1025)
);

CKINVDCx6p67_ASAP7_75t_R g1026 ( 
.A(n_1011),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_916),
.Y(n_1027)
);

AOI21xp33_ASAP7_75t_L g1028 ( 
.A1(n_917),
.A2(n_915),
.B(n_994),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_L g1029 ( 
.A(n_1017),
.B(n_903),
.C(n_1007),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_912),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_980),
.B(n_945),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_988),
.A2(n_998),
.B(n_995),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_SL g1033 ( 
.A1(n_943),
.A2(n_911),
.B(n_931),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1000),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1007),
.B(n_973),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_973),
.B(n_977),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_1012),
.A2(n_978),
.B1(n_982),
.B2(n_985),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_933),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_977),
.B(n_990),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_990),
.B(n_996),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_929),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_997),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_980),
.B(n_948),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_999),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_996),
.B(n_1008),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_919),
.A2(n_930),
.B(n_1008),
.C(n_943),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_927),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_993),
.A2(n_1018),
.B(n_938),
.C(n_950),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_927),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1003),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_904),
.Y(n_1051)
);

CKINVDCx16_ASAP7_75t_R g1052 ( 
.A(n_1015),
.Y(n_1052)
);

CKINVDCx8_ASAP7_75t_R g1053 ( 
.A(n_967),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_929),
.B(n_992),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_916),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_927),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_1004),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_911),
.A2(n_928),
.B1(n_931),
.B2(n_936),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_936),
.A2(n_938),
.B1(n_935),
.B2(n_944),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_992),
.B(n_1006),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_944),
.B(n_913),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_906),
.A2(n_983),
.B1(n_1001),
.B2(n_941),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_923),
.B(n_963),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_958),
.B(n_967),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_937),
.B(n_958),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_913),
.B(n_947),
.Y(n_1066)
);

BUFx8_ASAP7_75t_SL g1067 ( 
.A(n_967),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_904),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_946),
.A2(n_937),
.B1(n_947),
.B2(n_955),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_968),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_965),
.A2(n_1006),
.B1(n_952),
.B2(n_955),
.Y(n_1071)
);

AO21x1_ASAP7_75t_L g1072 ( 
.A1(n_957),
.A2(n_959),
.B(n_956),
.Y(n_1072)
);

AOI222xp33_ASAP7_75t_L g1073 ( 
.A1(n_969),
.A2(n_989),
.B1(n_957),
.B2(n_949),
.C1(n_959),
.C2(n_1010),
.Y(n_1073)
);

NAND2xp33_ASAP7_75t_L g1074 ( 
.A(n_908),
.B(n_934),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_908),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_1006),
.B(n_934),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_932),
.B(n_966),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_908),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_921),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_922),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_922),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_922),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_934),
.Y(n_1083)
);

INVx8_ASAP7_75t_L g1084 ( 
.A(n_940),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_940),
.B(n_942),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_940),
.B(n_942),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_965),
.A2(n_1002),
.B1(n_1016),
.B2(n_970),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_966),
.B(n_970),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_966),
.Y(n_1089)
);

AOI21xp33_ASAP7_75t_L g1090 ( 
.A1(n_1002),
.A2(n_972),
.B(n_926),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_SL g1091 ( 
.A1(n_964),
.A2(n_961),
.B(n_960),
.Y(n_1091)
);

BUFx12f_ASAP7_75t_L g1092 ( 
.A(n_970),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1016),
.B(n_991),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_1016),
.B(n_932),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_918),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_986),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_986),
.B(n_991),
.Y(n_1097)
);

OR2x6_ASAP7_75t_SL g1098 ( 
.A(n_909),
.B(n_1005),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_953),
.A2(n_939),
.B1(n_925),
.B2(n_962),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_974),
.B(n_1019),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_953),
.A2(n_954),
.B(n_924),
.C(n_920),
.Y(n_1101)
);

INVxp67_ASAP7_75t_SL g1102 ( 
.A(n_902),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_914),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_1009),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1013),
.B(n_1014),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_901),
.B(n_994),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_901),
.B(n_994),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_971),
.A2(n_976),
.B(n_975),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_929),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_904),
.Y(n_1110)
);

INVx3_ASAP7_75t_SL g1111 ( 
.A(n_951),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_971),
.A2(n_976),
.B(n_975),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_933),
.B(n_978),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_951),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_904),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_971),
.A2(n_976),
.B(n_975),
.Y(n_1116)
);

AND2x6_ASAP7_75t_L g1117 ( 
.A(n_903),
.B(n_774),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_901),
.B(n_994),
.Y(n_1118)
);

BUFx12f_ASAP7_75t_L g1119 ( 
.A(n_916),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_951),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_933),
.B(n_978),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_980),
.B(n_945),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_951),
.Y(n_1123)
);

BUFx12f_ASAP7_75t_L g1124 ( 
.A(n_916),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_901),
.B(n_994),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_901),
.B(n_994),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_951),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_916),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_971),
.A2(n_976),
.B(n_975),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_933),
.B(n_978),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_951),
.Y(n_1131)
);

CKINVDCx16_ASAP7_75t_R g1132 ( 
.A(n_951),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1017),
.A2(n_535),
.B1(n_917),
.B2(n_987),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_933),
.B(n_978),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_904),
.Y(n_1135)
);

BUFx12f_ASAP7_75t_L g1136 ( 
.A(n_916),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_971),
.A2(n_976),
.B(n_975),
.Y(n_1137)
);

OA21x2_ASAP7_75t_L g1138 ( 
.A1(n_907),
.A2(n_905),
.B(n_900),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_901),
.A2(n_919),
.B(n_772),
.C(n_903),
.Y(n_1139)
);

INVx5_ASAP7_75t_L g1140 ( 
.A(n_923),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_951),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_904),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_994),
.A2(n_893),
.B(n_894),
.C(n_882),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_971),
.A2(n_976),
.B(n_975),
.Y(n_1144)
);

OA21x2_ASAP7_75t_L g1145 ( 
.A1(n_907),
.A2(n_905),
.B(n_900),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_916),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_901),
.A2(n_1017),
.B1(n_896),
.B2(n_893),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_971),
.A2(n_976),
.B(n_975),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_980),
.B(n_945),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1039),
.B(n_1036),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1042),
.Y(n_1151)
);

BUFx12f_ASAP7_75t_L g1152 ( 
.A(n_1127),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1044),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1133),
.A2(n_1029),
.B1(n_1147),
.B2(n_1107),
.Y(n_1154)
);

BUFx4f_ASAP7_75t_SL g1155 ( 
.A(n_1120),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1050),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1113),
.B(n_1121),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_1132),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1020),
.Y(n_1159)
);

OAI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1025),
.A2(n_1147),
.B1(n_1106),
.B2(n_1023),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1112),
.A2(n_1144),
.B(n_1129),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1117),
.A2(n_1025),
.B1(n_1028),
.B2(n_1037),
.Y(n_1162)
);

AO21x1_ASAP7_75t_L g1163 ( 
.A1(n_1028),
.A2(n_1069),
.B(n_1059),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_1054),
.Y(n_1164)
);

CKINVDCx11_ASAP7_75t_R g1165 ( 
.A(n_1111),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1041),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1139),
.A2(n_1143),
.B(n_1046),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1117),
.A2(n_1062),
.B1(n_1063),
.B2(n_1073),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1109),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1081),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1036),
.B(n_1040),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1040),
.B(n_1045),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1045),
.B(n_1035),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1034),
.Y(n_1174)
);

INVx1_ASAP7_75t_SL g1175 ( 
.A(n_1022),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1067),
.Y(n_1176)
);

BUFx12f_ASAP7_75t_L g1177 ( 
.A(n_1057),
.Y(n_1177)
);

INVxp33_ASAP7_75t_L g1178 ( 
.A(n_1130),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1084),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1112),
.A2(n_1129),
.B(n_1148),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1134),
.B(n_1038),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1117),
.A2(n_1106),
.B1(n_1023),
.B2(n_1107),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1080),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_1030),
.B(n_1060),
.Y(n_1184)
);

AO21x2_ASAP7_75t_L g1185 ( 
.A1(n_1090),
.A2(n_1091),
.B(n_1024),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_SL g1186 ( 
.A1(n_1117),
.A2(n_1118),
.B1(n_1125),
.B2(n_1126),
.Y(n_1186)
);

INVx6_ASAP7_75t_L g1187 ( 
.A(n_1092),
.Y(n_1187)
);

CKINVDCx11_ASAP7_75t_R g1188 ( 
.A(n_1026),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1035),
.B(n_1066),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1078),
.Y(n_1190)
);

INVx4_ASAP7_75t_SL g1191 ( 
.A(n_1117),
.Y(n_1191)
);

AO21x2_ASAP7_75t_L g1192 ( 
.A1(n_1090),
.A2(n_1021),
.B(n_1137),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1118),
.A2(n_1126),
.B1(n_1125),
.B2(n_1069),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1032),
.A2(n_1116),
.B(n_1108),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1048),
.A2(n_1059),
.B(n_1033),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1080),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1131),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1114),
.B(n_1123),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1058),
.A2(n_1073),
.B(n_1065),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1096),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1058),
.A2(n_1071),
.B1(n_1066),
.B2(n_1061),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1097),
.Y(n_1202)
);

CKINVDCx11_ASAP7_75t_R g1203 ( 
.A(n_1053),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1105),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1082),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_1052),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1061),
.A2(n_1031),
.B1(n_1122),
.B2(n_1043),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1097),
.Y(n_1208)
);

BUFx12f_ASAP7_75t_L g1209 ( 
.A(n_1119),
.Y(n_1209)
);

BUFx4f_ASAP7_75t_SL g1210 ( 
.A(n_1124),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1149),
.A2(n_1072),
.B1(n_1070),
.B2(n_1047),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_1085),
.Y(n_1212)
);

OAI22xp33_ASAP7_75t_R g1213 ( 
.A1(n_1128),
.A2(n_1141),
.B1(n_1146),
.B2(n_1136),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1105),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1093),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1049),
.B(n_1056),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1027),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1093),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1088),
.B(n_1089),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1085),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1051),
.B(n_1135),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1140),
.A2(n_1055),
.B1(n_1079),
.B2(n_1098),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1051),
.B(n_1135),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1086),
.Y(n_1224)
);

INVxp67_ASAP7_75t_L g1225 ( 
.A(n_1086),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1140),
.A2(n_1068),
.B1(n_1083),
.B2(n_1095),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1075),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1075),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1110),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1101),
.A2(n_1099),
.B(n_1138),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1100),
.A2(n_1104),
.B(n_1102),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1087),
.A2(n_1145),
.B1(n_1094),
.B2(n_1110),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1103),
.A2(n_1074),
.B(n_1095),
.Y(n_1233)
);

BUFx4f_ASAP7_75t_SL g1234 ( 
.A(n_1115),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_1115),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1142),
.Y(n_1236)
);

BUFx2_ASAP7_75t_R g1237 ( 
.A(n_1077),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1142),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1054),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1042),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_SL g1241 ( 
.A1(n_1117),
.A2(n_917),
.B1(n_987),
.B2(n_433),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1113),
.B(n_1121),
.Y(n_1242)
);

INVx6_ASAP7_75t_L g1243 ( 
.A(n_1092),
.Y(n_1243)
);

CKINVDCx11_ASAP7_75t_R g1244 ( 
.A(n_1120),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1081),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1092),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1064),
.Y(n_1247)
);

INVx6_ASAP7_75t_L g1248 ( 
.A(n_1092),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1076),
.B(n_1081),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_1081),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1113),
.B(n_1121),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1076),
.B(n_1081),
.Y(n_1252)
);

OAI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1133),
.A2(n_917),
.B1(n_1017),
.B2(n_903),
.Y(n_1253)
);

AO21x1_ASAP7_75t_L g1254 ( 
.A1(n_1025),
.A2(n_917),
.B(n_915),
.Y(n_1254)
);

NAND3xp33_ASAP7_75t_SL g1255 ( 
.A(n_1133),
.B(n_1017),
.C(n_896),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1113),
.B(n_1121),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1147),
.B(n_1017),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1042),
.Y(n_1258)
);

OA21x2_ASAP7_75t_L g1259 ( 
.A1(n_1161),
.A2(n_1180),
.B(n_1194),
.Y(n_1259)
);

AND2x2_ASAP7_75t_SL g1260 ( 
.A(n_1168),
.B(n_1162),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1164),
.B(n_1239),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1182),
.B(n_1186),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1182),
.B(n_1204),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1157),
.B(n_1242),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1233),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1251),
.B(n_1256),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1244),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1204),
.B(n_1214),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1220),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1202),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1208),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1166),
.B(n_1169),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1155),
.B(n_1244),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1191),
.B(n_1178),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1200),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1233),
.Y(n_1276)
);

INVx5_ASAP7_75t_L g1277 ( 
.A(n_1245),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1205),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1159),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1199),
.B(n_1181),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1219),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1249),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1257),
.B(n_1193),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1257),
.B(n_1195),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1174),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1230),
.A2(n_1163),
.B(n_1167),
.Y(n_1286)
);

NOR2x1_ASAP7_75t_L g1287 ( 
.A(n_1222),
.B(n_1226),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1192),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1184),
.B(n_1173),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1151),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1153),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1156),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1230),
.A2(n_1231),
.B(n_1232),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1185),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1240),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1258),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1185),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1189),
.B(n_1160),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1212),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1225),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1215),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1218),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1224),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1171),
.B(n_1172),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1201),
.B(n_1162),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1201),
.B(n_1154),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1254),
.A2(n_1253),
.B(n_1255),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1150),
.B(n_1211),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1252),
.B(n_1232),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_SL g1310 ( 
.A(n_1237),
.B(n_1250),
.Y(n_1310)
);

AOI211xp5_ASAP7_75t_L g1311 ( 
.A1(n_1213),
.A2(n_1175),
.B(n_1198),
.C(n_1241),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1227),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1228),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1229),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1207),
.B(n_1236),
.Y(n_1315)
);

CKINVDCx14_ASAP7_75t_R g1316 ( 
.A(n_1176),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1238),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1284),
.B(n_1197),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1261),
.B(n_1216),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1284),
.B(n_1197),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1276),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1286),
.B(n_1221),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1299),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1286),
.B(n_1221),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1286),
.B(n_1221),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1298),
.B(n_1196),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1283),
.B(n_1306),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1298),
.B(n_1299),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1270),
.B(n_1271),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1286),
.B(n_1223),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1270),
.B(n_1196),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1275),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1261),
.B(n_1247),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1275),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1263),
.B(n_1190),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1279),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1279),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1285),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1271),
.B(n_1183),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1285),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1282),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1278),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1272),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1263),
.B(n_1190),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1283),
.B(n_1235),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1259),
.Y(n_1346)
);

INVx4_ASAP7_75t_L g1347 ( 
.A(n_1277),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1304),
.B(n_1170),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1276),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1272),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1306),
.B(n_1165),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1351),
.B(n_1165),
.Y(n_1352)
);

NAND3xp33_ASAP7_75t_L g1353 ( 
.A(n_1328),
.B(n_1311),
.C(n_1305),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1328),
.B(n_1300),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1351),
.A2(n_1260),
.B1(n_1305),
.B2(n_1262),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1318),
.B(n_1264),
.Y(n_1356)
);

NAND4xp25_ASAP7_75t_L g1357 ( 
.A(n_1326),
.B(n_1311),
.C(n_1273),
.D(n_1262),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1343),
.B(n_1281),
.Y(n_1358)
);

NAND4xp25_ASAP7_75t_L g1359 ( 
.A(n_1326),
.B(n_1280),
.C(n_1314),
.D(n_1313),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1318),
.B(n_1320),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1327),
.A2(n_1260),
.B(n_1287),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1343),
.B(n_1281),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1350),
.B(n_1289),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1327),
.A2(n_1260),
.B1(n_1307),
.B2(n_1308),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1318),
.B(n_1264),
.Y(n_1365)
);

OAI221xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1335),
.A2(n_1308),
.B1(n_1280),
.B2(n_1304),
.C(n_1265),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1350),
.B(n_1348),
.Y(n_1367)
);

NAND3xp33_ASAP7_75t_L g1368 ( 
.A(n_1342),
.B(n_1303),
.C(n_1301),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_SL g1369 ( 
.A1(n_1320),
.A2(n_1287),
.B(n_1321),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1342),
.B(n_1269),
.Y(n_1370)
);

OAI221xp5_ASAP7_75t_L g1371 ( 
.A1(n_1335),
.A2(n_1291),
.B1(n_1295),
.B2(n_1292),
.C(n_1296),
.Y(n_1371)
);

NAND3xp33_ASAP7_75t_L g1372 ( 
.A(n_1323),
.B(n_1303),
.C(n_1301),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1322),
.B(n_1266),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1319),
.B(n_1267),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1344),
.A2(n_1307),
.B1(n_1309),
.B2(n_1315),
.Y(n_1375)
);

AOI221xp5_ASAP7_75t_L g1376 ( 
.A1(n_1345),
.A2(n_1295),
.B1(n_1292),
.B2(n_1291),
.C(n_1290),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1323),
.B(n_1302),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1344),
.A2(n_1333),
.B1(n_1158),
.B2(n_1319),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1322),
.B(n_1293),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1344),
.A2(n_1158),
.B1(n_1206),
.B2(n_1217),
.Y(n_1380)
);

NAND3xp33_ASAP7_75t_L g1381 ( 
.A(n_1339),
.B(n_1302),
.C(n_1317),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1319),
.B(n_1307),
.Y(n_1382)
);

OAI21xp33_ASAP7_75t_L g1383 ( 
.A1(n_1339),
.A2(n_1314),
.B(n_1313),
.Y(n_1383)
);

NAND3xp33_ASAP7_75t_L g1384 ( 
.A(n_1331),
.B(n_1317),
.C(n_1345),
.Y(n_1384)
);

AND2x2_ASAP7_75t_SL g1385 ( 
.A(n_1321),
.B(n_1265),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1333),
.B(n_1268),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1333),
.B(n_1307),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1329),
.B(n_1290),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1329),
.B(n_1296),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1321),
.A2(n_1316),
.B(n_1274),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1332),
.B(n_1312),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1324),
.B(n_1293),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1324),
.B(n_1294),
.C(n_1297),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1346),
.B(n_1312),
.C(n_1288),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1391),
.Y(n_1395)
);

AND2x4_ASAP7_75t_SL g1396 ( 
.A(n_1360),
.B(n_1347),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1373),
.B(n_1349),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1377),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1382),
.B(n_1332),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1360),
.B(n_1324),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1383),
.B(n_1334),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1381),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1386),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1367),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1394),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1356),
.B(n_1325),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1356),
.B(n_1325),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1376),
.B(n_1334),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1385),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1386),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1363),
.B(n_1358),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1365),
.B(n_1325),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1365),
.B(n_1330),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1388),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1362),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1354),
.B(n_1336),
.Y(n_1417)
);

NAND2x1p5_ASAP7_75t_L g1418 ( 
.A(n_1385),
.B(n_1347),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1389),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1368),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1394),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1379),
.B(n_1330),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1372),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1379),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1384),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1392),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1384),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1392),
.B(n_1330),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1393),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1370),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1425),
.B(n_1369),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1396),
.B(n_1341),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1402),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1426),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1410),
.B(n_1374),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1403),
.A2(n_1353),
.B1(n_1361),
.B2(n_1355),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1410),
.B(n_1390),
.Y(n_1437)
);

NAND2x1_ASAP7_75t_L g1438 ( 
.A(n_1397),
.B(n_1347),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1402),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1426),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1395),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1395),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1404),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1407),
.B(n_1378),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1420),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1425),
.B(n_1337),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1426),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1427),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1407),
.B(n_1341),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1396),
.B(n_1341),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1407),
.B(n_1341),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1403),
.A2(n_1364),
.B1(n_1366),
.B2(n_1375),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1416),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1406),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1427),
.B(n_1420),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1423),
.B(n_1338),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1406),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1423),
.B(n_1338),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1405),
.B(n_1359),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1405),
.B(n_1371),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1415),
.B(n_1340),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1418),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1406),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1409),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1404),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1408),
.B(n_1380),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1416),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1411),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1411),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1408),
.B(n_1352),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1455),
.B(n_1400),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1432),
.Y(n_1472)
);

NAND2x2_ASAP7_75t_L g1473 ( 
.A(n_1431),
.B(n_1430),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1432),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1455),
.B(n_1400),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1456),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1456),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1445),
.B(n_1409),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1437),
.B(n_1408),
.Y(n_1479)
);

NOR2xp67_ASAP7_75t_L g1480 ( 
.A(n_1462),
.B(n_1429),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1435),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1435),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1445),
.B(n_1399),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1437),
.B(n_1470),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1464),
.B(n_1415),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1462),
.B(n_1396),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1443),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1470),
.B(n_1413),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1460),
.B(n_1399),
.Y(n_1489)
);

INVxp67_ASAP7_75t_SL g1490 ( 
.A(n_1464),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1444),
.B(n_1413),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1444),
.B(n_1413),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1434),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1460),
.B(n_1412),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1458),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1443),
.B(n_1412),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1448),
.B(n_1419),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1434),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1465),
.B(n_1417),
.Y(n_1499)
);

NOR2x1_ASAP7_75t_L g1500 ( 
.A(n_1431),
.B(n_1206),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1448),
.B(n_1419),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1458),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1453),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1467),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1434),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1466),
.B(n_1432),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1446),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1446),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1466),
.B(n_1414),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1459),
.B(n_1176),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1461),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1461),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1465),
.Y(n_1513)
);

INVx3_ASAP7_75t_SL g1514 ( 
.A(n_1481),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1490),
.B(n_1436),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1487),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1482),
.B(n_1436),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1500),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1471),
.B(n_1475),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1484),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1484),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1506),
.B(n_1454),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1493),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1487),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1493),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1494),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1478),
.B(n_1433),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1498),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1498),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1503),
.B(n_1433),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1513),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1504),
.B(n_1439),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1485),
.B(n_1439),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1506),
.B(n_1454),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1499),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1494),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1499),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1496),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1496),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1509),
.B(n_1462),
.Y(n_1540)
);

AOI22x1_ASAP7_75t_L g1541 ( 
.A1(n_1472),
.A2(n_1462),
.B1(n_1152),
.B2(n_1177),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1510),
.B(n_1209),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1473),
.A2(n_1452),
.B1(n_1429),
.B2(n_1463),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1473),
.A2(n_1452),
.B1(n_1429),
.B2(n_1463),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_L g1545 ( 
.A(n_1471),
.B(n_1438),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1483),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_SL g1547 ( 
.A(n_1486),
.B(n_1432),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1497),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1483),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1514),
.B(n_1509),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1515),
.A2(n_1480),
.B(n_1475),
.Y(n_1551)
);

OAI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1543),
.A2(n_1454),
.B1(n_1457),
.B2(n_1463),
.C(n_1489),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1526),
.B(n_1491),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1514),
.B(n_1491),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1536),
.B(n_1501),
.Y(n_1555)
);

NAND3xp33_ASAP7_75t_L g1556 ( 
.A(n_1544),
.B(n_1457),
.C(n_1476),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1517),
.A2(n_1459),
.B1(n_1474),
.B2(n_1472),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1518),
.A2(n_1457),
.B(n_1489),
.Y(n_1558)
);

AOI31xp33_ASAP7_75t_L g1559 ( 
.A1(n_1549),
.A2(n_1474),
.A3(n_1479),
.B(n_1492),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1546),
.B(n_1549),
.Y(n_1560)
);

AOI221xp5_ASAP7_75t_L g1561 ( 
.A1(n_1548),
.A2(n_1477),
.B1(n_1495),
.B2(n_1502),
.C(n_1508),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1546),
.Y(n_1562)
);

OAI32xp33_ASAP7_75t_L g1563 ( 
.A1(n_1519),
.A2(n_1507),
.A3(n_1479),
.B1(n_1511),
.B2(n_1512),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1516),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1514),
.B(n_1492),
.Y(n_1565)
);

A2O1A1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1527),
.A2(n_1421),
.B(n_1357),
.C(n_1505),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1520),
.A2(n_1488),
.B1(n_1418),
.B2(n_1486),
.Y(n_1567)
);

A2O1A1Ixp33_ASAP7_75t_L g1568 ( 
.A1(n_1548),
.A2(n_1421),
.B(n_1505),
.C(n_1486),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1520),
.A2(n_1488),
.B1(n_1418),
.B2(n_1424),
.Y(n_1569)
);

AOI221xp5_ASAP7_75t_L g1570 ( 
.A1(n_1538),
.A2(n_1421),
.B1(n_1441),
.B2(n_1442),
.C(n_1469),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1521),
.Y(n_1571)
);

O2A1O1Ixp33_ASAP7_75t_L g1572 ( 
.A1(n_1538),
.A2(n_1424),
.B(n_1442),
.C(n_1441),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1516),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1522),
.A2(n_1469),
.B1(n_1468),
.B2(n_1440),
.Y(n_1574)
);

AOI211xp5_ASAP7_75t_L g1575 ( 
.A1(n_1519),
.A2(n_1522),
.B(n_1534),
.C(n_1539),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1552),
.A2(n_1522),
.B1(n_1534),
.B2(n_1528),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1562),
.B(n_1521),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1550),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_SL g1579 ( 
.A1(n_1562),
.A2(n_1542),
.B1(n_1522),
.B2(n_1534),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1554),
.B(n_1547),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1565),
.B(n_1571),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1560),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1575),
.B(n_1534),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1553),
.B(n_1539),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1558),
.B(n_1535),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1564),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1555),
.B(n_1535),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1558),
.B(n_1537),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1559),
.B(n_1537),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1573),
.B(n_1530),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1557),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1556),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1572),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1566),
.B(n_1532),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1551),
.B(n_1540),
.Y(n_1595)
);

OAI31xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1592),
.A2(n_1545),
.A3(n_1561),
.B(n_1570),
.Y(n_1596)
);

AOI211xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1582),
.A2(n_1568),
.B(n_1567),
.C(n_1210),
.Y(n_1597)
);

NAND5xp2_ASAP7_75t_SL g1598 ( 
.A(n_1583),
.B(n_1572),
.C(n_1563),
.D(n_1540),
.E(n_1574),
.Y(n_1598)
);

OAI32xp33_ASAP7_75t_L g1599 ( 
.A1(n_1594),
.A2(n_1533),
.A3(n_1524),
.B1(n_1569),
.B2(n_1531),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1578),
.B(n_1531),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1585),
.A2(n_1545),
.B(n_1524),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1592),
.A2(n_1529),
.B1(n_1528),
.B2(n_1525),
.C(n_1523),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1593),
.A2(n_1588),
.B1(n_1594),
.B2(n_1591),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1577),
.B(n_1525),
.C(n_1523),
.Y(n_1604)
);

XNOR2xp5_ASAP7_75t_L g1605 ( 
.A(n_1579),
.B(n_1541),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1589),
.A2(n_1529),
.B1(n_1541),
.B2(n_1276),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1583),
.A2(n_1438),
.B(n_1468),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1600),
.Y(n_1608)
);

NOR3xp33_ASAP7_75t_L g1609 ( 
.A(n_1603),
.B(n_1587),
.C(n_1581),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1596),
.B(n_1578),
.Y(n_1610)
);

NOR2x1_ASAP7_75t_L g1611 ( 
.A(n_1604),
.B(n_1586),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1605),
.B(n_1580),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1599),
.B(n_1584),
.Y(n_1613)
);

NOR2x1_ASAP7_75t_L g1614 ( 
.A(n_1601),
.B(n_1586),
.Y(n_1614)
);

NAND3xp33_ASAP7_75t_L g1615 ( 
.A(n_1602),
.B(n_1597),
.C(n_1576),
.Y(n_1615)
);

NOR3x1_ASAP7_75t_L g1616 ( 
.A(n_1598),
.B(n_1590),
.C(n_1584),
.Y(n_1616)
);

NOR3xp33_ASAP7_75t_L g1617 ( 
.A(n_1607),
.B(n_1595),
.C(n_1590),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1606),
.Y(n_1618)
);

O2A1O1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1613),
.A2(n_1595),
.B(n_1217),
.C(n_1246),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1608),
.B(n_1440),
.Y(n_1620)
);

NAND3xp33_ASAP7_75t_SL g1621 ( 
.A(n_1609),
.B(n_1155),
.C(n_1188),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1612),
.B(n_1152),
.Y(n_1622)
);

NOR3xp33_ASAP7_75t_SL g1623 ( 
.A(n_1610),
.B(n_1210),
.C(n_1188),
.Y(n_1623)
);

NOR4xp75_ASAP7_75t_SL g1624 ( 
.A(n_1616),
.B(n_1209),
.C(n_1177),
.D(n_1450),
.Y(n_1624)
);

AOI211x1_ASAP7_75t_SL g1625 ( 
.A1(n_1615),
.A2(n_1447),
.B(n_1440),
.C(n_1346),
.Y(n_1625)
);

NOR2xp67_ASAP7_75t_L g1626 ( 
.A(n_1621),
.B(n_1618),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1620),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1620),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1622),
.A2(n_1611),
.B1(n_1614),
.B2(n_1617),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1619),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1625),
.B(n_1447),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1623),
.A2(n_1447),
.B1(n_1310),
.B2(n_1203),
.Y(n_1632)
);

AOI211x1_ASAP7_75t_L g1633 ( 
.A1(n_1624),
.A2(n_1398),
.B(n_1449),
.C(n_1451),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1629),
.Y(n_1634)
);

NOR2x1p5_ASAP7_75t_L g1635 ( 
.A(n_1630),
.B(n_1246),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1627),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1628),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_R g1638 ( 
.A(n_1626),
.B(n_1203),
.Y(n_1638)
);

XNOR2xp5_ASAP7_75t_L g1639 ( 
.A(n_1637),
.B(n_1634),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1636),
.Y(n_1640)
);

NOR3xp33_ASAP7_75t_L g1641 ( 
.A(n_1638),
.B(n_1632),
.C(n_1631),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1640),
.A2(n_1633),
.B1(n_1635),
.B2(n_1430),
.Y(n_1642)
);

OAI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1642),
.A2(n_1641),
.B1(n_1639),
.B2(n_1248),
.C(n_1243),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1643),
.A2(n_1248),
.B1(n_1243),
.B2(n_1187),
.Y(n_1644)
);

OAI31xp33_ASAP7_75t_L g1645 ( 
.A1(n_1643),
.A2(n_1310),
.A3(n_1418),
.B(n_1422),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1644),
.A2(n_1451),
.B(n_1449),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1645),
.A2(n_1243),
.B(n_1187),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1647),
.A2(n_1428),
.B(n_1422),
.Y(n_1648)
);

AOI221xp5_ASAP7_75t_L g1649 ( 
.A1(n_1646),
.A2(n_1430),
.B1(n_1422),
.B2(n_1428),
.C(n_1398),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_SL g1650 ( 
.A1(n_1648),
.A2(n_1248),
.B(n_1187),
.Y(n_1650)
);

AOI222xp33_ASAP7_75t_L g1651 ( 
.A1(n_1650),
.A2(n_1649),
.B1(n_1428),
.B2(n_1234),
.C1(n_1414),
.C2(n_1397),
.Y(n_1651)
);

OAI221xp5_ASAP7_75t_R g1652 ( 
.A1(n_1651),
.A2(n_1450),
.B1(n_1397),
.B2(n_1401),
.C(n_1414),
.Y(n_1652)
);

AOI211xp5_ASAP7_75t_L g1653 ( 
.A1(n_1652),
.A2(n_1179),
.B(n_1450),
.C(n_1417),
.Y(n_1653)
);


endmodule