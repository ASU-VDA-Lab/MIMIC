module fake_jpeg_18406_n_128 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_128);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_16),
.Y(n_36)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_23),
.Y(n_49)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_50),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_25),
.C(n_24),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_44),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_14),
.B1(n_18),
.B2(n_21),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR4xp25_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_11),
.C(n_10),
.D(n_4),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_52),
.Y(n_68)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_44),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_18),
.B1(n_19),
.B2(n_15),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_62),
.B1(n_71),
.B2(n_65),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_15),
.B1(n_19),
.B2(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_1),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_1),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_16),
.B(n_13),
.C(n_2),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_4),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_6),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_6),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_74),
.B1(n_70),
.B2(n_66),
.Y(n_86)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_84),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_89),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_77),
.A2(n_55),
.B(n_48),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_87),
.B(n_71),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g84 ( 
.A(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_76),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_55),
.B(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_48),
.B1(n_58),
.B2(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_58),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_87),
.B(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_96),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_77),
.B(n_65),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_62),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_86),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_95),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_92),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_110),
.B1(n_82),
.B2(n_91),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_112),
.Y(n_119)
);

OAI321xp33_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_97),
.A3(n_93),
.B1(n_64),
.B2(n_52),
.C(n_43),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_115),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_72),
.B(n_13),
.C(n_46),
.D(n_59),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_90),
.C(n_72),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_105),
.C(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_120),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_103),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_119),
.C(n_90),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_115),
.B1(n_103),
.B2(n_112),
.Y(n_123)
);

AOI31xp67_ASAP7_75t_SL g125 ( 
.A1(n_123),
.A2(n_46),
.A3(n_8),
.B(n_11),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_124),
.B(n_125),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_121),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_7),
.Y(n_128)
);


endmodule