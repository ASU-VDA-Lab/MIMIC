module fake_jpeg_25360_n_249 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_0),
.C(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_52),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_19),
.B1(n_20),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_32),
.Y(n_52)
);

CKINVDCx9p33_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_25),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_40),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_75),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_67),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_66),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_41),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_38),
.B1(n_19),
.B2(n_39),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_69),
.A2(n_87),
.B1(n_57),
.B2(n_28),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_73),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_34),
.B(n_26),
.C(n_30),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_17),
.Y(n_94)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_27),
.B1(n_32),
.B2(n_30),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_79),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_27),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_47),
.B(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_86),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_42),
.B1(n_35),
.B2(n_16),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_44),
.B1(n_35),
.B2(n_42),
.Y(n_102)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_45),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_33),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_43),
.A2(n_17),
.B1(n_33),
.B2(n_22),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_94),
.B(n_68),
.Y(n_129)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_73),
.B1(n_85),
.B2(n_64),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_45),
.B(n_1),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_112),
.B(n_115),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_33),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_86),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_35),
.B1(n_42),
.B2(n_49),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_89),
.B1(n_68),
.B2(n_77),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_22),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_13),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_110),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_29),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_35),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_28),
.A3(n_25),
.B1(n_24),
.B2(n_21),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_117),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_140),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_124),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_84),
.B1(n_82),
.B2(n_63),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_121),
.B1(n_138),
.B2(n_139),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_60),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_70),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_133),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_93),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_113),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_101),
.A2(n_88),
.B(n_78),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_136),
.B(n_92),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_98),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_137),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_61),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_132),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_83),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_94),
.B(n_29),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_96),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_97),
.A2(n_80),
.B(n_74),
.Y(n_136)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_74),
.B1(n_64),
.B2(n_25),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_97),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_112),
.C(n_111),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_148),
.C(n_162),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_158),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_100),
.C(n_103),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_146),
.B(n_152),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_165),
.B(n_131),
.Y(n_180)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_156),
.Y(n_178)
);

NOR4xp25_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_123),
.C(n_130),
.D(n_122),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_112),
.C(n_111),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_111),
.C(n_105),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_166),
.C(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_164),
.B(n_28),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_114),
.B(n_115),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_102),
.C(n_99),
.Y(n_166)
);

NAND4xp25_ASAP7_75t_SL g170 ( 
.A(n_144),
.B(n_116),
.C(n_57),
.D(n_137),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_170),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_181),
.Y(n_192)
);

XOR2x2_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_129),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_163),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_134),
.C(n_127),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_175),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_160),
.A2(n_127),
.B1(n_121),
.B2(n_139),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_174),
.A2(n_179),
.B1(n_180),
.B2(n_187),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_123),
.C(n_124),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_117),
.C(n_24),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_183),
.Y(n_190)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_21),
.C(n_16),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_166),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_0),
.B(n_1),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_185),
.A2(n_158),
.B1(n_154),
.B2(n_3),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_151),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_24),
.B1(n_21),
.B2(n_16),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_178),
.B(n_142),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_194),
.Y(n_215)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_168),
.B(n_181),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_200),
.B(n_180),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_185),
.B1(n_176),
.B2(n_172),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_202),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_161),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_169),
.A2(n_165),
.B1(n_149),
.B2(n_164),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_174),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_164),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_0),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_2),
.Y(n_209)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_207),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_167),
.C(n_173),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_208),
.A2(n_210),
.B(n_186),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_213),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_170),
.B(n_5),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_188),
.C(n_202),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_169),
.B1(n_167),
.B2(n_184),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_200),
.B1(n_197),
.B2(n_195),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_188),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_223),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_230)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_199),
.B(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_205),
.B(n_204),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_222),
.B(n_12),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_3),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_225),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_213),
.B(n_3),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_207),
.B(n_212),
.Y(n_227)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_212),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_230),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_5),
.B(n_6),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_233),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_217),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_238),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_218),
.C(n_7),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_10),
.C(n_6),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_12),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_231),
.C(n_7),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_239),
.A2(n_9),
.B1(n_10),
.B2(n_234),
.Y(n_242)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_238),
.B(n_9),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_10),
.B(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_245),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_247),
.Y(n_249)
);


endmodule