module fake_aes_1559_n_554 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_554);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_554;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_67;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_70;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_64;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_63;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g62 ( .A(n_48), .Y(n_62) );
INVx1_ASAP7_75t_L g63 ( .A(n_53), .Y(n_63) );
INVx1_ASAP7_75t_L g64 ( .A(n_56), .Y(n_64) );
INVxp67_ASAP7_75t_SL g65 ( .A(n_50), .Y(n_65) );
INVxp33_ASAP7_75t_SL g66 ( .A(n_18), .Y(n_66) );
INVxp67_ASAP7_75t_SL g67 ( .A(n_26), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_21), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_39), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_11), .Y(n_70) );
CKINVDCx16_ASAP7_75t_R g71 ( .A(n_19), .Y(n_71) );
CKINVDCx16_ASAP7_75t_R g72 ( .A(n_34), .Y(n_72) );
HB1xp67_ASAP7_75t_L g73 ( .A(n_57), .Y(n_73) );
INVx1_ASAP7_75t_SL g74 ( .A(n_47), .Y(n_74) );
BUFx2_ASAP7_75t_L g75 ( .A(n_36), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_13), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_49), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_3), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_40), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_25), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_45), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_42), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_30), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_55), .Y(n_84) );
INVxp33_ASAP7_75t_SL g85 ( .A(n_5), .Y(n_85) );
INVx1_ASAP7_75t_SL g86 ( .A(n_60), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_22), .Y(n_87) );
INVxp33_ASAP7_75t_SL g88 ( .A(n_29), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_61), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_15), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_2), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_16), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_0), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_38), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_10), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_8), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_28), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_10), .Y(n_98) );
HB1xp67_ASAP7_75t_L g99 ( .A(n_51), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_23), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_52), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_37), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_4), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_14), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_33), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_43), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_3), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_73), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_89), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_89), .Y(n_110) );
NOR2xp33_ASAP7_75t_R g111 ( .A(n_71), .B(n_32), .Y(n_111) );
NOR2xp33_ASAP7_75t_R g112 ( .A(n_71), .B(n_31), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_99), .Y(n_113) );
AND2x4_ASAP7_75t_L g114 ( .A(n_75), .B(n_0), .Y(n_114) );
NAND2xp33_ASAP7_75t_SL g115 ( .A(n_75), .B(n_1), .Y(n_115) );
AND2x6_ASAP7_75t_L g116 ( .A(n_89), .B(n_35), .Y(n_116) );
BUFx8_ASAP7_75t_L g117 ( .A(n_62), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_101), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_72), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_72), .B(n_1), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_79), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_79), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_95), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_70), .Y(n_124) );
BUFx3_ASAP7_75t_L g125 ( .A(n_62), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_101), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_63), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_95), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_105), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_107), .Y(n_130) );
BUFx10_ASAP7_75t_L g131 ( .A(n_84), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_63), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_64), .B(n_2), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_107), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_64), .Y(n_135) );
BUFx10_ASAP7_75t_L g136 ( .A(n_94), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_68), .B(n_4), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_68), .B(n_5), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_105), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_70), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_66), .Y(n_141) );
NOR2xp33_ASAP7_75t_R g142 ( .A(n_69), .B(n_44), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_88), .Y(n_143) );
INVxp67_ASAP7_75t_L g144 ( .A(n_76), .Y(n_144) );
XOR2xp5_ASAP7_75t_L g145 ( .A(n_85), .B(n_6), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_76), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_69), .B(n_6), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_78), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_110), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_109), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_109), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_108), .B(n_102), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_109), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_110), .Y(n_155) );
AO22x2_ASAP7_75t_L g156 ( .A1(n_114), .A2(n_106), .B1(n_77), .B2(n_80), .Y(n_156) );
INVx1_ASAP7_75t_SL g157 ( .A(n_119), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_116), .Y(n_158) );
OR2x2_ASAP7_75t_L g159 ( .A(n_124), .B(n_144), .Y(n_159) );
INVxp67_ASAP7_75t_SL g160 ( .A(n_125), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_113), .B(n_106), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_109), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_118), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_116), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_114), .B(n_90), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_125), .B(n_87), .Y(n_166) );
INVxp33_ASAP7_75t_L g167 ( .A(n_120), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_121), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_118), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_114), .B(n_93), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_118), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_146), .B(n_90), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_131), .B(n_80), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_111), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_146), .B(n_91), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_126), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_126), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_126), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_126), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_127), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_127), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_131), .B(n_87), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_130), .B(n_134), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_132), .Y(n_184) );
INVxp67_ASAP7_75t_SL g185 ( .A(n_117), .Y(n_185) );
INVx1_ASAP7_75t_SL g186 ( .A(n_129), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_131), .B(n_82), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_136), .Y(n_189) );
AO22x2_ASAP7_75t_L g190 ( .A1(n_145), .A2(n_82), .B1(n_97), .B2(n_77), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_135), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_135), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_116), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_136), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_116), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_140), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_139), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_123), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_128), .Y(n_199) );
NAND3x1_ASAP7_75t_L g200 ( .A(n_133), .B(n_96), .C(n_103), .Y(n_200) );
AO22x2_ASAP7_75t_L g201 ( .A1(n_137), .A2(n_97), .B1(n_103), .B2(n_78), .Y(n_201) );
NAND3xp33_ASAP7_75t_L g202 ( .A(n_138), .B(n_91), .C(n_92), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_148), .B(n_92), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_147), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_136), .B(n_98), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_142), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_159), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_192), .Y(n_208) );
OR2x2_ASAP7_75t_L g209 ( .A(n_159), .B(n_115), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_157), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_168), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_204), .B(n_93), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_204), .B(n_117), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_172), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_180), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_156), .A2(n_143), .B1(n_141), .B2(n_122), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_168), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_156), .Y(n_218) );
NOR2xp33_ASAP7_75t_R g219 ( .A(n_197), .B(n_115), .Y(n_219) );
OR2x6_ASAP7_75t_L g220 ( .A(n_156), .B(n_98), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g221 ( .A(n_164), .B(n_96), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_180), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_170), .B(n_104), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_184), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_184), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_192), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_198), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_191), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_191), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_183), .B(n_112), .Y(n_230) );
OR2x2_ASAP7_75t_L g231 ( .A(n_186), .B(n_7), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_172), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_176), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_196), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_156), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_177), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_170), .B(n_65), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_201), .A2(n_112), .B1(n_111), .B2(n_142), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_153), .B(n_86), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_149), .Y(n_240) );
NOR2xp33_ASAP7_75t_R g241 ( .A(n_197), .B(n_46), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_179), .Y(n_242) );
INVx5_ASAP7_75t_L g243 ( .A(n_193), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_149), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_179), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_206), .B(n_74), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_155), .Y(n_247) );
BUFx2_ASAP7_75t_L g248 ( .A(n_201), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_185), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_160), .B(n_100), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_155), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_175), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_206), .B(n_83), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_196), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_193), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_183), .B(n_67), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_193), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_196), .B(n_81), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_201), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_196), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_201), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_181), .Y(n_262) );
INVx5_ASAP7_75t_L g263 ( .A(n_220), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_220), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_232), .Y(n_265) );
OR2x6_ASAP7_75t_L g266 ( .A(n_220), .B(n_170), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_252), .Y(n_267) );
AND2x2_ASAP7_75t_SL g268 ( .A(n_218), .B(n_235), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_210), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_214), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_214), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_212), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_254), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_212), .B(n_170), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_212), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_230), .B(n_165), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_230), .B(n_165), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_254), .A2(n_164), .B(n_158), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_255), .Y(n_279) );
OAI22xp5_ASAP7_75t_SL g280 ( .A1(n_211), .A2(n_167), .B1(n_190), .B2(n_174), .Y(n_280) );
INVxp67_ASAP7_75t_L g281 ( .A(n_207), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_260), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_234), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_255), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_240), .Y(n_285) );
NAND3xp33_ASAP7_75t_L g286 ( .A(n_238), .B(n_202), .C(n_205), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_234), .Y(n_287) );
O2A1O1Ixp33_ASAP7_75t_L g288 ( .A1(n_261), .A2(n_161), .B(n_166), .C(n_202), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_208), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_207), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_213), .A2(n_164), .B(n_152), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_223), .B(n_175), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_218), .Y(n_293) );
INVx5_ASAP7_75t_L g294 ( .A(n_243), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_209), .B(n_173), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_221), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_221), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_209), .A2(n_190), .B1(n_182), .B2(n_187), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_256), .B(n_203), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_255), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_208), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_256), .B(n_203), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_223), .B(n_194), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_249), .Y(n_304) );
NAND2x1_ASAP7_75t_L g305 ( .A(n_240), .B(n_188), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_248), .B(n_190), .Y(n_306) );
INVx2_ASAP7_75t_SL g307 ( .A(n_221), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_248), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_289), .Y(n_309) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_286), .A2(n_259), .B(n_229), .C(n_228), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_265), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_263), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_290), .B(n_223), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_269), .A2(n_211), .B1(n_217), .B2(n_216), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_278), .A2(n_255), .B(n_257), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_266), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_269), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_281), .B(n_304), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_266), .B(n_259), .Y(n_319) );
BUFx12f_ASAP7_75t_L g320 ( .A(n_266), .Y(n_320) );
NAND2x1_ASAP7_75t_L g321 ( .A(n_266), .B(n_244), .Y(n_321) );
O2A1O1Ixp33_ASAP7_75t_L g322 ( .A1(n_276), .A2(n_231), .B(n_258), .C(n_246), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_263), .A2(n_237), .B1(n_244), .B2(n_247), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_263), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_299), .B(n_302), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_280), .Y(n_326) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_263), .B(n_247), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_263), .A2(n_237), .B1(n_251), .B2(n_215), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_274), .A2(n_237), .B1(n_251), .B2(n_215), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_306), .A2(n_222), .B1(n_225), .B2(n_228), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_267), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_306), .A2(n_219), .B1(n_231), .B2(n_239), .Y(n_332) );
NAND3xp33_ASAP7_75t_SL g333 ( .A(n_298), .B(n_241), .C(n_224), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_295), .B(n_189), .Y(n_334) );
NAND3xp33_ASAP7_75t_SL g335 ( .A(n_288), .B(n_229), .C(n_225), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_319), .B(n_316), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_311), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_327), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_331), .Y(n_339) );
AO21x2_ASAP7_75t_L g340 ( .A1(n_335), .A2(n_285), .B(n_291), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_325), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_326), .A2(n_268), .B1(n_272), .B2(n_275), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_318), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_313), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_315), .A2(n_305), .B(n_273), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_334), .B(n_277), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_309), .Y(n_347) );
INVxp67_ASAP7_75t_L g348 ( .A(n_317), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_330), .A2(n_308), .B1(n_271), .B2(n_270), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_335), .A2(n_273), .B(n_282), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_322), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_314), .A2(n_274), .B1(n_302), .B2(n_299), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_330), .A2(n_293), .B1(n_274), .B2(n_198), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_332), .B(n_198), .C(n_303), .Y(n_354) );
AO21x2_ASAP7_75t_L g355 ( .A1(n_333), .A2(n_224), .B(n_222), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_319), .A2(n_264), .B1(n_307), .B2(n_297), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_329), .A2(n_297), .B1(n_296), .B2(n_292), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_310), .A2(n_300), .B(n_279), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_327), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_343), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_337), .Y(n_361) );
OR2x6_ASAP7_75t_L g362 ( .A(n_338), .B(n_320), .Y(n_362) );
OAI211xp5_ASAP7_75t_SL g363 ( .A1(n_348), .A2(n_194), .B(n_316), .C(n_253), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_352), .B(n_333), .Y(n_364) );
NAND2x1p5_ASAP7_75t_SL g365 ( .A(n_338), .B(n_289), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_359), .B(n_312), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_341), .B(n_321), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_342), .A2(n_328), .B1(n_323), .B2(n_198), .Y(n_368) );
INVxp67_ASAP7_75t_SL g369 ( .A(n_359), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_350), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_350), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g372 ( .A1(n_346), .A2(n_250), .B1(n_297), .B2(n_296), .C(n_199), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_347), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_344), .B(n_199), .Y(n_374) );
NAND3xp33_ASAP7_75t_L g375 ( .A(n_351), .B(n_198), .C(n_171), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_336), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_345), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_339), .Y(n_378) );
OR2x6_ASAP7_75t_L g379 ( .A(n_357), .B(n_312), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_345), .Y(n_381) );
BUFx3_ASAP7_75t_L g382 ( .A(n_336), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
NAND2xp33_ASAP7_75t_R g384 ( .A(n_358), .B(n_296), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_349), .B(n_301), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_354), .A2(n_282), .B1(n_312), .B2(n_324), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_353), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_355), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_364), .A2(n_356), .B1(n_200), .B2(n_355), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_377), .Y(n_390) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_369), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_373), .Y(n_392) );
CKINVDCx16_ASAP7_75t_R g393 ( .A(n_362), .Y(n_393) );
INVx4_ASAP7_75t_L g394 ( .A(n_379), .Y(n_394) );
OAI31xp33_ASAP7_75t_SL g395 ( .A1(n_364), .A2(n_7), .A3(n_8), .B(n_9), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_361), .B(n_340), .Y(n_396) );
OAI33xp33_ASAP7_75t_L g397 ( .A1(n_360), .A2(n_178), .A3(n_163), .B1(n_169), .B2(n_262), .B3(n_150), .Y(n_397) );
OAI31xp33_ASAP7_75t_L g398 ( .A1(n_372), .A2(n_181), .A3(n_188), .B(n_283), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_378), .B(n_340), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_387), .B(n_324), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_376), .B(n_324), .Y(n_401) );
INVxp67_ASAP7_75t_SL g402 ( .A(n_385), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_388), .Y(n_403) );
NOR2x1_ASAP7_75t_SL g404 ( .A(n_379), .B(n_294), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_376), .B(n_54), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_377), .Y(n_406) );
NAND4xp25_ASAP7_75t_L g407 ( .A(n_383), .B(n_163), .C(n_169), .D(n_150), .Y(n_407) );
BUFx3_ASAP7_75t_L g408 ( .A(n_366), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_368), .A2(n_287), .B1(n_283), .B2(n_193), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_367), .Y(n_410) );
OAI21xp5_ASAP7_75t_SL g411 ( .A1(n_368), .A2(n_287), .B(n_283), .Y(n_411) );
OAI33xp33_ASAP7_75t_L g412 ( .A1(n_374), .A2(n_163), .A3(n_169), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_381), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_362), .B(n_12), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_370), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_376), .B(n_12), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_366), .B(n_13), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_370), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_371), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_371), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_362), .B(n_17), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_365), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_380), .B(n_17), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_380), .B(n_226), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_382), .B(n_226), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_365), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_382), .A2(n_287), .B1(n_158), .B2(n_195), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_388), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_388), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_414), .B(n_363), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_421), .B(n_379), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_410), .B(n_386), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_426), .B(n_386), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_394), .B(n_388), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_392), .B(n_375), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_405), .B(n_294), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_393), .B(n_20), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_391), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_417), .B(n_24), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_396), .B(n_171), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_396), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_399), .B(n_171), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_415), .Y(n_443) );
OAI221xp5_ASAP7_75t_L g444 ( .A1(n_395), .A2(n_384), .B1(n_171), .B2(n_151), .C(n_162), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_415), .Y(n_445) );
NAND2xp33_ASAP7_75t_R g446 ( .A(n_426), .B(n_27), .Y(n_446) );
INVxp67_ASAP7_75t_L g447 ( .A(n_423), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_415), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_393), .B(n_41), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_418), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_418), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_416), .Y(n_452) );
AND2x2_ASAP7_75t_SL g453 ( .A(n_394), .B(n_300), .Y(n_453) );
OAI31xp33_ASAP7_75t_L g454 ( .A1(n_398), .A2(n_227), .A3(n_152), .B(n_195), .Y(n_454) );
NOR2xp33_ASAP7_75t_R g455 ( .A(n_394), .B(n_58), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_408), .B(n_59), .Y(n_456) );
AOI21xp33_ASAP7_75t_L g457 ( .A1(n_422), .A2(n_171), .B(n_154), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_408), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_389), .B(n_294), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_424), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_412), .B(n_227), .C(n_245), .Y(n_462) );
AND2x2_ASAP7_75t_SL g463 ( .A(n_405), .B(n_300), .Y(n_463) );
INVx5_ASAP7_75t_L g464 ( .A(n_405), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_402), .B(n_151), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_400), .B(n_151), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_400), .B(n_151), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_401), .B(n_154), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g469 ( .A1(n_430), .A2(n_397), .B1(n_405), .B2(n_404), .C1(n_419), .C2(n_411), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_441), .B(n_389), .Y(n_470) );
NOR3xp33_ASAP7_75t_SL g471 ( .A(n_446), .B(n_398), .C(n_407), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_438), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g473 ( .A(n_464), .B(n_401), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_430), .A2(n_407), .B1(n_401), .B2(n_425), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_464), .A2(n_409), .B1(n_401), .B2(n_406), .Y(n_475) );
OAI31xp33_ASAP7_75t_L g476 ( .A1(n_444), .A2(n_429), .A3(n_403), .B(n_428), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_452), .Y(n_477) );
INVxp67_ASAP7_75t_L g478 ( .A(n_446), .Y(n_478) );
OAI32xp33_ASAP7_75t_L g479 ( .A1(n_436), .A2(n_413), .A3(n_428), .B1(n_390), .B2(n_404), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_432), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_447), .B(n_437), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_431), .A2(n_420), .B1(n_390), .B2(n_427), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_431), .A2(n_420), .B1(n_390), .B2(n_162), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_461), .Y(n_484) );
OAI322xp33_ASAP7_75t_L g485 ( .A1(n_459), .A2(n_154), .A3(n_162), .B1(n_227), .B2(n_245), .C1(n_242), .C2(n_233), .Y(n_485) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_465), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_458), .B(n_154), .Y(n_487) );
INVxp67_ASAP7_75t_L g488 ( .A(n_437), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_435), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_443), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_443), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_449), .B(n_284), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_445), .B(n_236), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_453), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_453), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_449), .A2(n_454), .B(n_463), .C(n_439), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_448), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_472), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_489), .B(n_450), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_484), .Y(n_500) );
OAI22xp33_ASAP7_75t_L g501 ( .A1(n_478), .A2(n_436), .B1(n_433), .B2(n_455), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_488), .B(n_433), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_477), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_480), .B(n_450), .Y(n_504) );
NOR3xp33_ASAP7_75t_SL g505 ( .A(n_496), .B(n_442), .C(n_440), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_486), .B(n_448), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_473), .Y(n_507) );
NAND3xp33_ASAP7_75t_L g508 ( .A(n_469), .B(n_468), .C(n_462), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_470), .B(n_460), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_481), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_490), .Y(n_511) );
NAND2xp33_ASAP7_75t_SL g512 ( .A(n_471), .B(n_456), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_491), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_497), .Y(n_514) );
NOR2xp33_ASAP7_75t_R g515 ( .A(n_494), .B(n_466), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_495), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_487), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_482), .B(n_434), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_474), .B(n_460), .Y(n_519) );
NOR2xp33_ASAP7_75t_R g520 ( .A(n_492), .B(n_467), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_493), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_483), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_512), .A2(n_502), .B1(n_508), .B2(n_505), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_500), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_499), .B(n_451), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_501), .A2(n_476), .B(n_479), .Y(n_526) );
NOR2x1p5_ASAP7_75t_L g527 ( .A(n_507), .B(n_469), .Y(n_527) );
NOR2x1_ASAP7_75t_L g528 ( .A(n_501), .B(n_485), .Y(n_528) );
BUFx2_ASAP7_75t_L g529 ( .A(n_515), .Y(n_529) );
NOR2xp67_ASAP7_75t_L g530 ( .A(n_507), .B(n_475), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_505), .A2(n_519), .B1(n_518), .B2(n_522), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_515), .Y(n_532) );
AOI322xp5_ASAP7_75t_L g533 ( .A1(n_523), .A2(n_510), .A3(n_503), .B1(n_516), .B2(n_498), .C1(n_506), .C2(n_509), .Y(n_533) );
AOI21xp33_ASAP7_75t_L g534 ( .A1(n_528), .A2(n_517), .B(n_521), .Y(n_534) );
AO22x2_ASAP7_75t_L g535 ( .A1(n_532), .A2(n_513), .B1(n_511), .B2(n_514), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_527), .A2(n_531), .B1(n_532), .B2(n_529), .Y(n_536) );
XNOR2x1_ASAP7_75t_L g537 ( .A(n_524), .B(n_517), .Y(n_537) );
NOR3xp33_ASAP7_75t_L g538 ( .A(n_526), .B(n_504), .C(n_457), .Y(n_538) );
NOR2xp67_ASAP7_75t_L g539 ( .A(n_530), .B(n_520), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_525), .A2(n_523), .B1(n_527), .B2(n_512), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_529), .A2(n_512), .B(n_526), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_524), .Y(n_542) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_542), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_537), .Y(n_544) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_539), .B(n_541), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_535), .Y(n_546) );
XNOR2x1_ASAP7_75t_L g547 ( .A(n_544), .B(n_536), .Y(n_547) );
NAND3xp33_ASAP7_75t_SL g548 ( .A(n_545), .B(n_540), .C(n_533), .Y(n_548) );
BUFx3_ASAP7_75t_L g549 ( .A(n_545), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_549), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_548), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_550), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_552), .A2(n_551), .B1(n_547), .B2(n_543), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_553), .A2(n_546), .B1(n_538), .B2(n_534), .Y(n_554) );
endmodule