module fake_netlist_1_9412_n_42 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_42);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
CKINVDCx16_ASAP7_75t_R g17 ( .A(n_11), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_12), .B(n_9), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_7), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_10), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_13), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_8), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_14), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_16), .B(n_0), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
NOR2xp67_ASAP7_75t_L g26 ( .A(n_19), .B(n_0), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_21), .B(n_1), .Y(n_27) );
BUFx6f_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
OA21x2_ASAP7_75t_L g29 ( .A1(n_24), .A2(n_20), .B(n_21), .Y(n_29) );
AOI22xp33_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_25), .B1(n_26), .B2(n_20), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
NAND2x1p5_ASAP7_75t_L g32 ( .A(n_31), .B(n_28), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_28), .Y(n_33) );
OAI22xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_28), .B1(n_17), .B2(n_29), .Y(n_34) );
AOI22xp33_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_28), .B1(n_29), .B2(n_23), .Y(n_35) );
O2A1O1Ixp33_ASAP7_75t_SL g36 ( .A1(n_35), .A2(n_18), .B(n_15), .C(n_22), .Y(n_36) );
NOR4xp25_ASAP7_75t_L g37 ( .A(n_34), .B(n_1), .C(n_2), .D(n_3), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_37), .B(n_2), .Y(n_38) );
A2O1A1Ixp33_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_22), .B(n_4), .C(n_5), .Y(n_39) );
NAND2xp5_ASAP7_75t_R g40 ( .A(n_38), .B(n_6), .Y(n_40) );
AOI22x1_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_7), .B1(n_38), .B2(n_39), .Y(n_41) );
BUFx2_ASAP7_75t_SL g42 ( .A(n_41), .Y(n_42) );
endmodule