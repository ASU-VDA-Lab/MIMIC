module fake_jpeg_17892_n_31 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_31;

wire n_13;
wire n_21;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_15;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_8),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_3),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_2),
.Y(n_15)
);

INVx4_ASAP7_75t_SL g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_0),
.B1(n_6),
.B2(n_9),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_5),
.A2(n_3),
.B(n_4),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_0),
.C(n_7),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.C(n_23),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_12),
.C(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_16),
.A2(n_18),
.B1(n_17),
.B2(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_11),
.A2(n_15),
.B1(n_12),
.B2(n_18),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_16),
.B1(n_22),
.B2(n_20),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_15),
.Y(n_30)
);

AOI332xp33_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_13),
.A3(n_14),
.B1(n_21),
.B2(n_26),
.B3(n_28),
.C1(n_29),
.C2(n_25),
.Y(n_31)
);


endmodule