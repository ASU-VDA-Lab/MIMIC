module real_jpeg_6014_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_1),
.Y(n_107)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_1),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_2),
.A2(n_66),
.B1(n_80),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_2),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_2),
.A2(n_149),
.B1(n_237),
.B2(n_256),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_2),
.A2(n_237),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_2),
.A2(n_185),
.B1(n_237),
.B2(n_380),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_3),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_4),
.A2(n_79),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_4),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_4),
.A2(n_86),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_4),
.A2(n_86),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_4),
.A2(n_86),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_5),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_5),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_5),
.A2(n_81),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_5),
.A2(n_81),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_5),
.A2(n_81),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_7),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_7),
.Y(n_190)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_7),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_7),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g395 ( 
.A(n_7),
.Y(n_395)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_8),
.Y(n_272)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_10),
.Y(n_442)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_11),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_12),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_12),
.A2(n_51),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_12),
.A2(n_51),
.B1(n_192),
.B2(n_195),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_12),
.B(n_68),
.Y(n_285)
);

O2A1O1Ixp33_ASAP7_75t_L g340 ( 
.A1(n_12),
.A2(n_23),
.B(n_341),
.C(n_348),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_12),
.B(n_370),
.C(n_371),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_12),
.B(n_21),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_12),
.B(n_290),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_12),
.B(n_101),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_13),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_13),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_440),
.B(n_443),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_155),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_153),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_18),
.B(n_133),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_55),
.B1(n_56),
.B2(n_87),
.Y(n_19)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_20),
.A2(n_87),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_34),
.B(n_48),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_21),
.B(n_123),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_21),
.A2(n_121),
.B(n_147),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_21),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_22),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx5_ASAP7_75t_L g356 ( 
.A(n_25),
.Y(n_356)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_27),
.Y(n_178)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_27),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_27),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_29),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_29),
.Y(n_199)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_29),
.Y(n_347)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_34),
.A2(n_147),
.B(n_151),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_34),
.B(n_48),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_34),
.B(n_255),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_35),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_38),
.Y(n_344)
);

AOI32xp33_ASAP7_75t_L g261 ( 
.A1(n_39),
.A2(n_262),
.A3(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_261)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_41),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_45),
.Y(n_148)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_47),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_47),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_48),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_51),
.A2(n_60),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_51),
.B(n_144),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g341 ( 
.A1(n_51),
.A2(n_342),
.B(n_345),
.Y(n_341)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_78),
.B(n_82),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_57),
.A2(n_131),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_58),
.B(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_58),
.B(n_236),
.Y(n_235)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_68),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_63),
.Y(n_262)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_68),
.B(n_142),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_68),
.B(n_236),
.Y(n_250)
);

AO22x2_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_75),
.Y(n_269)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_78),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_82),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_82),
.B(n_235),
.Y(n_302)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_87),
.B(n_311),
.C(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_118),
.C(n_129),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_118),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_89),
.A2(n_139),
.B1(n_146),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_89),
.A2(n_139),
.B1(n_252),
.B2(n_258),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_89),
.B(n_249),
.C(n_252),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_112),
.B(n_113),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_90),
.A2(n_197),
.B(n_204),
.Y(n_196)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_91),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_91),
.B(n_114),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_91),
.B(n_355),
.Y(n_354)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_101),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_97),
.B2(n_100),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AO22x2_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_102),
.B1(n_104),
.B2(n_108),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_101),
.B(n_173),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_101),
.B(n_355),
.Y(n_374)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_107),
.Y(n_227)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_110),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_111),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_112),
.B(n_113),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_112),
.A2(n_172),
.B(n_197),
.Y(n_230)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_119),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_121),
.Y(n_253)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_124),
.Y(n_257)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_130),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_132),
.B(n_250),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_140),
.C(n_145),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_134),
.A2(n_135),
.B1(n_140),
.B2(n_163),
.Y(n_240)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_140),
.C(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_141),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_143),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_145),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_152),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_152),
.B(n_283),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_242),
.B(n_436),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_238),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_208),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_159),
.B(n_208),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_180),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_167),
.B2(n_168),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_162),
.B(n_167),
.C(n_180),
.Y(n_241)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_168),
.A2(n_169),
.B(n_179),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_179),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_170),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_172),
.B(n_374),
.Y(n_416)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_205),
.B(n_206),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_182),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_196),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_205),
.B1(n_206),
.B2(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_183),
.A2(n_196),
.B1(n_205),
.B2(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_183),
.B(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_183),
.A2(n_205),
.B1(n_340),
.B2(n_419),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_189),
.B(n_191),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_184),
.B(n_191),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_184),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_184),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_186),
.Y(n_381)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_194),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_196),
.Y(n_323)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_204),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_204),
.B(n_354),
.Y(n_383)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.C(n_215),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_209),
.A2(n_213),
.B1(n_214),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_209),
.Y(n_327)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_215),
.B(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_231),
.C(n_233),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_216),
.A2(n_217),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_230),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_218),
.B(n_230),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_219),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_223),
.B(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_224),
.A2(n_274),
.B(n_279),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_225),
.B(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_227),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_231),
.B(n_233),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_232),
.B(n_254),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_238),
.A2(n_438),
.B(n_439),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_239),
.B(n_241),
.Y(n_439)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_428),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_316),
.C(n_330),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_305),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_291),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_247),
.B(n_291),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_259),
.C(n_281),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_248),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_259),
.A2(n_260),
.B1(n_281),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_273),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_261),
.B(n_273),
.Y(n_300)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp33_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_274),
.A2(n_288),
.B(n_296),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_281),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.C(n_286),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_287),
.B(n_393),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_288),
.B(n_378),
.Y(n_406)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_299),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_294),
.C(n_299),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_297),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_298),
.B(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_302),
.C(n_303),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_305),
.A2(n_431),
.B(n_432),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_315),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_306),
.B(n_315),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_309),
.C(n_310),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_328),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_317),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_325),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_318),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_318),
.B(n_329),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_318),
.B(n_325),
.Y(n_435)
);

FAx1_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_322),
.CI(n_324),
.CON(n_318),
.SN(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_328),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_360),
.B(n_427),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_332),
.B(n_335),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.C(n_351),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_336),
.B(n_423),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_339),
.A2(n_351),
.B1(n_352),
.B2(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_339),
.Y(n_424)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx8_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_SL g345 ( 
.A(n_346),
.Y(n_345)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx12f_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_421),
.B(n_426),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_411),
.B(n_420),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_387),
.B(n_410),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_375),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_375),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_373),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_365),
.A2(n_366),
.B1(n_373),
.B2(n_390),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_373),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_382),
.Y(n_375)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_376),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_383),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_382)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_383),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_384),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_385),
.C(n_413),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_396),
.B(n_409),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_391),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_391),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_405),
.B(n_408),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_404),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_403),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_406),
.B(n_407),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_414),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_418),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_417),
.C(n_418),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_425),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_425),
.Y(n_426)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g428 ( 
.A1(n_429),
.A2(n_430),
.B(n_433),
.C(n_434),
.D(n_435),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx5_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx8_ASAP7_75t_L g444 ( 
.A(n_442),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);


endmodule