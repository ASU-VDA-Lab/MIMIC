module real_jpeg_26743_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_335, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_335;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_0),
.B(n_49),
.Y(n_91)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_0),
.Y(n_249)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_2),
.A2(n_27),
.B1(n_49),
.B2(n_51),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_2),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_4),
.A2(n_44),
.B1(n_55),
.B2(n_56),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_4),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_44),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_5),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_117),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_117),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_5),
.A2(n_49),
.B1(n_51),
.B2(n_117),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_6),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_6),
.A2(n_29),
.B(n_33),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_121),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_6),
.B(n_31),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_6),
.A2(n_55),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_6),
.B(n_55),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_6),
.B(n_71),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_6),
.A2(n_90),
.B1(n_245),
.B2(n_249),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_6),
.A2(n_32),
.B(n_261),
.Y(n_260)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_8),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_111),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_111),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_8),
.A2(n_49),
.B1(n_51),
.B2(n_111),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_9),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_9),
.A2(n_46),
.B1(n_55),
.B2(n_56),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_46),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_10),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_106),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_106),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_10),
.A2(n_49),
.B1(n_51),
.B2(n_106),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_48)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_12),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_108),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_12),
.A2(n_49),
.B1(n_51),
.B2(n_108),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_108),
.Y(n_265)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_15),
.A2(n_37),
.B1(n_55),
.B2(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_15),
.A2(n_37),
.B1(n_49),
.B2(n_51),
.Y(n_130)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_16),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_17),
.A2(n_55),
.B1(n_56),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_17),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_101),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_101),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_17),
.A2(n_49),
.B1(n_51),
.B2(n_101),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_79),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_38),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_23),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_25),
.A2(n_35),
.B(n_121),
.C(n_122),
.Y(n_120)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_31),
.B1(n_42),
.B2(n_45),
.Y(n_41)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_28),
.A2(n_31),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_28),
.A2(n_31),
.B1(n_107),
.B2(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_28),
.A2(n_31),
.B1(n_116),
.B2(n_188),
.Y(n_187)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_31),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_63),
.B(n_65),
.C(n_66),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_63),
.Y(n_65)
);

OAI32xp33_ASAP7_75t_L g269 ( 
.A1(n_32),
.A2(n_56),
.A3(n_67),
.B1(n_262),
.B2(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_33),
.B(n_121),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_72),
.C(n_74),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_39),
.A2(n_40),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.C(n_60),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_41),
.B(n_318),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_43),
.A2(n_76),
.B1(n_78),
.B2(n_168),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_47),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_47),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_47),
.A2(n_60),
.B1(n_312),
.B2(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_53),
.B(n_59),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_53),
.B1(n_99),
.B2(n_102),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_48),
.A2(n_53),
.B1(n_102),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_48),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_48),
.A2(n_53),
.B1(n_59),
.B2(n_141),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_48),
.A2(n_53),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_48),
.A2(n_53),
.B1(n_219),
.B2(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_48),
.B(n_121),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_48),
.A2(n_53),
.B1(n_186),
.B2(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_49),
.B(n_52),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_49),
.B(n_251),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g221 ( 
.A1(n_51),
.A2(n_55),
.A3(n_58),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_54)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_53),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_56),
.B1(n_64),
.B2(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_55),
.B(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_60),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_61),
.A2(n_71),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_61),
.A2(n_71),
.B1(n_112),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_61),
.A2(n_71),
.B1(n_182),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_61),
.A2(n_69),
.B1(n_71),
.B2(n_310),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_66),
.B(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_62),
.A2(n_66),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_62),
.A2(n_66),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_62),
.A2(n_66),
.B1(n_126),
.B2(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_62),
.A2(n_66),
.B1(n_194),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_67),
.Y(n_271)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_70),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_72),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_78),
.B1(n_115),
.B2(n_118),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_76),
.A2(n_78),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_326),
.B(n_332),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_303),
.A3(n_322),
.B1(n_324),
.B2(n_325),
.C(n_335),
.Y(n_82)
);

AOI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_152),
.A3(n_174),
.B1(n_297),
.B2(n_302),
.C(n_336),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_85),
.A2(n_298),
.B(n_301),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_133),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_86),
.B(n_133),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_113),
.C(n_128),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_87),
.B(n_128),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_103),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_104),
.C(n_109),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_98),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_89),
.B(n_98),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B1(n_94),
.B2(n_97),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_94),
.B1(n_97),
.B2(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_90),
.A2(n_94),
.B(n_130),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_90),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_90),
.A2(n_96),
.B1(n_239),
.B2(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_90),
.A2(n_233),
.B1(n_234),
.B2(n_273),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_93),
.B1(n_95),
.B2(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_91),
.A2(n_95),
.B1(n_124),
.B2(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_91),
.A2(n_95),
.B1(n_238),
.B2(n_240),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g234 ( 
.A(n_95),
.Y(n_234)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_96),
.B(n_121),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_100),
.A2(n_139),
.B1(n_142),
.B2(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_105),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_113),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.C(n_125),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_114),
.B(n_125),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_119),
.B(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_120),
.B(n_123),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_131),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_132),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_151),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_145),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_145),
.C(n_151),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_143),
.B2(n_144),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_136),
.B(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_139),
.A2(n_142),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_144),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_143),
.A2(n_166),
.B(n_169),
.Y(n_314)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_145),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.CI(n_150),
.CON(n_145),
.SN(n_145)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_148),
.C(n_150),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_153),
.B(n_154),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_172),
.B2(n_173),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_157),
.B(n_163),
.C(n_173),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_161),
.B(n_162),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_161),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_160),
.Y(n_310)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_162),
.B(n_305),
.CI(n_314),
.CON(n_304),
.SN(n_304)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_172),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_204),
.C(n_209),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_198),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_176),
.B(n_198),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_189),
.C(n_190),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_177),
.B(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_187),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_184),
.C(n_187),
.Y(n_201)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_295),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_189),
.Y(n_295)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.C(n_197),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_192),
.B(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_195),
.B(n_197),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_196),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_201),
.C(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_205),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_206),
.B(n_207),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_291),
.B(n_296),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_277),
.B(n_290),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_255),
.B(n_276),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_235),
.B(n_254),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_224),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_214),
.B(n_224),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_216),
.B1(n_220),
.B2(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_231),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_229),
.C(n_231),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_230),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_232),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_242),
.B(n_253),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_237),
.B(n_241),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_247),
.B(n_252),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_244),
.B(n_246),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_256),
.B(n_257),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_268),
.B1(n_274),
.B2(n_275),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_267),
.C(n_275),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_265),
.Y(n_287)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_268),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_272),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_279),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_286),
.C(n_288),
.Y(n_292)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_315),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_304),
.B(n_323),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_315),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_313),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_307),
.B1(n_317),
.B2(n_320),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_309),
.C(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_320),
.C(n_321),
.Y(n_327)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_308),
.Y(n_313)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule