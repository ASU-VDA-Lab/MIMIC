module fake_jpeg_17428_n_166 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_166);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx8_ASAP7_75t_SL g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_58),
.Y(n_91)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_54),
.B1(n_65),
.B2(n_59),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_0),
.B(n_1),
.Y(n_102)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_77),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_61),
.B1(n_54),
.B2(n_51),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_87),
.B1(n_0),
.B2(n_1),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_46),
.B(n_58),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_89),
.Y(n_101)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_64),
.B1(n_50),
.B2(n_62),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_53),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_91),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_60),
.B1(n_57),
.B2(n_63),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_96),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_56),
.C(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

HAxp5_ASAP7_75t_SL g99 ( 
.A(n_88),
.B(n_47),
.CON(n_99),
.SN(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_107),
.Y(n_117)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_103),
.B1(n_8),
.B2(n_9),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_2),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_108),
.B(n_8),
.Y(n_123)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_112),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_116),
.B(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_97),
.B(n_7),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_124),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_101),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_94),
.C(n_117),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_130),
.B1(n_124),
.B2(n_128),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_126),
.B(n_125),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_137),
.B1(n_109),
.B2(n_111),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_105),
.B1(n_104),
.B2(n_94),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_135),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_143),
.C(n_95),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_141),
.Y(n_144)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_146),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_143),
.A2(n_122),
.B1(n_118),
.B2(n_120),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_147),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_148),
.A2(n_98),
.B1(n_26),
.B2(n_10),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_151),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_149),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_144),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_144),
.B(n_153),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_27),
.B1(n_41),
.B2(n_13),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_25),
.B(n_39),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_23),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_31),
.B(n_38),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_22),
.B(n_37),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_21),
.C(n_35),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_19),
.B(n_34),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_164),
.A2(n_17),
.B1(n_32),
.B2(n_14),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_16),
.Y(n_166)
);


endmodule