module fake_jpeg_10790_n_631 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_631);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_631;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_10),
.B(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_4),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_60),
.Y(n_151)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_62),
.B(n_66),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_21),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_67),
.B(n_75),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_22),
.B(n_0),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_77),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_78),
.B(n_80),
.Y(n_162)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_82),
.Y(n_183)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_34),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_85),
.B(n_93),
.Y(n_168)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_88),
.Y(n_202)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_1),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_43),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

INVx11_ASAP7_75t_SL g98 ( 
.A(n_59),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_100),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_101),
.Y(n_212)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_102),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_104),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_22),
.B(n_3),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_105),
.B(n_106),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_26),
.B(n_3),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_20),
.Y(n_110)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_41),
.Y(n_112)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_31),
.Y(n_114)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_37),
.Y(n_117)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_23),
.Y(n_121)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_35),
.Y(n_122)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_35),
.Y(n_123)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_54),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_52),
.Y(n_137)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_35),
.Y(n_125)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_31),
.Y(n_126)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_31),
.Y(n_127)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_37),
.Y(n_128)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_128),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_125),
.B1(n_101),
.B2(n_99),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_135),
.A2(n_142),
.B1(n_122),
.B2(n_123),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_26),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_136),
.B(n_144),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_137),
.B(n_187),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_37),
.B1(n_56),
.B2(n_36),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_55),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_109),
.A2(n_49),
.B1(n_56),
.B2(n_36),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_148),
.A2(n_154),
.B1(n_204),
.B2(n_210),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_86),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_110),
.A2(n_49),
.B1(n_56),
.B2(n_36),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_88),
.B(n_58),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g246 ( 
.A1(n_159),
.A2(n_191),
.B(n_130),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_76),
.B(n_29),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_165),
.B(n_201),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_98),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_166),
.B(n_208),
.Y(n_257)
);

AOI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_72),
.A2(n_33),
.B(n_54),
.Y(n_186)
);

NAND2xp67_ASAP7_75t_SL g238 ( 
.A(n_186),
.B(n_5),
.Y(n_238)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_203),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_63),
.B(n_50),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g197 ( 
.A(n_65),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_103),
.B(n_55),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_68),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_115),
.A2(n_47),
.B1(n_45),
.B2(n_49),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_73),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_71),
.B(n_40),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_119),
.A2(n_45),
.B1(n_47),
.B2(n_29),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_73),
.Y(n_211)
);

CKINVDCx6p67_ASAP7_75t_R g248 ( 
.A(n_211),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_81),
.A2(n_45),
.B1(n_47),
.B2(n_58),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_215),
.A2(n_80),
.B1(n_82),
.B2(n_53),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_SL g321 ( 
.A1(n_216),
.A2(n_223),
.B(n_238),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_133),
.B(n_53),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_218),
.B(n_222),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_219),
.A2(n_229),
.B1(n_260),
.B2(n_265),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_221),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_133),
.B(n_50),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_40),
.B1(n_121),
.B2(n_89),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_4),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_224),
.B(n_252),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_202),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_226),
.B(n_264),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_172),
.A2(n_174),
.B1(n_156),
.B2(n_194),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_135),
.A2(n_33),
.B1(n_6),
.B2(n_7),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_228),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_168),
.A2(n_33),
.B1(n_6),
.B2(n_7),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_172),
.A2(n_174),
.B1(n_141),
.B2(n_139),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_230),
.A2(n_273),
.B1(n_281),
.B2(n_286),
.Y(n_341)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_231),
.Y(n_329)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_232),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_233),
.Y(n_322)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_234),
.Y(n_326)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_239),
.Y(n_305)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_178),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_240),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_130),
.B(n_5),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_241),
.B(n_250),
.Y(n_340)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_242),
.Y(n_298)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_138),
.Y(n_244)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_244),
.Y(n_333)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_246),
.Y(n_325)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_138),
.Y(n_247)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_247),
.Y(n_346)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_5),
.Y(n_250)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_189),
.Y(n_251)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_251),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_5),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_175),
.Y(n_253)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_253),
.Y(n_293)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

INVx2_ASAP7_75t_R g255 ( 
.A(n_211),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_255),
.B(n_256),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_129),
.B(n_6),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_132),
.B(n_7),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_267),
.Y(n_304)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_199),
.Y(n_259)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_151),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_178),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g343 ( 
.A(n_261),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_159),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_262),
.A2(n_290),
.B1(n_287),
.B2(n_216),
.Y(n_292)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_161),
.Y(n_263)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_263),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_147),
.B(n_11),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_169),
.A2(n_18),
.B1(n_13),
.B2(n_15),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

INVx11_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_158),
.B(n_12),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_173),
.B(n_17),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_268),
.B(n_270),
.C(n_176),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_167),
.B(n_17),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_271),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_181),
.B(n_17),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_171),
.B(n_17),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_185),
.Y(n_272)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_160),
.A2(n_198),
.B1(n_134),
.B2(n_150),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_162),
.B(n_18),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_284),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_162),
.B(n_157),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_276),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_197),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_277),
.B(n_280),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_131),
.B(n_143),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_164),
.A2(n_177),
.B1(n_213),
.B2(n_149),
.Y(n_281)
);

O2A1O1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_152),
.A2(n_206),
.B(n_145),
.C(n_164),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_287),
.B(n_219),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_157),
.B(n_163),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_283),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_170),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_184),
.B(n_188),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_285),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_157),
.A2(n_195),
.B1(n_192),
.B2(n_183),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_140),
.A2(n_146),
.B1(n_153),
.B2(n_214),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_192),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_207),
.Y(n_314)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_214),
.Y(n_289)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_289),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_195),
.A2(n_140),
.B1(n_146),
.B2(n_153),
.Y(n_290)
);

AOI32xp33_ASAP7_75t_L g291 ( 
.A1(n_218),
.A2(n_161),
.A3(n_176),
.B1(n_179),
.B2(n_183),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_291),
.A2(n_282),
.B(n_248),
.C(n_263),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_292),
.A2(n_242),
.B1(n_261),
.B2(n_243),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_301),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_235),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_314),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_258),
.B(n_212),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_317),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_267),
.B(n_279),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_225),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_320),
.B(n_344),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_238),
.A2(n_179),
.B(n_212),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_330),
.A2(n_301),
.B(n_341),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_237),
.A2(n_228),
.B1(n_229),
.B2(n_265),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_331),
.A2(n_303),
.B1(n_300),
.B2(n_237),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_274),
.B(n_268),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_338),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_246),
.B(n_236),
.C(n_245),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_336),
.C(n_332),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_222),
.B(n_224),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_268),
.B(n_270),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_270),
.B(n_252),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_345),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_239),
.B(n_259),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_254),
.B(n_217),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_295),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_257),
.A2(n_221),
.B1(n_244),
.B2(n_233),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_349),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_345),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_350),
.B(n_362),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_351),
.A2(n_367),
.B1(n_373),
.B2(n_385),
.Y(n_396)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_305),
.Y(n_354)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_356),
.B(n_336),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_284),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_357),
.B(n_363),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_304),
.B(n_234),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_358),
.B(n_365),
.Y(n_405)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_305),
.Y(n_359)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_359),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_314),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_308),
.B(n_220),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_300),
.A2(n_260),
.B1(n_288),
.B2(n_221),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_366),
.A2(n_386),
.B(n_322),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_303),
.A2(n_228),
.B1(n_289),
.B2(n_231),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_220),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_368),
.B(n_379),
.Y(n_431)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_369),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_370),
.A2(n_299),
.B(n_328),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_334),
.B(n_272),
.C(n_276),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_320),
.C(n_311),
.Y(n_399)
);

INVx13_ASAP7_75t_L g372 ( 
.A(n_318),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_372),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_330),
.A2(n_228),
.B1(n_251),
.B2(n_278),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_323),
.Y(n_374)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_374),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_304),
.B(n_253),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_375),
.B(n_376),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_315),
.B(n_255),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_378),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_309),
.B(n_232),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_324),
.B(n_248),
.Y(n_379)
);

INVx13_ASAP7_75t_L g380 ( 
.A(n_318),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_380),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_309),
.B(n_249),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_381),
.B(n_383),
.Y(n_423)
);

INVx13_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_382),
.Y(n_414)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_325),
.B(n_248),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_306),
.Y(n_384)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_384),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_317),
.A2(n_247),
.B1(n_248),
.B2(n_243),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_340),
.B(n_240),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_387),
.A2(n_294),
.B1(n_337),
.B2(n_339),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_295),
.B(n_243),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_388),
.B(n_322),
.Y(n_419)
);

AO22x1_ASAP7_75t_SL g389 ( 
.A1(n_292),
.A2(n_266),
.B1(n_321),
.B2(n_306),
.Y(n_389)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_338),
.B(n_266),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_R g411 ( 
.A(n_390),
.B(n_342),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_327),
.Y(n_418)
);

INVx13_ASAP7_75t_L g393 ( 
.A(n_343),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_393),
.Y(n_422)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_394),
.A2(n_343),
.B1(n_335),
.B2(n_329),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_395),
.A2(n_404),
.B(n_410),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_367),
.A2(n_299),
.B1(n_312),
.B2(n_333),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_398),
.A2(n_416),
.B1(n_427),
.B2(n_387),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_399),
.B(n_402),
.C(n_403),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_400),
.A2(n_401),
.B1(n_391),
.B2(n_350),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_352),
.A2(n_310),
.B1(n_302),
.B2(n_294),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_302),
.C(n_311),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_370),
.A2(n_296),
.B(n_298),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_356),
.B(n_297),
.C(n_293),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_407),
.B(n_408),
.C(n_424),
.Y(n_454)
);

MAJx2_ASAP7_75t_L g408 ( 
.A(n_360),
.B(n_327),
.C(n_348),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_364),
.A2(n_298),
.B(n_342),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_411),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_351),
.A2(n_337),
.B1(n_339),
.B2(n_346),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_418),
.B(n_390),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_419),
.A2(n_425),
.B(n_429),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_420),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_360),
.B(n_307),
.Y(n_424)
);

OAI22x1_ASAP7_75t_L g425 ( 
.A1(n_352),
.A2(n_346),
.B1(n_329),
.B2(n_326),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_377),
.A2(n_335),
.B(n_343),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_430),
.B(n_391),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_433),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_405),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_434),
.B(n_457),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_353),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_435),
.B(n_436),
.C(n_438),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_353),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_397),
.Y(n_437)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_437),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_371),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_419),
.Y(n_439)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_439),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_440),
.Y(n_490)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_397),
.Y(n_441)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_441),
.Y(n_471)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_443),
.Y(n_484)
);

NOR3xp33_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_357),
.C(n_386),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_445),
.B(n_456),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_399),
.B(n_365),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_452),
.C(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_406),
.Y(n_448)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_448),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_395),
.A2(n_362),
.B(n_378),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_449),
.Y(n_491)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_406),
.Y(n_450)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_450),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_361),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_407),
.B(n_361),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_430),
.A2(n_373),
.B1(n_375),
.B2(n_389),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_455),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_415),
.B(n_388),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_412),
.B(n_355),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_421),
.A2(n_389),
.B1(n_381),
.B2(n_383),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_458),
.A2(n_421),
.B1(n_417),
.B2(n_423),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_405),
.B(n_358),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_459),
.Y(n_492)
);

OR2x4_ASAP7_75t_L g460 ( 
.A(n_411),
.B(n_389),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_460),
.B(n_366),
.Y(n_500)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_431),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_465),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_463),
.B(n_401),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_419),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_464),
.B(n_467),
.Y(n_476)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_426),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_355),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_431),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_468),
.B(n_470),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_469),
.A2(n_368),
.B1(n_409),
.B2(n_359),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_438),
.B(n_423),
.Y(n_470)
);

FAx1_ASAP7_75t_SL g474 ( 
.A(n_459),
.B(n_417),
.CI(n_408),
.CON(n_474),
.SN(n_474)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_474),
.B(n_475),
.Y(n_526)
);

XOR2x2_ASAP7_75t_L g475 ( 
.A(n_463),
.B(n_396),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_435),
.B(n_363),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_494),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_442),
.A2(n_446),
.B(n_444),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_480),
.A2(n_495),
.B(n_500),
.Y(n_518)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_483),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_447),
.B(n_412),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_485),
.B(n_496),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_439),
.A2(n_400),
.B1(n_396),
.B2(n_429),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_486),
.A2(n_432),
.B1(n_422),
.B2(n_414),
.Y(n_524)
);

OAI21x1_ASAP7_75t_R g487 ( 
.A1(n_462),
.A2(n_404),
.B(n_414),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_487),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_433),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_442),
.A2(n_420),
.B(n_410),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_379),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_433),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_497),
.B(n_425),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_SL g502 ( 
.A(n_473),
.B(n_451),
.C(n_444),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_502),
.A2(n_514),
.B1(n_491),
.B2(n_495),
.Y(n_533)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_477),
.Y(n_503)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_503),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_472),
.B(n_451),
.C(n_454),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_504),
.B(n_507),
.C(n_513),
.Y(n_531)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_476),
.Y(n_506)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_506),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_454),
.C(n_436),
.Y(n_507)
);

XNOR2x1_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_458),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_527),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_482),
.B(n_449),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_510),
.B(n_511),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_482),
.B(n_452),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_490),
.A2(n_446),
.B1(n_455),
.B2(n_462),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_512),
.A2(n_516),
.B1(n_521),
.B2(n_486),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_468),
.B(n_408),
.C(n_443),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_490),
.A2(n_493),
.B1(n_484),
.B2(n_491),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_475),
.B(n_376),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_515),
.B(n_474),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_493),
.A2(n_460),
.B1(n_437),
.B2(n_383),
.Y(n_516)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_517),
.Y(n_540)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_471),
.Y(n_520)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_520),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_484),
.A2(n_385),
.B1(n_432),
.B2(n_416),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_522),
.A2(n_524),
.B1(n_481),
.B2(n_525),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_475),
.B(n_409),
.C(n_425),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_489),
.C(n_492),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_469),
.B(n_354),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_499),
.A2(n_422),
.B1(n_413),
.B2(n_384),
.Y(n_528)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_528),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_497),
.B(n_394),
.Y(n_529)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_529),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_532),
.A2(n_523),
.B1(n_527),
.B2(n_518),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_533),
.Y(n_564)
);

FAx1_ASAP7_75t_SL g537 ( 
.A(n_526),
.B(n_474),
.CI(n_480),
.CON(n_537),
.SN(n_537)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_537),
.B(n_549),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_538),
.A2(n_512),
.B1(n_516),
.B2(n_518),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_501),
.B(n_499),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_539),
.B(n_550),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_481),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_541),
.B(n_542),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_507),
.B(n_489),
.C(n_492),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_544),
.B(n_545),
.C(n_546),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_487),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_504),
.B(n_479),
.C(n_487),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_508),
.B(n_500),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_505),
.B(n_498),
.Y(n_551)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_551),
.Y(n_573)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_529),
.Y(n_552)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_552),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_514),
.A2(n_498),
.B1(n_488),
.B2(n_471),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_553),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_555),
.A2(n_569),
.B1(n_571),
.B2(n_394),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_538),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_557),
.B(n_560),
.Y(n_589)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_543),
.Y(n_558)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_558),
.Y(n_588)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_540),
.Y(n_559)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_559),
.Y(n_590)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_548),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_562),
.B(n_550),
.Y(n_579)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_547),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_566),
.B(n_567),
.Y(n_575)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_536),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_544),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_568),
.B(n_570),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_542),
.A2(n_529),
.B(n_515),
.Y(n_569)
);

OAI21xp33_ASAP7_75t_L g570 ( 
.A1(n_537),
.A2(n_509),
.B(n_519),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_546),
.A2(n_513),
.B1(n_505),
.B2(n_479),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_563),
.B(n_531),
.C(n_534),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_574),
.B(n_576),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_563),
.B(n_531),
.C(n_534),
.Y(n_576)
);

FAx1_ASAP7_75t_SL g578 ( 
.A(n_572),
.B(n_537),
.CI(n_549),
.CON(n_578),
.SN(n_578)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_578),
.B(n_585),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_579),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_556),
.B(n_541),
.C(n_551),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_580),
.B(n_582),
.C(n_583),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_SL g581 ( 
.A(n_565),
.B(n_545),
.C(n_530),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_581),
.B(n_569),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_556),
.B(n_535),
.C(n_521),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_571),
.B(n_535),
.C(n_488),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_564),
.B(n_413),
.C(n_369),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_584),
.B(n_587),
.C(n_554),
.Y(n_600)
);

FAx1_ASAP7_75t_SL g585 ( 
.A(n_572),
.B(n_372),
.CI(n_380),
.CON(n_585),
.SN(n_585)
);

AOI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_586),
.A2(n_562),
.B1(n_582),
.B2(n_584),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_564),
.B(n_326),
.C(n_382),
.Y(n_587)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_588),
.Y(n_591)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_591),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_575),
.A2(n_561),
.B1(n_566),
.B2(n_559),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_592),
.B(n_596),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_597),
.B(n_585),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_574),
.B(n_567),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_599),
.B(n_603),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_600),
.B(n_587),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_576),
.B(n_573),
.C(n_555),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_601),
.B(n_602),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_577),
.B(n_573),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_578),
.B(n_558),
.Y(n_603)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_604),
.Y(n_617)
);

AOI31xp67_ASAP7_75t_L g605 ( 
.A1(n_595),
.A2(n_575),
.A3(n_589),
.B(n_590),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_605),
.B(n_560),
.C(n_600),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_601),
.A2(n_583),
.B(n_580),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_607),
.B(n_608),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_579),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_593),
.B(n_554),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_610),
.B(n_593),
.Y(n_614)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_613),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_614),
.B(n_618),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_615),
.A2(n_612),
.B1(n_594),
.B2(n_609),
.Y(n_621)
);

BUFx24_ASAP7_75t_SL g618 ( 
.A(n_606),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_SL g619 ( 
.A1(n_611),
.A2(n_594),
.B1(n_596),
.B2(n_372),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_619),
.A2(n_613),
.B1(n_604),
.B2(n_380),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_621),
.B(n_622),
.Y(n_626)
);

AO21x2_ASAP7_75t_SL g623 ( 
.A1(n_620),
.A2(n_382),
.B(n_393),
.Y(n_623)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_623),
.A2(n_393),
.B(n_617),
.C(n_619),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_625),
.B(n_623),
.Y(n_627)
);

AO21x1_ASAP7_75t_L g628 ( 
.A1(n_627),
.A2(n_626),
.B(n_621),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_628),
.B(n_624),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_629),
.B(n_616),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_630),
.B(n_623),
.Y(n_631)
);


endmodule