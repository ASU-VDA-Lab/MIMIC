module fake_jpeg_15647_n_172 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_35),
.Y(n_40)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_41),
.B1(n_43),
.B2(n_47),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_23),
.B1(n_31),
.B2(n_34),
.Y(n_41)
);

HAxp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_22),
.CON(n_42),
.SN(n_42)
);

NAND3xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_39),
.C(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_43)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_29),
.B(n_25),
.CI(n_26),
.CON(n_45),
.SN(n_45)
);

NOR2xp67_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_21),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_14),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_13),
.B1(n_25),
.B2(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_20),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_28),
.B1(n_31),
.B2(n_27),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_56),
.B1(n_36),
.B2(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_55),
.Y(n_73)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_59),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_60),
.B(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_61),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_18),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_74),
.B(n_51),
.C(n_27),
.D(n_65),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_56),
.B(n_52),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_32),
.B(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_44),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_43),
.B1(n_47),
.B2(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_72),
.Y(n_88)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_37),
.A3(n_32),
.B1(n_27),
.B2(n_49),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_52),
.B1(n_48),
.B2(n_34),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_78),
.B1(n_48),
.B2(n_54),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_48),
.B1(n_44),
.B2(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_90),
.B1(n_94),
.B2(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_67),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_79),
.Y(n_108)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_93),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_63),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_53),
.B1(n_37),
.B2(n_65),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_96),
.B(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_105),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_69),
.C(n_70),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_101),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_74),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_109),
.B1(n_85),
.B2(n_101),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_88),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_93),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_76),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_18),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_32),
.B(n_77),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_122),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_85),
.B1(n_94),
.B2(n_90),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_124),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_95),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_111),
.Y(n_121)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_79),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_110),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_108),
.C(n_14),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_113),
.C(n_122),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_32),
.C(n_110),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_135),
.C(n_16),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_79),
.C(n_26),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_124),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_139),
.C(n_143),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_115),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_140),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_146),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_119),
.B1(n_123),
.B2(n_12),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_16),
.C(n_12),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_145),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

OAI21x1_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_126),
.B(n_136),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_4),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_144),
.A2(n_132),
.B1(n_134),
.B2(n_133),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_1),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_156),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_1),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_1),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_153),
.B(n_152),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_148),
.C(n_5),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_154),
.B(n_5),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_4),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_159),
.A2(n_148),
.B1(n_5),
.B2(n_6),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_165),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_167),
.C(n_8),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_6),
.B(n_8),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_162),
.B(n_8),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_169),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_170),
.Y(n_172)
);


endmodule