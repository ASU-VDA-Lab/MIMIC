module fake_jpeg_5360_n_181 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_181);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_SL g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx12_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_31),
.Y(n_40)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_32),
.B1(n_24),
.B2(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_0),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_13),
.B1(n_20),
.B2(n_22),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_49),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_17),
.B1(n_25),
.B2(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_13),
.B1(n_25),
.B2(n_17),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_16),
.B1(n_24),
.B2(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_14),
.Y(n_60)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_33),
.B1(n_27),
.B2(n_15),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_33),
.B1(n_32),
.B2(n_29),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_44),
.B1(n_40),
.B2(n_43),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_19),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_63),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_42),
.B1(n_37),
.B2(n_39),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_41),
.B1(n_32),
.B2(n_49),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_47),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_19),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_27),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_40),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_53),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_72),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_62),
.B1(n_64),
.B2(n_58),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_80),
.B1(n_58),
.B2(n_62),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_46),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_65),
.C(n_54),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_43),
.B1(n_45),
.B2(n_35),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_65),
.B1(n_60),
.B2(n_51),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_82),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_66),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_94),
.B1(n_96),
.B2(n_92),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_64),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_72),
.B(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_26),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_26),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

AO21x2_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_59),
.B(n_68),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_108),
.B(n_114),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_91),
.C(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_98),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_78),
.B(n_76),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_113),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_70),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_56),
.A3(n_34),
.B1(n_35),
.B2(n_29),
.C1(n_31),
.C2(n_26),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_15),
.B(n_19),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_116),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_128),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_123),
.C(n_127),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_103),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_96),
.C(n_87),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_85),
.B(n_90),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_126),
.B(n_103),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_61),
.B(n_70),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_34),
.C(n_35),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_120),
.Y(n_140)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_133),
.B1(n_35),
.B2(n_34),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_126),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_103),
.B1(n_99),
.B2(n_112),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_31),
.B(n_29),
.C(n_26),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_140),
.B1(n_141),
.B2(n_127),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_100),
.C(n_108),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_123),
.C(n_124),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_26),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_103),
.B1(n_114),
.B2(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_145),
.C(n_151),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_124),
.C(n_115),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_138),
.A2(n_120),
.B1(n_115),
.B2(n_56),
.Y(n_146)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_56),
.B1(n_3),
.B2(n_4),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_150),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_148),
.A2(n_149),
.B1(n_130),
.B2(n_139),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_48),
.Y(n_151)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_137),
.C(n_134),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_156),
.C(n_157),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_132),
.C(n_135),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_48),
.C(n_31),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_31),
.C(n_26),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_158),
.B(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_6),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_167),
.Y(n_168)
);

OAI211xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_164),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_11),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_2),
.B(n_5),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_171),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_163),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_166),
.B(n_6),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_174),
.B1(n_10),
.B2(n_176),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_7),
.C(n_8),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_168),
.B(n_7),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_SL g177 ( 
.A1(n_175),
.A2(n_8),
.B(n_9),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_10),
.Y(n_181)
);


endmodule