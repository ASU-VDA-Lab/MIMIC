module fake_jpeg_15062_n_146 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_146);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_21),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_28),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_27),
.B(n_23),
.C(n_16),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_17),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_29),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_29),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_29),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_30),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_32),
.A2(n_14),
.B1(n_16),
.B2(n_25),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_63),
.B1(n_18),
.B2(n_20),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_14),
.B1(n_25),
.B2(n_22),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_22),
.B(n_20),
.C(n_18),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_79),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_1),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_72),
.Y(n_99)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_24),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_45),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_74),
.Y(n_95)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_50),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_93),
.Y(n_101)
);

OAI22x1_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_26),
.B1(n_58),
.B2(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_92),
.B1(n_100),
.B2(n_99),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_49),
.B1(n_45),
.B2(n_51),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_58),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_79),
.C(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_107),
.C(n_113),
.Y(n_114)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_70),
.B(n_67),
.Y(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_111),
.B(n_85),
.C(n_26),
.D(n_46),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_68),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_68),
.B1(n_72),
.B2(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_92),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_80),
.B1(n_66),
.B2(n_50),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_77),
.B1(n_65),
.B2(n_66),
.Y(n_110)
);

NOR4xp25_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_72),
.C(n_58),
.D(n_74),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_26),
.C(n_46),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_120),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_105),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_90),
.C(n_87),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_106),
.C(n_104),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_102),
.A2(n_100),
.B1(n_87),
.B2(n_85),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_108),
.B(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_109),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_113),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_118),
.B1(n_4),
.B2(n_5),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_114),
.C(n_106),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_114),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_126),
.B(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_2),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_116),
.B(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_131),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_134),
.Y(n_137)
);

AOI31xp67_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_123),
.A3(n_127),
.B(n_129),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

XOR2x2_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_131),
.C(n_124),
.Y(n_139)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_138),
.A3(n_137),
.B1(n_134),
.B2(n_125),
.C1(n_11),
.C2(n_12),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_9),
.C1(n_11),
.C2(n_140),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_143),
.C(n_3),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_3),
.Y(n_146)
);


endmodule