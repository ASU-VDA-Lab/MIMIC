module real_jpeg_10394_n_17 (n_8, n_0, n_2, n_10, n_9, n_333, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_334, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_333;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_334;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_1),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_1),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_1),
.A2(n_16),
.B(n_35),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_2),
.A2(n_37),
.B1(n_69),
.B2(n_72),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_2),
.A2(n_37),
.B1(n_46),
.B2(n_47),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_3),
.A2(n_61),
.B1(n_69),
.B2(n_72),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_61),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g125 ( 
.A(n_4),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_9),
.A2(n_50),
.B1(n_69),
.B2(n_72),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_10),
.A2(n_28),
.B1(n_69),
.B2(n_72),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_10),
.A2(n_28),
.B1(n_46),
.B2(n_47),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_11),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_11),
.A2(n_69),
.B1(n_72),
.B2(n_84),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_84),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_84),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_12),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_12),
.A2(n_69),
.B1(n_72),
.B2(n_105),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_105),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_105),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_13),
.A2(n_69),
.B1(n_72),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_13),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_122),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_122),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_122),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_14),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_14),
.A2(n_69),
.B1(n_72),
.B2(n_117),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_117),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_117),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_16),
.A2(n_47),
.B(n_64),
.C(n_102),
.D(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_16),
.B(n_47),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_16),
.B(n_45),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_16),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_16),
.A2(n_123),
.B(n_126),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_16),
.A2(n_34),
.B(n_41),
.C(n_158),
.D(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_16),
.B(n_34),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_16),
.B(n_38),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_16),
.A2(n_26),
.B1(n_27),
.B2(n_139),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_90),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_20),
.B(n_76),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_51),
.B1(n_52),
.B2(n_75),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_21),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_39),
.B2(n_40),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_25),
.A2(n_30),
.B1(n_33),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_31),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_27),
.A2(n_31),
.B(n_139),
.C(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_29),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_29),
.B(n_220),
.Y(n_229)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_30),
.A2(n_33),
.B1(n_60),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_30),
.A2(n_33),
.B1(n_228),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_30),
.A2(n_219),
.B(n_257),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_33),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_33),
.A2(n_83),
.B(n_229),
.Y(n_299)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_38),
.B(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_48),
.Y(n_40)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_41),
.B(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_41),
.A2(n_45),
.B1(n_254),
.B2(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_41),
.A2(n_45),
.B1(n_89),
.B2(n_273),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_42),
.B(n_47),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_44),
.A2(n_46),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_65),
.B(n_67),
.C(n_68),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_65),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.C(n_62),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_54),
.B1(n_62),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_55),
.A2(n_57),
.B1(n_178),
.B2(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_55),
.A2(n_214),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_57),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_57),
.A2(n_178),
.B(n_179),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_57),
.A2(n_179),
.B(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_59),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_62),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_73),
.B(n_74),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_63),
.A2(n_73),
.B1(n_116),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_63),
.A2(n_156),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_63),
.A2(n_73),
.B1(n_211),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_63),
.A2(n_73),
.B1(n_239),
.B2(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_63),
.A2(n_73),
.B1(n_248),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_64),
.B(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_64),
.A2(n_68),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_72),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_65),
.B(n_72),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_67),
.A2(n_69),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_69),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_72),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_72),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_116),
.B(n_118),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_73),
.B(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_73),
.A2(n_118),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_74),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.C(n_85),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_318),
.Y(n_324)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.C(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_82),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_82),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_85),
.B(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI321xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_315),
.A3(n_325),
.B1(n_330),
.B2(n_331),
.C(n_333),
.Y(n_92)
);

AOI321xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_265),
.A3(n_303),
.B1(n_309),
.B2(n_314),
.C(n_334),
.Y(n_93)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_222),
.C(n_261),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_193),
.B(n_221),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_172),
.B(n_192),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_150),
.B(n_171),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_128),
.B(n_149),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_110),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_100),
.B(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_106),
.B1(n_107),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_103),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_115),
.C(n_120),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_123),
.B(n_126),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_123),
.A2(n_141),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_123),
.A2(n_141),
.B1(n_204),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_123),
.A2(n_141),
.B1(n_237),
.B2(n_246),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_123),
.A2(n_141),
.B(n_246),
.Y(n_278)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_124),
.A2(n_125),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_124),
.B(n_127),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_124),
.A2(n_125),
.B1(n_169),
.B2(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_136),
.B(n_148),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_134),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_143),
.B(n_147),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_140),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_141),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_142),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_152),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_163),
.B2(n_170),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_155),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_162),
.C(n_170),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_159),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_167),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_174),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_186),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_188),
.C(n_190),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_181),
.B2(n_185),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_182),
.C(n_183),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_187),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_188),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_194),
.B(n_195),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_208),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_197),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_197),
.B(n_207),
.C(n_208),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_202),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_205),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_216),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_210),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_215),
.C(n_216),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g310 ( 
.A1(n_223),
.A2(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_241),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_224),
.B(n_241),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.C(n_240),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_227),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_233),
.C(n_234),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_240),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_238),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_259),
.B2(n_260),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_249),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_244),
.B(n_249),
.C(n_260),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_247),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_255),
.C(n_258),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_252),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_263),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_283),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_266),
.B(n_283),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_276),
.C(n_282),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_267),
.A2(n_268),
.B1(n_276),
.B2(n_308),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_272),
.C(n_274),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_276),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_281),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_277),
.A2(n_278),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_277),
.A2(n_295),
.B(n_299),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_279),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_279),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_280),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_307),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_301),
.B2(n_302),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_293),
.B2(n_294),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_294),
.C(n_302),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_291),
.B(n_292),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_291),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_292),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_292),
.A2(n_317),
.B1(n_321),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_300),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_297),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_301),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_304),
.A2(n_310),
.B(n_313),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_323),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_323),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_321),
.C(n_322),
.Y(n_316)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);


endmodule