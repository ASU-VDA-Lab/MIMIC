module fake_jpeg_25172_n_249 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_21),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_61),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_35),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_27),
.C(n_30),
.Y(n_83)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_33),
.B1(n_31),
.B2(n_18),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_64),
.B1(n_32),
.B2(n_25),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_23),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_33),
.B1(n_18),
.B2(n_23),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_18),
.B1(n_33),
.B2(n_24),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_29),
.B1(n_19),
.B2(n_34),
.Y(n_87)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_1),
.C(n_3),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_69),
.B(n_84),
.C(n_3),
.Y(n_114)
);

AO22x1_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_40),
.B1(n_38),
.B2(n_44),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_66),
.B(n_68),
.Y(n_110)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_82),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_40),
.B1(n_27),
.B2(n_30),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_93),
.B1(n_60),
.B2(n_47),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_28),
.B1(n_24),
.B2(n_29),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_55),
.B1(n_56),
.B2(n_5),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_90),
.Y(n_96)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_28),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_19),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_44),
.B1(n_41),
.B2(n_30),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_50),
.B(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_51),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_27),
.B1(n_34),
.B2(n_25),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_96),
.B1(n_99),
.B2(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_107),
.Y(n_129)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_60),
.B1(n_52),
.B2(n_63),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_4),
.Y(n_142)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_105),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_59),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_108),
.B(n_81),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_52),
.B1(n_63),
.B2(n_49),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_80),
.B1(n_89),
.B2(n_75),
.Y(n_127)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_71),
.B(n_54),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_67),
.B(n_49),
.C(n_68),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_73),
.B1(n_85),
.B2(n_53),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_78),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_115),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_114),
.A2(n_53),
.B1(n_5),
.B2(n_6),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_4),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_87),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_124),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_134),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_94),
.Y(n_152)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_130),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_132),
.B1(n_139),
.B2(n_141),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_114),
.C(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_81),
.B1(n_92),
.B2(n_66),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_100),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_102),
.B(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_142),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_92),
.B1(n_74),
.B2(n_7),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_4),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_137),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_74),
.B1(n_6),
.B2(n_7),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_96),
.B1(n_107),
.B2(n_104),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_139),
.B1(n_138),
.B2(n_119),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_102),
.C(n_96),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_158),
.C(n_161),
.Y(n_177)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_155),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_148),
.B(n_8),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_151),
.B(n_154),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_153),
.B(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_164),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_102),
.C(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_95),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_165),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_108),
.C(n_113),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_121),
.A2(n_119),
.B(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_137),
.B(n_115),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_178),
.B1(n_166),
.B2(n_183),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_144),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_169),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_123),
.B1(n_108),
.B2(n_142),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_171),
.A2(n_178),
.B1(n_160),
.B2(n_10),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_173),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_142),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_185),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_123),
.B(n_130),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_175),
.A2(n_180),
.B(n_182),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_123),
.B1(n_124),
.B2(n_105),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_149),
.A2(n_98),
.B(n_101),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_8),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_120),
.B(n_9),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_106),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_106),
.B1(n_120),
.B2(n_10),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_155),
.B1(n_154),
.B2(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_193),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_191),
.B1(n_196),
.B2(n_203),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_143),
.B1(n_151),
.B2(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_161),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_176),
.B1(n_168),
.B2(n_182),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_166),
.B1(n_163),
.B2(n_150),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_159),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_201),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_202),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_145),
.C(n_150),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_173),
.C(n_168),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_145),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_210),
.C(n_197),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_179),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_176),
.C(n_175),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_172),
.B(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_179),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_193),
.B1(n_194),
.B2(n_200),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_202),
.B(n_203),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_221),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_219),
.A2(n_223),
.B(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_220),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_226),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_194),
.B(n_195),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_186),
.B1(n_171),
.B2(n_201),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_212),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_204),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_228),
.B(n_232),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_231),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_211),
.Y(n_232)
);

NAND4xp25_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_9),
.C(n_12),
.D(n_13),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g239 ( 
.A(n_233),
.Y(n_239)
);

AOI21x1_ASAP7_75t_SL g240 ( 
.A1(n_234),
.A2(n_225),
.B(n_222),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_223),
.B(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_229),
.A2(n_226),
.B1(n_218),
.B2(n_234),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_240),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_230),
.C(n_206),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_244),
.B(n_239),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_230),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_246),
.B(n_241),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_233),
.B(n_15),
.C(n_16),
.Y(n_246)
);

OAI311xp33_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_14),
.A3(n_16),
.B1(n_239),
.C1(n_246),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_14),
.Y(n_249)
);


endmodule