module real_jpeg_17325_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OA22x2_ASAP7_75t_L g12 ( 
.A1(n_0),
.A2(n_3),
.B1(n_13),
.B2(n_14),
.Y(n_12)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

AO22x1_ASAP7_75t_SL g18 ( 
.A1(n_0),
.A2(n_5),
.B1(n_14),
.B2(n_19),
.Y(n_18)
);

INVx2_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

OR2x4_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_20),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_20),
.Y(n_29)
);

INVx2_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

A2O1A1O1Ixp25_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_8),
.B(n_21),
.C(n_23),
.D(n_25),
.Y(n_6)
);

OR2x4_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_20),
.Y(n_22)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_20),
.Y(n_9)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_15),
.B(n_16),
.Y(n_10)
);

INVx1_ASAP7_75t_SL g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_15),
.B(n_17),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_15),
.A2(n_18),
.B(n_31),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);


endmodule