module real_jpeg_5758_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_1),
.B(n_37),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_1),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_1),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_1),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_1),
.B(n_81),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_1),
.B(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_2),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_2),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_3),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_3),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_3),
.B(n_128),
.Y(n_127)
);

NAND2x1p5_ASAP7_75t_L g170 ( 
.A(n_3),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_3),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_4),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_4),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_4),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_5),
.B(n_61),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_5),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_5),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_5),
.B(n_114),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_5),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_5),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_6),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_6),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_6),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_6),
.B(n_145),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_6),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_6),
.B(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_6),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_6),
.B(n_380),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_7),
.Y(n_187)
);

INVx8_ASAP7_75t_L g276 ( 
.A(n_7),
.Y(n_276)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_8),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_9),
.B(n_37),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_9),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_9),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_9),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_9),
.B(n_260),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_9),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_9),
.B(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_10),
.B(n_36),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_10),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_10),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_10),
.B(n_367),
.Y(n_366)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_11),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_11),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_11),
.Y(n_361)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_13),
.Y(n_193)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_13),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_13),
.Y(n_269)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_13),
.Y(n_329)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_13),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_14),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_14),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_14),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_14),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_14),
.B(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_15),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_15),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_16),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_16),
.B(n_114),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_16),
.B(n_173),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_16),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_17),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_17),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_17),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_17),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_17),
.B(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_340),
.Y(n_18)
);

AOI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_296),
.B(n_339),
.Y(n_19)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_249),
.B(n_295),
.Y(n_20)
);

AOI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_205),
.B(n_248),
.Y(n_21)
);

OAI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_157),
.B(n_204),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_122),
.B(n_156),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_86),
.B(n_121),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_68),
.B(n_85),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_46),
.B(n_67),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_42),
.B(n_45),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_38),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_38),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_35),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_32),
.Y(n_218)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_40),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_48),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_57),
.B2(n_58),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_60),
.C(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_53),
.Y(n_272)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_66),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_84),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_84),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_77),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_76),
.C(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_74),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_77),
.Y(n_389)
);

FAx1_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.CI(n_83),
.CON(n_77),
.SN(n_77)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_106),
.C(n_107),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_81),
.Y(n_365)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_82),
.Y(n_261)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_89),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_104),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_90),
.B(n_105),
.C(n_108),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_93),
.C(n_96),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_94),
.B(n_139),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_103),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_102),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_117),
.C(n_119),
.Y(n_154)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_115),
.Y(n_288)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_116),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_155),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_155),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_135),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_125),
.B(n_134),
.C(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_133),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_131),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_182),
.C(n_183),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_147),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_149),
.C(n_153),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g390 ( 
.A(n_136),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_141),
.CI(n_144),
.CON(n_136),
.SN(n_136)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_141),
.C(n_144),
.Y(n_179)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_140),
.Y(n_236)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_143),
.Y(n_244)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_143),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_143),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_146),
.Y(n_232)
);

INVx6_ASAP7_75t_L g320 ( 
.A(n_146),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_146),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_153),
.B2(n_154),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_202),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_202),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_180),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_160),
.B(n_161),
.C(n_180),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_176),
.B2(n_177),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_162),
.B(n_225),
.C(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_166),
.C(n_175),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_170),
.B2(n_175),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx8_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_172),
.B(n_308),
.Y(n_307)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_185),
.C(n_201),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_190),
.B1(n_200),
.B2(n_201),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_188),
.B(n_189),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_188),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_189),
.B(n_209),
.C(n_220),
.Y(n_279)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_191),
.B(n_196),
.C(n_198),
.Y(n_246)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_196),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_247),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_SL g248 ( 
.A(n_206),
.B(n_247),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_223),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_222),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_208),
.B(n_222),
.C(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_219),
.B2(n_221),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_211),
.B(n_215),
.C(n_290),
.Y(n_289)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_223),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_228),
.C(n_239),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_239),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_234),
.C(n_237),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_246),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_245),
.Y(n_240)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_241),
.B(n_245),
.C(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_246),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_293),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_293),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_251),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_278),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_253),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_263),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_254),
.B(n_264),
.C(n_267),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_255),
.B(n_259),
.C(n_262),
.Y(n_335)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_271),
.C(n_274),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_273),
.B1(n_274),
.B2(n_277),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_271),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_273),
.A2(n_274),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_273),
.B(n_305),
.C(n_307),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_278),
.B(n_337),
.C(n_338),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_283),
.B1(n_291),
.B2(n_292),
.Y(n_280)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_292),
.C(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_287),
.C(n_289),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_336),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_297),
.B(n_336),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_298),
.B(n_386),
.C(n_387),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_321),
.Y(n_300)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_301),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_309),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_302),
.B(n_310),
.C(n_311),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_307),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_304),
.A2(n_305),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_312),
.B(n_317),
.C(n_318),
.Y(n_356)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_324),
.C(n_325),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_335),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_330),
.B1(n_333),
.B2(n_334),
.Y(n_326)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_330),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_333),
.C(n_375),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_330),
.A2(n_334),
.B1(n_379),
.B2(n_383),
.Y(n_378)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_335),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_388),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_385),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_385),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_372),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_355),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_370),
.B2(n_371),
.Y(n_355)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_357),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_362),
.Y(n_357)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx11_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_384),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_379),
.Y(n_383)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx8_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);


endmodule