module fake_jpeg_16040_n_86 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_29),
.A2(n_1),
.B1(n_3),
.B2(n_11),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_32),
.A2(n_13),
.B1(n_16),
.B2(n_19),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_22),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_56),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_70),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_60),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_66),
.C(n_42),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_79),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_57),
.B(n_61),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_55),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_80),
.C(n_63),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g84 ( 
.A(n_83),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_57),
.C(n_62),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_63),
.Y(n_86)
);


endmodule