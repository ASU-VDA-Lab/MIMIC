module fake_aes_2840_n_1355 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_376, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_378, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1355);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_378;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1355;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_533;
wire n_1010;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_688;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_401;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_1275;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_653;
wire n_881;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_600;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g379 ( .A(n_276), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_5), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_245), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_0), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_152), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_370), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_134), .Y(n_385) );
CKINVDCx16_ASAP7_75t_R g386 ( .A(n_163), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_172), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_272), .Y(n_388) );
CKINVDCx14_ASAP7_75t_R g389 ( .A(n_12), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_146), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_355), .Y(n_391) );
NOR2xp67_ASAP7_75t_L g392 ( .A(n_131), .B(n_307), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_261), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_205), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_156), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_371), .Y(n_396) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_227), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_4), .Y(n_398) );
CKINVDCx14_ASAP7_75t_R g399 ( .A(n_296), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_310), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_297), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_200), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_244), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_232), .Y(n_404) );
NOR2xp67_ASAP7_75t_L g405 ( .A(n_334), .B(n_172), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_366), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_364), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g408 ( .A(n_372), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_368), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_14), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g411 ( .A(n_285), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_308), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_134), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_26), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_195), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_279), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_218), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_100), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_234), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_213), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_363), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_260), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_132), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_313), .Y(n_424) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_155), .Y(n_425) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_50), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_135), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_145), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_139), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_349), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_263), .Y(n_431) );
INVxp67_ASAP7_75t_L g432 ( .A(n_286), .Y(n_432) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_229), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_177), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_362), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_155), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_13), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_41), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_122), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_31), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_38), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_37), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_273), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_91), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_115), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_148), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_42), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_314), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_196), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_133), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_5), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_164), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_167), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_75), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g455 ( .A(n_303), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_243), .Y(n_456) );
INVxp33_ASAP7_75t_SL g457 ( .A(n_267), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_228), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_278), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_335), .Y(n_460) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_190), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_361), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_341), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_369), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_233), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_351), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_321), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_192), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_365), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_188), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_338), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_235), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_241), .Y(n_473) );
INVxp33_ASAP7_75t_SL g474 ( .A(n_93), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_6), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_12), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_46), .Y(n_477) );
INVxp33_ASAP7_75t_L g478 ( .A(n_238), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_118), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_348), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_105), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_298), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_322), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_248), .Y(n_484) );
INVx1_ASAP7_75t_SL g485 ( .A(n_7), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_257), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_183), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_270), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_331), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_210), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_113), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_56), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_84), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_208), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_258), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_266), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_123), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_281), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_311), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_211), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_242), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_58), .Y(n_502) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_32), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_280), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_293), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_377), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_189), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g508 ( .A(n_283), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_6), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_187), .Y(n_510) );
BUFx2_ASAP7_75t_SL g511 ( .A(n_151), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_121), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_367), .Y(n_513) );
XNOR2x1_ASAP7_75t_L g514 ( .A(n_48), .B(n_343), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_4), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_46), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_64), .Y(n_517) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_374), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_304), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_299), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_87), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_130), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_264), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_153), .B(n_289), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_166), .Y(n_525) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_115), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_317), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_346), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_262), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_26), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_329), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_125), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_102), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_77), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_290), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_225), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_112), .Y(n_537) );
INVxp33_ASAP7_75t_L g538 ( .A(n_309), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_128), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_325), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_209), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_25), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_120), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_124), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_330), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_324), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_221), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_173), .Y(n_548) );
INVxp33_ASAP7_75t_SL g549 ( .A(n_358), .Y(n_549) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_96), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_48), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_50), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_207), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_33), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_66), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_40), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_93), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_352), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_89), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_85), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_251), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_37), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_57), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_300), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_141), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_295), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_418), .Y(n_567) );
INVx3_ASAP7_75t_L g568 ( .A(n_425), .Y(n_568) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_384), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_418), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_383), .B(n_1), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_487), .B(n_1), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_438), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_533), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_408), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_487), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_384), .Y(n_577) );
AND2x2_ASAP7_75t_SL g578 ( .A(n_480), .B(n_378), .Y(n_578) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_384), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_438), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_475), .Y(n_581) );
BUFx8_ASAP7_75t_L g582 ( .A(n_384), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_433), .Y(n_583) );
OA21x2_ASAP7_75t_L g584 ( .A1(n_406), .A2(n_185), .B(n_184), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_389), .Y(n_585) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_433), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_411), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_455), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_479), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_402), .B(n_2), .Y(n_590) );
BUFx2_ASAP7_75t_L g591 ( .A(n_389), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_508), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_386), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_520), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_479), .B(n_2), .Y(n_595) );
OAI22xp5_ASAP7_75t_SL g596 ( .A1(n_437), .A2(n_8), .B1(n_3), .B2(n_7), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_536), .B(n_3), .Y(n_597) );
BUFx3_ASAP7_75t_L g598 ( .A(n_421), .Y(n_598) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_433), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_562), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_572), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_572), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_572), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_576), .B(n_541), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_591), .B(n_574), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_598), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_572), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_576), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_576), .B(n_478), .Y(n_609) );
INVx3_ASAP7_75t_L g610 ( .A(n_595), .Y(n_610) );
INVx4_ASAP7_75t_SL g611 ( .A(n_598), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_578), .A2(n_439), .B1(n_440), .B2(n_437), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_591), .B(n_497), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_595), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_595), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_569), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_595), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_568), .Y(n_618) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_569), .Y(n_619) );
INVx3_ASAP7_75t_L g620 ( .A(n_568), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_569), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_569), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_568), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_581), .B(n_478), .Y(n_624) );
BUFx2_ASAP7_75t_L g625 ( .A(n_600), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_598), .B(n_538), .Y(n_626) );
AND2x4_ASAP7_75t_L g627 ( .A(n_567), .B(n_497), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_568), .Y(n_628) );
AND2x6_ASAP7_75t_L g629 ( .A(n_590), .B(n_421), .Y(n_629) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_569), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_577), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_567), .B(n_538), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_570), .B(n_537), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_569), .Y(n_634) );
INVx3_ASAP7_75t_L g635 ( .A(n_627), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_613), .B(n_590), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_624), .A2(n_578), .B1(n_587), .B2(n_575), .Y(n_637) );
INVx5_ASAP7_75t_L g638 ( .A(n_629), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_613), .B(n_597), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_626), .B(n_578), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_601), .B(n_379), .Y(n_641) );
BUFx3_ASAP7_75t_L g642 ( .A(n_606), .Y(n_642) );
INVx2_ASAP7_75t_SL g643 ( .A(n_605), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_631), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_625), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_605), .A2(n_592), .B1(n_594), .B2(n_588), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_606), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_601), .B(n_381), .Y(n_648) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_610), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_614), .A2(n_474), .B1(n_573), .B2(n_570), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_602), .B(n_391), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_609), .B(n_597), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_608), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_606), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_632), .B(n_571), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_631), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_632), .B(n_571), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_602), .B(n_394), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_627), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_613), .B(n_396), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_604), .B(n_564), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_614), .A2(n_474), .B1(n_580), .B2(n_573), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_613), .B(n_457), .Y(n_663) );
BUFx2_ASAP7_75t_L g664 ( .A(n_625), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_627), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_633), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_633), .Y(n_667) );
INVx3_ASAP7_75t_L g668 ( .A(n_633), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_612), .A2(n_585), .B1(n_401), .B2(n_412), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_604), .B(n_564), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_603), .A2(n_584), .B(n_449), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_617), .B(n_457), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_617), .Y(n_673) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_610), .Y(n_674) );
INVx2_ASAP7_75t_SL g675 ( .A(n_629), .Y(n_675) );
INVx5_ASAP7_75t_L g676 ( .A(n_629), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_603), .B(n_566), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_612), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_629), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_620), .Y(n_680) );
AO22x1_ASAP7_75t_L g681 ( .A1(n_629), .A2(n_549), .B1(n_382), .B2(n_548), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_607), .B(n_566), .Y(n_682) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_607), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_610), .A2(n_589), .B1(n_580), .B2(n_387), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_610), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_615), .B(n_399), .Y(n_686) );
AND3x2_ASAP7_75t_SL g687 ( .A(n_629), .B(n_514), .C(n_596), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_615), .A2(n_589), .B1(n_395), .B2(n_398), .Y(n_688) );
BUFx10_ASAP7_75t_L g689 ( .A(n_629), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_629), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_629), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_611), .Y(n_692) );
INVx5_ASAP7_75t_L g693 ( .A(n_620), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_611), .B(n_432), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_611), .B(n_400), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_611), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_628), .B(n_582), .Y(n_697) );
AND2x4_ASAP7_75t_L g698 ( .A(n_628), .B(n_396), .Y(n_698) );
AND2x4_ASAP7_75t_L g699 ( .A(n_628), .B(n_401), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_664), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_640), .A2(n_596), .B1(n_514), .B2(n_582), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_652), .B(n_412), .Y(n_702) );
INVx3_ASAP7_75t_L g703 ( .A(n_649), .Y(n_703) );
INVx4_ASAP7_75t_L g704 ( .A(n_649), .Y(n_704) );
OAI21xp33_ASAP7_75t_SL g705 ( .A1(n_655), .A2(n_503), .B(n_426), .Y(n_705) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_674), .Y(n_706) );
INVx1_ASAP7_75t_SL g707 ( .A(n_645), .Y(n_707) );
OAI21x1_ASAP7_75t_L g708 ( .A1(n_671), .A2(n_584), .B(n_616), .Y(n_708) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_674), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_674), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_635), .Y(n_711) );
AOI21x1_ASAP7_75t_L g712 ( .A1(n_681), .A2(n_584), .B(n_618), .Y(n_712) );
OAI21x1_ASAP7_75t_L g713 ( .A1(n_690), .A2(n_584), .B(n_616), .Y(n_713) );
O2A1O1Ixp5_ASAP7_75t_SL g714 ( .A1(n_695), .A2(n_403), .B(n_407), .C(n_404), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_657), .B(n_382), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_636), .A2(n_582), .B1(n_511), .B2(n_439), .Y(n_716) );
AOI222xp33_ASAP7_75t_L g717 ( .A1(n_678), .A2(n_440), .B1(n_542), .B2(n_442), .C1(n_526), .C2(n_593), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_636), .B(n_434), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_685), .A2(n_623), .B(n_618), .Y(n_719) );
OAI22x1_ASAP7_75t_L g720 ( .A1(n_669), .A2(n_551), .B1(n_555), .B2(n_548), .Y(n_720) );
BUFx12f_ASAP7_75t_L g721 ( .A(n_660), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g722 ( .A1(n_660), .A2(n_442), .B1(n_542), .B2(n_522), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_643), .Y(n_723) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_698), .Y(n_724) );
INVxp67_ASAP7_75t_L g725 ( .A(n_639), .Y(n_725) );
NAND2x1p5_ASAP7_75t_L g726 ( .A(n_668), .B(n_537), .Y(n_726) );
O2A1O1Ixp33_ASAP7_75t_L g727 ( .A1(n_639), .A2(n_410), .B(n_413), .C(n_380), .Y(n_727) );
AND2x4_ASAP7_75t_L g728 ( .A(n_659), .B(n_435), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_683), .B(n_551), .Y(n_729) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_698), .Y(n_730) );
INVx5_ASAP7_75t_L g731 ( .A(n_689), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_683), .A2(n_471), .B1(n_495), .B2(n_468), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_646), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_665), .Y(n_734) );
OAI21xp5_ASAP7_75t_L g735 ( .A1(n_673), .A2(n_623), .B(n_524), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_684), .A2(n_546), .B1(n_561), .B2(n_495), .Y(n_736) );
INVx3_ASAP7_75t_L g737 ( .A(n_693), .Y(n_737) );
INVxp67_ASAP7_75t_L g738 ( .A(n_699), .Y(n_738) );
INVx3_ASAP7_75t_L g739 ( .A(n_693), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_666), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_667), .B(n_546), .Y(n_741) );
INVxp67_ASAP7_75t_L g742 ( .A(n_661), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_653), .Y(n_743) );
O2A1O1Ixp33_ASAP7_75t_L g744 ( .A1(n_663), .A2(n_423), .B(n_427), .C(n_414), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_641), .A2(n_461), .B(n_397), .Y(n_745) );
BUFx3_ASAP7_75t_L g746 ( .A(n_693), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_677), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_663), .A2(n_561), .B1(n_555), .B2(n_390), .Y(n_748) );
BUFx2_ASAP7_75t_L g749 ( .A(n_670), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_637), .B(n_385), .Y(n_750) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_642), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_644), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_672), .A2(n_428), .B1(n_436), .B2(n_429), .Y(n_753) );
INVx3_ASAP7_75t_L g754 ( .A(n_693), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_672), .A2(n_509), .B1(n_530), .B2(n_517), .Y(n_755) );
NAND2xp33_ASAP7_75t_L g756 ( .A(n_638), .B(n_388), .Y(n_756) );
BUFx3_ASAP7_75t_L g757 ( .A(n_656), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_684), .A2(n_444), .B1(n_445), .B2(n_441), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_682), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_641), .A2(n_518), .B(n_469), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_648), .Y(n_761) );
BUFx10_ASAP7_75t_L g762 ( .A(n_694), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_648), .Y(n_763) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_650), .A2(n_447), .B1(n_451), .B2(n_450), .C(n_446), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g765 ( .A(n_638), .B(n_393), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_650), .B(n_485), .Y(n_766) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_642), .Y(n_767) );
BUFx2_ASAP7_75t_L g768 ( .A(n_679), .Y(n_768) );
INVx3_ASAP7_75t_L g769 ( .A(n_689), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_688), .A2(n_453), .B1(n_454), .B2(n_452), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_662), .B(n_476), .Y(n_771) );
INVx3_ASAP7_75t_L g772 ( .A(n_692), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_651), .Y(n_773) );
INVxp33_ASAP7_75t_SL g774 ( .A(n_662), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_675), .B(n_539), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_688), .A2(n_481), .B1(n_491), .B2(n_477), .Y(n_776) );
BUFx2_ASAP7_75t_L g777 ( .A(n_638), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_651), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_680), .Y(n_779) );
NAND2x1p5_ASAP7_75t_L g780 ( .A(n_676), .B(n_492), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_647), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_658), .A2(n_502), .B1(n_512), .B2(n_493), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_658), .B(n_515), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_686), .Y(n_784) );
INVx2_ASAP7_75t_SL g785 ( .A(n_676), .Y(n_785) );
BUFx3_ASAP7_75t_L g786 ( .A(n_696), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_654), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_694), .A2(n_521), .B1(n_525), .B2(n_516), .Y(n_788) );
AOI22xp33_ASAP7_75t_SL g789 ( .A1(n_687), .A2(n_534), .B1(n_543), .B2(n_532), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_697), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_691), .B(n_544), .Y(n_791) );
A2O1A1Ixp33_ASAP7_75t_L g792 ( .A1(n_695), .A2(n_554), .B(n_556), .C(n_552), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_687), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_676), .B(n_557), .Y(n_794) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_649), .Y(n_795) );
NAND2x1p5_ASAP7_75t_L g796 ( .A(n_635), .B(n_559), .Y(n_796) );
AO32x1_ASAP7_75t_L g797 ( .A1(n_690), .A2(n_583), .A3(n_577), .B1(n_415), .B2(n_416), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_757), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_707), .B(n_560), .Y(n_799) );
OR2x2_ASAP7_75t_L g800 ( .A(n_732), .B(n_563), .Y(n_800) );
OAI21x1_ASAP7_75t_L g801 ( .A1(n_713), .A2(n_449), .B(n_406), .Y(n_801) );
OR2x2_ASAP7_75t_L g802 ( .A(n_732), .B(n_565), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_774), .B(n_494), .Y(n_803) );
INVx1_ASAP7_75t_SL g804 ( .A(n_707), .Y(n_804) );
AO21x2_ASAP7_75t_L g805 ( .A1(n_712), .A2(n_405), .B(n_392), .Y(n_805) );
OAI21x1_ASAP7_75t_L g806 ( .A1(n_708), .A2(n_463), .B(n_462), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_752), .Y(n_807) );
INVx8_ASAP7_75t_L g808 ( .A(n_721), .Y(n_808) );
OAI21x1_ASAP7_75t_L g809 ( .A1(n_714), .A2(n_501), .B(n_472), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_700), .Y(n_810) );
INVx4_ASAP7_75t_L g811 ( .A(n_706), .Y(n_811) );
OAI21x1_ASAP7_75t_L g812 ( .A1(n_772), .A2(n_510), .B(n_507), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g813 ( .A1(n_784), .A2(n_510), .B(n_507), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_725), .A2(n_736), .B1(n_793), .B2(n_743), .Y(n_814) );
OA21x2_ASAP7_75t_L g815 ( .A1(n_791), .A2(n_545), .B(n_531), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_796), .Y(n_816) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_736), .Y(n_817) );
OAI21x1_ASAP7_75t_L g818 ( .A1(n_772), .A2(n_545), .B(n_531), .Y(n_818) );
O2A1O1Ixp33_ASAP7_75t_SL g819 ( .A1(n_791), .A2(n_417), .B(n_420), .C(n_419), .Y(n_819) );
OAI21x1_ASAP7_75t_L g820 ( .A1(n_780), .A2(n_424), .B(n_422), .Y(n_820) );
AO32x2_ASAP7_75t_L g821 ( .A1(n_758), .A2(n_579), .A3(n_599), .B1(n_586), .B2(n_550), .Y(n_821) );
OAI21x1_ASAP7_75t_L g822 ( .A1(n_780), .A2(n_431), .B(n_430), .Y(n_822) );
NOR2x1_ASAP7_75t_R g823 ( .A(n_728), .B(n_409), .Y(n_823) );
OAI21x1_ASAP7_75t_L g824 ( .A1(n_719), .A2(n_448), .B(n_443), .Y(n_824) );
AOI222xp33_ASAP7_75t_L g825 ( .A1(n_701), .A2(n_425), .B1(n_550), .B2(n_456), .C1(n_460), .C2(n_459), .Y(n_825) );
XOR2xp5_ASAP7_75t_L g826 ( .A(n_722), .B(n_8), .Y(n_826) );
OAI21xp5_ASAP7_75t_L g827 ( .A1(n_790), .A2(n_464), .B(n_458), .Y(n_827) );
OAI21x1_ASAP7_75t_SL g828 ( .A1(n_704), .A2(n_466), .B(n_465), .Y(n_828) );
O2A1O1Ixp33_ASAP7_75t_L g829 ( .A1(n_744), .A2(n_467), .B(n_473), .C(n_470), .Y(n_829) );
NAND2xp33_ASAP7_75t_SL g830 ( .A(n_751), .B(n_425), .Y(n_830) );
OA21x2_ASAP7_75t_L g831 ( .A1(n_735), .A2(n_484), .B(n_482), .Y(n_831) );
OAI21x1_ASAP7_75t_L g832 ( .A1(n_719), .A2(n_489), .B(n_488), .Y(n_832) );
BUFx2_ASAP7_75t_L g833 ( .A(n_741), .Y(n_833) );
OAI21x1_ASAP7_75t_L g834 ( .A1(n_726), .A2(n_496), .B(n_490), .Y(n_834) );
BUFx3_ASAP7_75t_L g835 ( .A(n_746), .Y(n_835) );
OAI21x1_ASAP7_75t_L g836 ( .A1(n_726), .A2(n_500), .B(n_498), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_742), .B(n_504), .Y(n_837) );
INVx3_ASAP7_75t_L g838 ( .A(n_751), .Y(n_838) );
INVxp67_ASAP7_75t_L g839 ( .A(n_723), .Y(n_839) );
AO32x2_ASAP7_75t_L g840 ( .A1(n_758), .A2(n_599), .A3(n_586), .B1(n_579), .B2(n_577), .Y(n_840) );
OAI21x1_ASAP7_75t_L g841 ( .A1(n_703), .A2(n_506), .B(n_505), .Y(n_841) );
OAI21x1_ASAP7_75t_L g842 ( .A1(n_703), .A2(n_519), .B(n_513), .Y(n_842) );
OAI21x1_ASAP7_75t_L g843 ( .A1(n_794), .A2(n_527), .B(n_523), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_747), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_759), .Y(n_845) );
OAI21x1_ASAP7_75t_L g846 ( .A1(n_794), .A2(n_540), .B(n_528), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_789), .A2(n_547), .B1(n_558), .B2(n_553), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_715), .B(n_483), .Y(n_848) );
INVx4_ASAP7_75t_SL g849 ( .A(n_767), .Y(n_849) );
INVx6_ASAP7_75t_L g850 ( .A(n_706), .Y(n_850) );
AO31x2_ASAP7_75t_L g851 ( .A1(n_792), .A2(n_583), .A3(n_622), .B(n_621), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_715), .A2(n_535), .B1(n_433), .B2(n_583), .Y(n_852) );
NAND2xp33_ASAP7_75t_L g853 ( .A(n_767), .B(n_486), .Y(n_853) );
OR2x6_ASAP7_75t_L g854 ( .A(n_738), .B(n_535), .Y(n_854) );
NAND2x1p5_ASAP7_75t_L g855 ( .A(n_706), .B(n_535), .Y(n_855) );
OR2x2_ASAP7_75t_L g856 ( .A(n_702), .B(n_9), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_734), .Y(n_857) );
AO21x2_ASAP7_75t_L g858 ( .A1(n_735), .A2(n_622), .B(n_621), .Y(n_858) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_724), .Y(n_859) );
AO21x2_ASAP7_75t_L g860 ( .A1(n_761), .A2(n_634), .B(n_622), .Y(n_860) );
INVx6_ASAP7_75t_L g861 ( .A(n_709), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_749), .B(n_9), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_748), .B(n_10), .Y(n_863) );
INVx3_ASAP7_75t_L g864 ( .A(n_737), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_740), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_729), .Y(n_866) );
BUFx6f_ASAP7_75t_L g867 ( .A(n_709), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_718), .B(n_499), .Y(n_868) );
BUFx10_ASAP7_75t_L g869 ( .A(n_730), .Y(n_869) );
O2A1O1Ixp33_ASAP7_75t_L g870 ( .A1(n_727), .A2(n_634), .B(n_13), .C(n_10), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_783), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_770), .A2(n_529), .B1(n_586), .B2(n_579), .Y(n_872) );
BUFx3_ASAP7_75t_L g873 ( .A(n_739), .Y(n_873) );
INVx4_ASAP7_75t_L g874 ( .A(n_709), .Y(n_874) );
AND2x4_ASAP7_75t_L g875 ( .A(n_711), .B(n_11), .Y(n_875) );
AO21x2_ASAP7_75t_L g876 ( .A1(n_763), .A2(n_586), .B(n_579), .Y(n_876) );
BUFx2_ASAP7_75t_L g877 ( .A(n_705), .Y(n_877) );
AO21x1_ASAP7_75t_L g878 ( .A1(n_773), .A2(n_599), .B(n_579), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_783), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_733), .Y(n_880) );
INVxp67_ASAP7_75t_SL g881 ( .A(n_710), .Y(n_881) );
OR2x2_ASAP7_75t_L g882 ( .A(n_718), .B(n_14), .Y(n_882) );
OAI21x1_ASAP7_75t_L g883 ( .A1(n_754), .A2(n_599), .B(n_191), .Y(n_883) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_797), .A2(n_630), .B(n_619), .Y(n_884) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_710), .Y(n_885) );
OAI21x1_ASAP7_75t_SL g886 ( .A1(n_778), .A2(n_15), .B(n_16), .Y(n_886) );
AO31x2_ASAP7_75t_L g887 ( .A1(n_771), .A2(n_599), .A3(n_630), .B(n_619), .Y(n_887) );
NAND3xp33_ASAP7_75t_L g888 ( .A(n_753), .B(n_599), .C(n_619), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_771), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_766), .A2(n_630), .B1(n_619), .B2(n_17), .Y(n_890) );
OR2x2_ASAP7_75t_L g891 ( .A(n_720), .B(n_15), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_764), .B(n_16), .Y(n_892) );
NAND3xp33_ASAP7_75t_SL g893 ( .A(n_717), .B(n_17), .C(n_18), .Y(n_893) );
OAI21x1_ASAP7_75t_L g894 ( .A1(n_754), .A2(n_193), .B(n_186), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_781), .Y(n_895) );
NOR3xp33_ASAP7_75t_L g896 ( .A(n_750), .B(n_18), .C(n_19), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_764), .B(n_19), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_782), .Y(n_898) );
OAI21x1_ASAP7_75t_L g899 ( .A1(n_769), .A2(n_197), .B(n_194), .Y(n_899) );
OAI21x1_ASAP7_75t_L g900 ( .A1(n_769), .A2(n_199), .B(n_198), .Y(n_900) );
OAI21x1_ASAP7_75t_L g901 ( .A1(n_787), .A2(n_202), .B(n_201), .Y(n_901) );
O2A1O1Ixp33_ASAP7_75t_L g902 ( .A1(n_716), .A2(n_22), .B(n_20), .C(n_21), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g903 ( .A1(n_776), .A2(n_22), .B1(n_20), .B2(n_21), .Y(n_903) );
AO31x2_ASAP7_75t_L g904 ( .A1(n_797), .A2(n_619), .A3(n_630), .B(n_25), .Y(n_904) );
OAI21x1_ASAP7_75t_L g905 ( .A1(n_765), .A2(n_204), .B(n_203), .Y(n_905) );
OAI21x1_ASAP7_75t_L g906 ( .A1(n_779), .A2(n_760), .B(n_745), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_788), .Y(n_907) );
CKINVDCx8_ASAP7_75t_R g908 ( .A(n_777), .Y(n_908) );
OAI21x1_ASAP7_75t_L g909 ( .A1(n_775), .A2(n_212), .B(n_206), .Y(n_909) );
OA21x2_ASAP7_75t_L g910 ( .A1(n_797), .A2(n_768), .B(n_785), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_762), .A2(n_630), .B1(n_619), .B2(n_27), .Y(n_911) );
BUFx3_ASAP7_75t_L g912 ( .A(n_786), .Y(n_912) );
AND2x4_ASAP7_75t_L g913 ( .A(n_731), .B(n_23), .Y(n_913) );
AND2x4_ASAP7_75t_L g914 ( .A(n_731), .B(n_23), .Y(n_914) );
AOI22xp33_ASAP7_75t_SL g915 ( .A1(n_814), .A2(n_717), .B1(n_795), .B2(n_710), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_889), .B(n_795), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_844), .Y(n_917) );
A2O1A1Ixp33_ASAP7_75t_L g918 ( .A1(n_902), .A2(n_755), .B(n_756), .C(n_795), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g919 ( .A(n_896), .B(n_630), .C(n_731), .Y(n_919) );
OAI22xp33_ASAP7_75t_L g920 ( .A1(n_817), .A2(n_28), .B1(n_24), .B2(n_27), .Y(n_920) );
AOI21xp5_ASAP7_75t_L g921 ( .A1(n_806), .A2(n_215), .B(n_214), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_845), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_814), .A2(n_30), .B1(n_28), .B2(n_29), .C(n_31), .Y(n_923) );
AOI22xp33_ASAP7_75t_SL g924 ( .A1(n_817), .A2(n_36), .B1(n_34), .B2(n_35), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_857), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_893), .A2(n_36), .B1(n_34), .B2(n_35), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_903), .A2(n_40), .B1(n_38), .B2(n_39), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_893), .A2(n_42), .B1(n_39), .B2(n_41), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_803), .A2(n_45), .B1(n_43), .B2(n_44), .Y(n_929) );
OAI221xp5_ASAP7_75t_L g930 ( .A1(n_803), .A2(n_45), .B1(n_43), .B2(n_44), .C(n_47), .Y(n_930) );
OAI21xp33_ASAP7_75t_L g931 ( .A1(n_837), .A2(n_47), .B(n_49), .Y(n_931) );
INVx2_ASAP7_75t_SL g932 ( .A(n_808), .Y(n_932) );
AND2x4_ASAP7_75t_L g933 ( .A(n_816), .B(n_51), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_903), .A2(n_54), .B1(n_52), .B2(n_53), .Y(n_934) );
AOI221xp5_ASAP7_75t_L g935 ( .A1(n_866), .A2(n_55), .B1(n_53), .B2(n_54), .C(n_56), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_804), .Y(n_936) );
AO21x2_ASAP7_75t_L g937 ( .A1(n_805), .A2(n_217), .B(n_216), .Y(n_937) );
OAI21xp5_ASAP7_75t_L g938 ( .A1(n_813), .A2(n_59), .B(n_60), .Y(n_938) );
OAI211xp5_ASAP7_75t_L g939 ( .A1(n_825), .A2(n_826), .B(n_896), .C(n_847), .Y(n_939) );
AOI221xp5_ASAP7_75t_L g940 ( .A1(n_907), .A2(n_63), .B1(n_61), .B2(n_62), .C(n_64), .Y(n_940) );
INVx3_ASAP7_75t_L g941 ( .A(n_811), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_799), .B(n_62), .Y(n_942) );
A2O1A1Ixp33_ASAP7_75t_SL g943 ( .A1(n_837), .A2(n_66), .B(n_63), .C(n_65), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_833), .A2(n_68), .B1(n_65), .B2(n_67), .Y(n_944) );
AOI21xp33_ASAP7_75t_L g945 ( .A1(n_870), .A2(n_67), .B(n_68), .Y(n_945) );
AOI21xp5_ASAP7_75t_L g946 ( .A1(n_801), .A2(n_220), .B(n_219), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g947 ( .A1(n_829), .A2(n_71), .B1(n_69), .B2(n_70), .C(n_72), .Y(n_947) );
OR2x2_ASAP7_75t_L g948 ( .A(n_800), .B(n_69), .Y(n_948) );
AOI221xp5_ASAP7_75t_L g949 ( .A1(n_829), .A2(n_72), .B1(n_70), .B2(n_71), .C(n_73), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_807), .Y(n_950) );
AOI21xp5_ASAP7_75t_L g951 ( .A1(n_858), .A2(n_223), .B(n_222), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_854), .A2(n_75), .B1(n_73), .B2(n_74), .Y(n_952) );
NAND2x1p5_ASAP7_75t_L g953 ( .A(n_913), .B(n_74), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_877), .A2(n_79), .B1(n_76), .B2(n_78), .Y(n_954) );
INVx3_ASAP7_75t_L g955 ( .A(n_811), .Y(n_955) );
AO31x2_ASAP7_75t_L g956 ( .A1(n_878), .A2(n_81), .A3(n_79), .B(n_80), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_863), .A2(n_82), .B1(n_80), .B2(n_81), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_898), .A2(n_84), .B1(n_82), .B2(n_83), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_865), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_875), .Y(n_960) );
AND2x4_ASAP7_75t_L g961 ( .A(n_849), .B(n_912), .Y(n_961) );
NOR2x1_ASAP7_75t_SL g962 ( .A(n_854), .B(n_83), .Y(n_962) );
OAI221xp5_ASAP7_75t_L g963 ( .A1(n_802), .A2(n_87), .B1(n_85), .B2(n_86), .C(n_88), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g964 ( .A1(n_810), .A2(n_92), .B1(n_90), .B2(n_91), .Y(n_964) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_808), .Y(n_965) );
INVx3_ASAP7_75t_L g966 ( .A(n_874), .Y(n_966) );
AND2x2_ASAP7_75t_L g967 ( .A(n_862), .B(n_92), .Y(n_967) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_854), .A2(n_96), .B1(n_94), .B2(n_95), .Y(n_968) );
AOI221xp5_ASAP7_75t_L g969 ( .A1(n_892), .A2(n_94), .B1(n_95), .B2(n_97), .C(n_98), .Y(n_969) );
OAI21xp5_ASAP7_75t_L g970 ( .A1(n_813), .A2(n_99), .B(n_100), .Y(n_970) );
AOI22xp5_ASAP7_75t_L g971 ( .A1(n_880), .A2(n_103), .B1(n_101), .B2(n_102), .Y(n_971) );
OAI221xp5_ASAP7_75t_L g972 ( .A1(n_839), .A2(n_103), .B1(n_104), .B2(n_105), .C(n_106), .Y(n_972) );
INVxp33_ASAP7_75t_L g973 ( .A(n_823), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_890), .A2(n_107), .B1(n_104), .B2(n_106), .Y(n_974) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_880), .A2(n_109), .B1(n_107), .B2(n_108), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_859), .B(n_110), .Y(n_976) );
AOI21xp5_ASAP7_75t_L g977 ( .A1(n_858), .A2(n_226), .B(n_224), .Y(n_977) );
CKINVDCx5p33_ASAP7_75t_R g978 ( .A(n_808), .Y(n_978) );
AOI21x1_ASAP7_75t_L g979 ( .A1(n_884), .A2(n_231), .B(n_230), .Y(n_979) );
OAI22xp33_ASAP7_75t_L g980 ( .A1(n_892), .A2(n_114), .B1(n_111), .B2(n_113), .Y(n_980) );
INVx2_ASAP7_75t_L g981 ( .A(n_895), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_897), .B(n_114), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_856), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_891), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_882), .Y(n_985) );
OAI221xp5_ASAP7_75t_L g986 ( .A1(n_827), .A2(n_116), .B1(n_117), .B2(n_119), .C(n_120), .Y(n_986) );
NOR2xp33_ASAP7_75t_L g987 ( .A(n_848), .B(n_122), .Y(n_987) );
AOI21xp33_ASAP7_75t_L g988 ( .A1(n_805), .A2(n_123), .B(n_124), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_913), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_871), .B(n_125), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_879), .A2(n_128), .B1(n_126), .B2(n_127), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_914), .Y(n_992) );
AO22x2_ASAP7_75t_L g993 ( .A1(n_828), .A2(n_131), .B1(n_129), .B2(n_130), .Y(n_993) );
AND2x4_ASAP7_75t_L g994 ( .A(n_849), .B(n_132), .Y(n_994) );
OAI221xp5_ASAP7_75t_SL g995 ( .A1(n_890), .A2(n_133), .B1(n_135), .B2(n_136), .C(n_137), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_868), .A2(n_141), .B1(n_138), .B2(n_140), .Y(n_996) );
AOI21xp5_ASAP7_75t_L g997 ( .A1(n_881), .A2(n_237), .B(n_236), .Y(n_997) );
INVx8_ASAP7_75t_L g998 ( .A(n_867), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_868), .A2(n_798), .B1(n_869), .B2(n_872), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_911), .A2(n_144), .B1(n_142), .B2(n_143), .Y(n_1000) );
INVx2_ASAP7_75t_L g1001 ( .A(n_906), .Y(n_1001) );
OAI221xp5_ASAP7_75t_L g1002 ( .A1(n_911), .A2(n_142), .B1(n_143), .B2(n_144), .C(n_145), .Y(n_1002) );
OAI221xp5_ASAP7_75t_L g1003 ( .A1(n_852), .A2(n_146), .B1(n_147), .B2(n_148), .C(n_149), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_835), .B(n_147), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_886), .Y(n_1005) );
OAI22xp33_ASAP7_75t_L g1006 ( .A1(n_908), .A2(n_149), .B1(n_150), .B2(n_151), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_873), .B(n_153), .Y(n_1007) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_819), .A2(n_154), .B1(n_156), .B2(n_157), .C(n_158), .Y(n_1008) );
INVx2_ASAP7_75t_SL g1009 ( .A(n_864), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_834), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_836), .Y(n_1011) );
AND2x4_ASAP7_75t_L g1012 ( .A(n_849), .B(n_154), .Y(n_1012) );
INVx3_ASAP7_75t_L g1013 ( .A(n_874), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_819), .Y(n_1014) );
OAI21xp5_ASAP7_75t_L g1015 ( .A1(n_824), .A2(n_832), .B(n_888), .Y(n_1015) );
BUFx3_ASAP7_75t_L g1016 ( .A(n_838), .Y(n_1016) );
INVx2_ASAP7_75t_L g1017 ( .A(n_815), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_831), .B(n_159), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_831), .B(n_160), .Y(n_1019) );
AOI221xp5_ASAP7_75t_L g1020 ( .A1(n_888), .A2(n_161), .B1(n_162), .B2(n_163), .C(n_164), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_864), .Y(n_1021) );
OAI211xp5_ASAP7_75t_L g1022 ( .A1(n_830), .A2(n_161), .B(n_162), .C(n_165), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_910), .A2(n_165), .B1(n_166), .B2(n_167), .Y(n_1023) );
A2O1A1Ixp33_ASAP7_75t_L g1024 ( .A1(n_843), .A2(n_168), .B(n_169), .C(n_170), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_851), .Y(n_1025) );
NAND2x1_ASAP7_75t_L g1026 ( .A(n_1017), .B(n_1010), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_925), .B(n_821), .Y(n_1027) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_976), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_950), .B(n_904), .Y(n_1029) );
INVx2_ASAP7_75t_SL g1030 ( .A(n_998), .Y(n_1030) );
BUFx3_ASAP7_75t_L g1031 ( .A(n_965), .Y(n_1031) );
INVx3_ASAP7_75t_L g1032 ( .A(n_998), .Y(n_1032) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1001), .Y(n_1033) );
BUFx3_ASAP7_75t_L g1034 ( .A(n_961), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_917), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_922), .Y(n_1036) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_941), .B(n_838), .Y(n_1037) );
HB1xp67_ASAP7_75t_L g1038 ( .A(n_936), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_959), .Y(n_1039) );
OR2x2_ASAP7_75t_L g1040 ( .A(n_984), .B(n_887), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_981), .B(n_840), .Y(n_1041) );
INVx2_ASAP7_75t_L g1042 ( .A(n_916), .Y(n_1042) );
AND2x4_ASAP7_75t_L g1043 ( .A(n_941), .B(n_867), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1044 ( .A(n_955), .B(n_867), .Y(n_1044) );
AND2x4_ASAP7_75t_L g1045 ( .A(n_955), .B(n_885), .Y(n_1045) );
NOR2x1_ASAP7_75t_SL g1046 ( .A(n_952), .B(n_885), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_982), .B(n_840), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_915), .B(n_840), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_939), .B(n_853), .Y(n_1049) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_948), .B(n_910), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_933), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_1018), .B(n_851), .Y(n_1052) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_1011), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1019), .B(n_851), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_985), .B(n_809), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_938), .B(n_812), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_938), .B(n_818), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_1025), .Y(n_1058) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_990), .B(n_846), .Y(n_1059) );
NOR2xp67_ASAP7_75t_L g1060 ( .A(n_978), .B(n_171), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_983), .B(n_820), .Y(n_1061) );
INVx3_ASAP7_75t_L g1062 ( .A(n_966), .Y(n_1062) );
BUFx2_ASAP7_75t_L g1063 ( .A(n_953), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_970), .B(n_860), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_970), .B(n_860), .Y(n_1065) );
BUFx2_ASAP7_75t_L g1066 ( .A(n_953), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_942), .B(n_822), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_993), .B(n_885), .Y(n_1068) );
INVx3_ASAP7_75t_L g1069 ( .A(n_966), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_956), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_987), .B(n_841), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_967), .B(n_842), .Y(n_1072) );
NOR3xp33_ASAP7_75t_L g1073 ( .A(n_930), .B(n_830), .C(n_909), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1004), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1007), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_960), .Y(n_1076) );
INVx2_ASAP7_75t_L g1077 ( .A(n_979), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_961), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_927), .B(n_894), .Y(n_1079) );
AND2x2_ASAP7_75t_SL g1080 ( .A(n_994), .B(n_899), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_927), .B(n_934), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_952), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_937), .Y(n_1083) );
INVx2_ASAP7_75t_SL g1084 ( .A(n_932), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_968), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_994), .B(n_850), .Y(n_1086) );
BUFx6f_ASAP7_75t_L g1087 ( .A(n_1013), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1012), .B(n_861), .Y(n_1088) );
AND2x4_ASAP7_75t_L g1089 ( .A(n_989), .B(n_900), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_968), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_992), .B(n_876), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_986), .Y(n_1092) );
INVx2_ASAP7_75t_L g1093 ( .A(n_937), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_986), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_923), .B(n_861), .Y(n_1095) );
INVx2_ASAP7_75t_L g1096 ( .A(n_1014), .Y(n_1096) );
INVxp67_ASAP7_75t_SL g1097 ( .A(n_962), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1021), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_924), .B(n_855), .Y(n_1099) );
OR2x2_ASAP7_75t_L g1100 ( .A(n_1005), .B(n_174), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1016), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_926), .B(n_883), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_980), .Y(n_1103) );
BUFx3_ASAP7_75t_L g1104 ( .A(n_1009), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_928), .B(n_901), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_974), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_969), .B(n_174), .Y(n_1107) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_1000), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_945), .B(n_175), .Y(n_1109) );
BUFx3_ASAP7_75t_L g1110 ( .A(n_919), .Y(n_1110) );
INVx2_ASAP7_75t_L g1111 ( .A(n_1015), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_957), .B(n_176), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_999), .A2(n_905), .B1(n_177), .B2(n_178), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_963), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_920), .Y(n_1115) );
INVx2_ASAP7_75t_L g1116 ( .A(n_1015), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_931), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_919), .Y(n_1118) );
BUFx6f_ASAP7_75t_L g1119 ( .A(n_921), .Y(n_1119) );
NOR2xp33_ASAP7_75t_L g1120 ( .A(n_973), .B(n_178), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_954), .B(n_179), .Y(n_1121) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1002), .Y(n_1122) );
INVx2_ASAP7_75t_L g1123 ( .A(n_1003), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_929), .B(n_179), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1008), .B(n_180), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_991), .B(n_180), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_972), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_971), .Y(n_1128) );
OR2x2_ASAP7_75t_L g1129 ( .A(n_995), .B(n_181), .Y(n_1129) );
BUFx2_ASAP7_75t_L g1130 ( .A(n_918), .Y(n_1130) );
INVx2_ASAP7_75t_L g1131 ( .A(n_975), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1023), .B(n_181), .Y(n_1132) );
AO21x2_ASAP7_75t_L g1133 ( .A1(n_988), .A2(n_182), .B(n_239), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_988), .B(n_240), .Y(n_1134) );
BUFx3_ASAP7_75t_L g1135 ( .A(n_1022), .Y(n_1135) );
AND2x4_ASAP7_75t_L g1136 ( .A(n_1034), .B(n_1024), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_1081), .A2(n_947), .B1(n_949), .B2(n_1006), .Y(n_1137) );
NAND3xp33_ASAP7_75t_L g1138 ( .A(n_1049), .B(n_1020), .C(n_940), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1074), .B(n_964), .Y(n_1139) );
NAND2xp5_ASAP7_75t_SL g1140 ( .A(n_1063), .B(n_935), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1028), .B(n_944), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1035), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1036), .Y(n_1143) );
AND2x4_ASAP7_75t_L g1144 ( .A(n_1034), .B(n_958), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1075), .B(n_996), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1039), .Y(n_1146) );
AOI211xp5_ASAP7_75t_L g1147 ( .A1(n_1066), .A2(n_943), .B(n_977), .C(n_951), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1038), .B(n_997), .Y(n_1148) );
CKINVDCx5p33_ASAP7_75t_R g1149 ( .A(n_1031), .Y(n_1149) );
OAI33xp33_ASAP7_75t_L g1150 ( .A1(n_1129), .A2(n_246), .A3(n_247), .B1(n_249), .B2(n_250), .B3(n_252), .Y(n_1150) );
AND2x6_ASAP7_75t_SL g1151 ( .A(n_1120), .B(n_253), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1040), .Y(n_1152) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_1108), .A2(n_946), .B1(n_255), .B2(n_256), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1084), .B(n_254), .Y(n_1154) );
NAND2xp5_ASAP7_75t_SL g1155 ( .A(n_1087), .B(n_259), .Y(n_1155) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1042), .Y(n_1156) );
INVx5_ASAP7_75t_L g1157 ( .A(n_1087), .Y(n_1157) );
NAND5xp2_ASAP7_75t_L g1158 ( .A(n_1073), .B(n_265), .C(n_268), .D(n_269), .E(n_271), .Y(n_1158) );
OAI22xp5_ASAP7_75t_L g1159 ( .A1(n_1129), .A2(n_274), .B1(n_275), .B2(n_277), .Y(n_1159) );
INVx2_ASAP7_75t_SL g1160 ( .A(n_1031), .Y(n_1160) );
NOR2xp33_ASAP7_75t_SL g1161 ( .A(n_1080), .B(n_1079), .Y(n_1161) );
AND2x4_ASAP7_75t_L g1162 ( .A(n_1062), .B(n_282), .Y(n_1162) );
INVx5_ASAP7_75t_L g1163 ( .A(n_1032), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1040), .Y(n_1164) );
INVx5_ASAP7_75t_L g1165 ( .A(n_1032), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1104), .B(n_284), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1076), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1128), .B(n_287), .Y(n_1168) );
INVx5_ASAP7_75t_L g1169 ( .A(n_1043), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1101), .B(n_288), .Y(n_1170) );
BUFx6f_ASAP7_75t_L g1171 ( .A(n_1030), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1098), .Y(n_1172) );
OR2x6_ASAP7_75t_L g1173 ( .A(n_1068), .B(n_291), .Y(n_1173) );
AND2x4_ASAP7_75t_L g1174 ( .A(n_1062), .B(n_292), .Y(n_1174) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1058), .Y(n_1175) );
OAI322xp33_ASAP7_75t_SL g1176 ( .A1(n_1082), .A2(n_1085), .A3(n_1090), .B1(n_1094), .B2(n_1092), .C1(n_1114), .C2(n_1127), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1058), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1178 ( .A1(n_1115), .A2(n_1103), .B1(n_1106), .B2(n_1107), .C(n_1131), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1067), .B(n_294), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1067), .B(n_301), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1100), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1078), .B(n_302), .Y(n_1182) );
INVx4_ASAP7_75t_L g1183 ( .A(n_1069), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1050), .B(n_376), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1051), .Y(n_1185) );
OAI211xp5_ASAP7_75t_L g1186 ( .A1(n_1060), .A2(n_305), .B(n_306), .C(n_312), .Y(n_1186) );
OAI21xp5_ASAP7_75t_L g1187 ( .A1(n_1122), .A2(n_375), .B(n_316), .Y(n_1187) );
OAI221xp5_ASAP7_75t_L g1188 ( .A1(n_1122), .A2(n_315), .B1(n_318), .B2(n_319), .C(n_320), .Y(n_1188) );
AND2x4_ASAP7_75t_L g1189 ( .A(n_1069), .B(n_323), .Y(n_1189) );
AO21x2_ASAP7_75t_L g1190 ( .A1(n_1077), .A2(n_326), .B(n_327), .Y(n_1190) );
INVxp67_ASAP7_75t_SL g1191 ( .A(n_1053), .Y(n_1191) );
AND2x4_ASAP7_75t_L g1192 ( .A(n_1069), .B(n_328), .Y(n_1192) );
BUFx2_ASAP7_75t_L g1193 ( .A(n_1043), .Y(n_1193) );
HB1xp67_ASAP7_75t_L g1194 ( .A(n_1026), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1050), .Y(n_1195) );
AOI21xp5_ASAP7_75t_L g1196 ( .A1(n_1080), .A2(n_332), .B(n_333), .Y(n_1196) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1029), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1072), .B(n_336), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1061), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1059), .B(n_373), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1112), .B(n_337), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1052), .B(n_1054), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1052), .B(n_339), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1121), .B(n_340), .Y(n_1204) );
HB1xp67_ASAP7_75t_L g1205 ( .A(n_1026), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1047), .B(n_1064), .Y(n_1206) );
AO21x2_ASAP7_75t_L g1207 ( .A1(n_1077), .A2(n_342), .B(n_344), .Y(n_1207) );
AOI221xp5_ASAP7_75t_L g1208 ( .A1(n_1125), .A2(n_345), .B1(n_347), .B2(n_350), .C(n_353), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1109), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1121), .B(n_354), .Y(n_1210) );
NOR2xp33_ASAP7_75t_L g1211 ( .A(n_1139), .B(n_1135), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1212 ( .A(n_1202), .B(n_1091), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1195), .B(n_1064), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1142), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1143), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1152), .B(n_1065), .Y(n_1216) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1172), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1146), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1164), .B(n_1065), .Y(n_1219) );
NOR2xp33_ASAP7_75t_L g1220 ( .A(n_1140), .B(n_1135), .Y(n_1220) );
NAND5xp2_ASAP7_75t_SL g1221 ( .A(n_1149), .B(n_1125), .C(n_1048), .D(n_1132), .E(n_1126), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1167), .Y(n_1222) );
HB1xp67_ASAP7_75t_L g1223 ( .A(n_1191), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1209), .B(n_1055), .Y(n_1224) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1175), .Y(n_1225) );
AND2x4_ASAP7_75t_L g1226 ( .A(n_1191), .B(n_1046), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1185), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1193), .B(n_1046), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1179), .B(n_1047), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1178), .B(n_1070), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1180), .B(n_1079), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1178), .B(n_1070), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1199), .B(n_1130), .Y(n_1233) );
AND2x4_ASAP7_75t_L g1234 ( .A(n_1169), .B(n_1110), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1181), .B(n_1088), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1177), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1156), .B(n_1086), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1169), .B(n_1045), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1206), .B(n_1111), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1169), .B(n_1044), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1206), .B(n_1111), .Y(n_1241) );
AND2x4_ASAP7_75t_L g1242 ( .A(n_1173), .B(n_1097), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1197), .Y(n_1243) );
HB1xp67_ASAP7_75t_L g1244 ( .A(n_1194), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1145), .B(n_1116), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1184), .Y(n_1246) );
HB1xp67_ASAP7_75t_L g1247 ( .A(n_1205), .Y(n_1247) );
INVx2_ASAP7_75t_L g1248 ( .A(n_1183), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1141), .B(n_1116), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1160), .B(n_1037), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1148), .B(n_1117), .Y(n_1251) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_1205), .Y(n_1252) );
NOR2xp33_ASAP7_75t_L g1253 ( .A(n_1151), .B(n_1123), .Y(n_1253) );
NAND2x1p5_ASAP7_75t_L g1254 ( .A(n_1163), .B(n_1099), .Y(n_1254) );
INVxp67_ASAP7_75t_L g1255 ( .A(n_1200), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1136), .B(n_1118), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1136), .B(n_1118), .Y(n_1257) );
OR2x6_ASAP7_75t_L g1258 ( .A(n_1196), .B(n_1089), .Y(n_1258) );
AND2x4_ASAP7_75t_L g1259 ( .A(n_1157), .B(n_1089), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1171), .B(n_1027), .Y(n_1260) );
NAND2x1_ASAP7_75t_L g1261 ( .A(n_1162), .B(n_1089), .Y(n_1261) );
NOR2xp33_ASAP7_75t_L g1262 ( .A(n_1144), .B(n_1095), .Y(n_1262) );
AND2x4_ASAP7_75t_L g1263 ( .A(n_1163), .B(n_1096), .Y(n_1263) );
NOR3xp33_ASAP7_75t_L g1264 ( .A(n_1158), .B(n_1124), .C(n_1071), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1203), .B(n_1056), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1137), .B(n_1057), .Y(n_1266) );
OAI322xp33_ASAP7_75t_L g1267 ( .A1(n_1161), .A2(n_1113), .A3(n_1095), .B1(n_1096), .B2(n_1093), .C1(n_1083), .C2(n_1134), .Y(n_1267) );
OAI21xp33_ASAP7_75t_L g1268 ( .A1(n_1158), .A2(n_1134), .B(n_1105), .Y(n_1268) );
NAND2xp33_ASAP7_75t_SL g1269 ( .A(n_1261), .B(n_1159), .Y(n_1269) );
NOR2xp33_ASAP7_75t_L g1270 ( .A(n_1220), .B(n_1138), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1271 ( .A(n_1212), .B(n_1033), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1214), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1262), .B(n_1057), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1224), .B(n_1093), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1215), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1231), .B(n_1041), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1218), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1243), .B(n_1176), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1222), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1229), .B(n_1260), .Y(n_1280) );
NOR3xp33_ASAP7_75t_L g1281 ( .A(n_1253), .B(n_1208), .C(n_1186), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1249), .B(n_1198), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1249), .B(n_1166), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1216), .B(n_1162), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1266), .B(n_1176), .Y(n_1285) );
HB1xp67_ASAP7_75t_L g1286 ( .A(n_1223), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1265), .B(n_1102), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1235), .B(n_1163), .Y(n_1288) );
NOR2xp33_ASAP7_75t_L g1289 ( .A(n_1211), .B(n_1168), .Y(n_1289) );
INVx2_ASAP7_75t_L g1290 ( .A(n_1217), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_1216), .B(n_1174), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1250), .B(n_1163), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1227), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1245), .B(n_1201), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1295 ( .A(n_1219), .B(n_1189), .Y(n_1295) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1225), .Y(n_1296) );
INVx2_ASAP7_75t_L g1297 ( .A(n_1236), .Y(n_1297) );
HB1xp67_ASAP7_75t_L g1298 ( .A(n_1223), .Y(n_1298) );
NAND2x1p5_ASAP7_75t_L g1299 ( .A(n_1242), .B(n_1165), .Y(n_1299) );
INVxp67_ASAP7_75t_SL g1300 ( .A(n_1244), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1213), .B(n_1174), .Y(n_1301) );
AOI22xp5_ASAP7_75t_L g1302 ( .A1(n_1270), .A2(n_1264), .B1(n_1268), .B2(n_1242), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1280), .B(n_1228), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1272), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1275), .Y(n_1305) );
OAI322xp33_ASAP7_75t_L g1306 ( .A1(n_1285), .A2(n_1255), .A3(n_1233), .B1(n_1251), .B2(n_1256), .C1(n_1257), .C2(n_1232), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1277), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1279), .Y(n_1308) );
OAI322xp33_ASAP7_75t_L g1309 ( .A1(n_1278), .A2(n_1233), .A3(n_1256), .B1(n_1257), .B2(n_1230), .C1(n_1232), .C2(n_1213), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1297), .B(n_1286), .Y(n_1310) );
INVx2_ASAP7_75t_L g1311 ( .A(n_1298), .Y(n_1311) );
OAI32xp33_ASAP7_75t_L g1312 ( .A1(n_1269), .A2(n_1254), .A3(n_1248), .B1(n_1247), .B2(n_1252), .Y(n_1312) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_1281), .A2(n_1221), .B1(n_1258), .B2(n_1246), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1276), .B(n_1226), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1276), .B(n_1259), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1297), .B(n_1293), .Y(n_1316) );
AOI21xp5_ASAP7_75t_L g1317 ( .A1(n_1299), .A2(n_1150), .B(n_1267), .Y(n_1317) );
AOI22xp5_ASAP7_75t_L g1318 ( .A1(n_1289), .A2(n_1237), .B1(n_1239), .B2(n_1241), .Y(n_1318) );
XNOR2x1_ASAP7_75t_L g1319 ( .A(n_1302), .B(n_1282), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1316), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1310), .Y(n_1321) );
INVx2_ASAP7_75t_L g1322 ( .A(n_1311), .Y(n_1322) );
NAND2x1p5_ASAP7_75t_L g1323 ( .A(n_1317), .B(n_1234), .Y(n_1323) );
INVx2_ASAP7_75t_L g1324 ( .A(n_1304), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1305), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1318), .B(n_1287), .Y(n_1326) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1307), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1308), .Y(n_1328) );
OAI221xp5_ASAP7_75t_L g1329 ( .A1(n_1313), .A2(n_1294), .B1(n_1300), .B2(n_1273), .C(n_1284), .Y(n_1329) );
OAI32xp33_ASAP7_75t_L g1330 ( .A1(n_1315), .A2(n_1301), .A3(n_1295), .B1(n_1291), .B2(n_1283), .Y(n_1330) );
AOI22xp33_ASAP7_75t_SL g1331 ( .A1(n_1323), .A2(n_1312), .B1(n_1288), .B2(n_1292), .Y(n_1331) );
AOI31xp33_ASAP7_75t_L g1332 ( .A1(n_1323), .A2(n_1150), .A3(n_1314), .B(n_1303), .Y(n_1332) );
NOR2xp33_ASAP7_75t_L g1333 ( .A(n_1319), .B(n_1309), .Y(n_1333) );
O2A1O1Ixp33_ASAP7_75t_L g1334 ( .A1(n_1329), .A2(n_1306), .B(n_1188), .C(n_1153), .Y(n_1334) );
OAI22xp5_ASAP7_75t_L g1335 ( .A1(n_1319), .A2(n_1271), .B1(n_1296), .B2(n_1290), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1321), .B(n_1274), .Y(n_1336) );
OAI21xp5_ASAP7_75t_SL g1337 ( .A1(n_1326), .A2(n_1210), .B(n_1204), .Y(n_1337) );
NAND4xp25_ASAP7_75t_L g1338 ( .A(n_1333), .B(n_1147), .C(n_1330), .D(n_1187), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1336), .Y(n_1339) );
OAI21xp5_ASAP7_75t_SL g1340 ( .A1(n_1332), .A2(n_1328), .B(n_1327), .Y(n_1340) );
OAI22xp5_ASAP7_75t_L g1341 ( .A1(n_1331), .A2(n_1320), .B1(n_1325), .B2(n_1324), .Y(n_1341) );
A2O1A1Ixp33_ASAP7_75t_L g1342 ( .A1(n_1331), .A2(n_1322), .B(n_1240), .C(n_1238), .Y(n_1342) );
AOI211xp5_ASAP7_75t_SL g1343 ( .A1(n_1335), .A2(n_1153), .B(n_1154), .C(n_1182), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1339), .Y(n_1344) );
AOI21xp33_ASAP7_75t_SL g1345 ( .A1(n_1340), .A2(n_1334), .B(n_1337), .Y(n_1345) );
NOR2x1_ASAP7_75t_L g1346 ( .A(n_1341), .B(n_1192), .Y(n_1346) );
OR4x2_ASAP7_75t_L g1347 ( .A(n_1345), .B(n_1342), .C(n_1338), .D(n_1343), .Y(n_1347) );
NOR3xp33_ASAP7_75t_L g1348 ( .A(n_1346), .B(n_1155), .C(n_1170), .Y(n_1348) );
NOR3xp33_ASAP7_75t_SL g1349 ( .A(n_1344), .B(n_1133), .C(n_357), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1347), .Y(n_1350) );
AOI22xp5_ASAP7_75t_L g1351 ( .A1(n_1350), .A2(n_1349), .B1(n_1348), .B2(n_1263), .Y(n_1351) );
BUFx3_ASAP7_75t_L g1352 ( .A(n_1351), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_1352), .A2(n_1119), .B1(n_1207), .B2(n_1190), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1353), .Y(n_1354) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_1354), .A2(n_356), .B1(n_359), .B2(n_360), .Y(n_1355) );
endmodule