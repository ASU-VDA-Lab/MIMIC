module fake_netlist_5_953_n_1954 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_389, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_397, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_400, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_395, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_402, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_66, n_177, n_60, n_403, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_409, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_391, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1954);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_389;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_400;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_402;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_403;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_391;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1954;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1360;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1728;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_1948;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_550;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_464;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_1538;
wire n_1162;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_512;
wire n_1591;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_824;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_815;
wire n_1795;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_1437;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_507;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_1457;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_1937;
wire n_585;
wire n_1739;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_437;
wire n_1642;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_289),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_43),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_16),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_55),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_88),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_132),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_177),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_312),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_284),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_15),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_410),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_329),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_393),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_70),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_202),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_84),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_407),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_230),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_378),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_330),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_45),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_98),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_152),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_309),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_332),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_386),
.Y(n_438)
);

BUFx10_ASAP7_75t_L g439 ( 
.A(n_217),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_240),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_272),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_256),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_38),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_165),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_362),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_53),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_279),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_367),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_233),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_262),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_57),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_201),
.Y(n_452)
);

BUFx10_ASAP7_75t_L g453 ( 
.A(n_108),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_155),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_142),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_96),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_363),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_302),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_228),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_214),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_13),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_134),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_186),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_133),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_189),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_328),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_184),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_131),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_86),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_168),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_151),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_377),
.Y(n_474)
);

BUFx8_ASAP7_75t_SL g475 ( 
.A(n_15),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_120),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_71),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_28),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_31),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_394),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_169),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_344),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_396),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_296),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_10),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_3),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_327),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_382),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_263),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_65),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_297),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_318),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_255),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_275),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_3),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_379),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_107),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_325),
.Y(n_498)
);

INVxp33_ASAP7_75t_L g499 ( 
.A(n_308),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_79),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_31),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_10),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_102),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_23),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_269),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_234),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_203),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_49),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_323),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_209),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_178),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_361),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_167),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_399),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_42),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_128),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_298),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_374),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_226),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_163),
.Y(n_520)
);

BUFx2_ASAP7_75t_SL g521 ( 
.A(n_95),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_171),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_101),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_277),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_220),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_317),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_409),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_114),
.Y(n_528)
);

BUFx8_ASAP7_75t_SL g529 ( 
.A(n_337),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_221),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_345),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_391),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_41),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_360),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_395),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_260),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_343),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_231),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_349),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_405),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_257),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_144),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_352),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_138),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_406),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_271),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_370),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_58),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_310),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_143),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_404),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_156),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_303),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_38),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_339),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_375),
.Y(n_556)
);

INVxp33_ASAP7_75t_R g557 ( 
.A(n_194),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_77),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_331),
.Y(n_559)
);

BUFx10_ASAP7_75t_L g560 ( 
.A(n_173),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_12),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_195),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_290),
.Y(n_563)
);

BUFx5_ASAP7_75t_L g564 ( 
.A(n_99),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_56),
.Y(n_565)
);

BUFx10_ASAP7_75t_L g566 ( 
.A(n_253),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_12),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_389),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_187),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_29),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_9),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_40),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_261),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_398),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_113),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_222),
.Y(n_576)
);

BUFx10_ASAP7_75t_L g577 ( 
.A(n_9),
.Y(n_577)
);

CKINVDCx14_ASAP7_75t_R g578 ( 
.A(n_23),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_381),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_164),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_376),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_11),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_273),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_354),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_250),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_118),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_20),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_47),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_304),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_238),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_229),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_91),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_51),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_254),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_176),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_116),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_316),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_150),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_196),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_44),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_294),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_180),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_388),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_129),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_73),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_350),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_11),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_369),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_258),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_123),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_39),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_353),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_25),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_244),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_110),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_14),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_59),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_32),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_39),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_46),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_392),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_371),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_124),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_342),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_402),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_66),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_32),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_268),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_291),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_351),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_355),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_280),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_170),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_340),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_115),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_243),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_35),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_242),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_162),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_247),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_341),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_37),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_237),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_174),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_365),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_35),
.Y(n_646)
);

BUFx10_ASAP7_75t_L g647 ( 
.A(n_232),
.Y(n_647)
);

CKINVDCx16_ASAP7_75t_R g648 ( 
.A(n_246),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_125),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_248),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_356),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_364),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_18),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_210),
.Y(n_654)
);

INVx1_ASAP7_75t_SL g655 ( 
.A(n_358),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_181),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_74),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_68),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_218),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_111),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_83),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_18),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_239),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_276),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_182),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_2),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_92),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_5),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_383),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_72),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_282),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_172),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_153),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_366),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_8),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_48),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_274),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_28),
.Y(n_678)
);

INVxp33_ASAP7_75t_R g679 ( 
.A(n_198),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_40),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_20),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_4),
.Y(n_682)
);

CKINVDCx14_ASAP7_75t_R g683 ( 
.A(n_121),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_390),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_105),
.Y(n_685)
);

BUFx8_ASAP7_75t_SL g686 ( 
.A(n_385),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_245),
.Y(n_687)
);

CKINVDCx14_ASAP7_75t_R g688 ( 
.A(n_24),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_285),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_313),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_89),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_387),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_2),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_314),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_213),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_17),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_97),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_249),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_135),
.Y(n_699)
);

BUFx8_ASAP7_75t_SL g700 ( 
.A(n_69),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_300),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_288),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_397),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_306),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_223),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_207),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_348),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_227),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_219),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_336),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_161),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_368),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_30),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_67),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_301),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_200),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_145),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_357),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_158),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_82),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_359),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_384),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_37),
.Y(n_723)
);

BUFx8_ASAP7_75t_SL g724 ( 
.A(n_27),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_251),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_414),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_666),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_723),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_666),
.Y(n_729)
);

CKINVDCx16_ASAP7_75t_R g730 ( 
.A(n_606),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_511),
.Y(n_731)
);

INVxp33_ASAP7_75t_SL g732 ( 
.A(n_413),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_567),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_439),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_439),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_666),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_529),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_682),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_686),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_427),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_700),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_696),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_570),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_587),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_475),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_627),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_724),
.Y(n_747)
);

CKINVDCx16_ASAP7_75t_R g748 ( 
.A(n_640),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_637),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_681),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_433),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_693),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_713),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_411),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_437),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_416),
.Y(n_756)
);

CKINVDCx16_ASAP7_75t_R g757 ( 
.A(n_648),
.Y(n_757)
);

INVxp33_ASAP7_75t_L g758 ( 
.A(n_653),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_412),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_415),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_419),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_425),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_564),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_426),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_417),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_577),
.Y(n_766)
);

CKINVDCx16_ASAP7_75t_R g767 ( 
.A(n_578),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_430),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_432),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_577),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_449),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_494),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_441),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_420),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_447),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_564),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_454),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_514),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_458),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_443),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_564),
.Y(n_781)
);

INVxp33_ASAP7_75t_L g782 ( 
.A(n_537),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_418),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_421),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_461),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_422),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_532),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_466),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_618),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_469),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_472),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_473),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_482),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_484),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_423),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_489),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_428),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_429),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_493),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_434),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_453),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_462),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_662),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_565),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_505),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_506),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_435),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_478),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_513),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_720),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_438),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_564),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_516),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_440),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_517),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_442),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_520),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_527),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_533),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_444),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_585),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_445),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_431),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_535),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_536),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_544),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_546),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_551),
.Y(n_828)
);

INVxp33_ASAP7_75t_L g829 ( 
.A(n_424),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_556),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_479),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_446),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_448),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_568),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_451),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_575),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_601),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_576),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_452),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_431),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_580),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_455),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_597),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_605),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_459),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_620),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_626),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_464),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_628),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_468),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_631),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_688),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_471),
.Y(n_853)
);

INVxp67_ASAP7_75t_SL g854 ( 
.A(n_470),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_485),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_632),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_474),
.Y(n_857)
);

INVxp67_ASAP7_75t_SL g858 ( 
.A(n_593),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_476),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_645),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_649),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_650),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_608),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_629),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_657),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_659),
.Y(n_866)
);

INVxp67_ASAP7_75t_SL g867 ( 
.A(n_634),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_669),
.Y(n_868)
);

CKINVDCx16_ASAP7_75t_R g869 ( 
.A(n_683),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_453),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_677),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_684),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_685),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_486),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_689),
.Y(n_875)
);

BUFx10_ASAP7_75t_L g876 ( 
.A(n_495),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_692),
.Y(n_877)
);

CKINVDCx16_ASAP7_75t_R g878 ( 
.A(n_635),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_651),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_480),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_695),
.Y(n_881)
);

INVxp67_ASAP7_75t_SL g882 ( 
.A(n_530),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_481),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_697),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_698),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_703),
.Y(n_886)
);

CKINVDCx16_ASAP7_75t_R g887 ( 
.A(n_694),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_483),
.Y(n_888)
);

INVxp33_ASAP7_75t_L g889 ( 
.A(n_499),
.Y(n_889)
);

CKINVDCx14_ASAP7_75t_R g890 ( 
.A(n_490),
.Y(n_890)
);

INVxp67_ASAP7_75t_SL g891 ( 
.A(n_542),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_715),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_488),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_711),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_501),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_712),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_714),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_594),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_431),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_717),
.Y(n_900)
);

INVxp33_ASAP7_75t_SL g901 ( 
.A(n_502),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_504),
.Y(n_902)
);

INVxp33_ASAP7_75t_SL g903 ( 
.A(n_554),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_603),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_436),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_490),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_491),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_496),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_497),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_467),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_561),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_498),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_564),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_487),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_508),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_510),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_509),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_523),
.Y(n_918)
);

INVxp67_ASAP7_75t_SL g919 ( 
.A(n_460),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_573),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_512),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_571),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_515),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_589),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_518),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_600),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_667),
.Y(n_927)
);

CKINVDCx16_ASAP7_75t_R g928 ( 
.A(n_522),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_522),
.Y(n_929)
);

CKINVDCx16_ASAP7_75t_R g930 ( 
.A(n_540),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_710),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_457),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_540),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_457),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_564),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_519),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_457),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_492),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_572),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_525),
.Y(n_940)
);

BUFx2_ASAP7_75t_SL g941 ( 
.A(n_560),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_526),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_492),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_492),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_531),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_639),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_507),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_534),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_538),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_507),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_507),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_528),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_582),
.Y(n_953)
);

CKINVDCx16_ASAP7_75t_R g954 ( 
.A(n_560),
.Y(n_954)
);

INVxp33_ASAP7_75t_L g955 ( 
.A(n_528),
.Y(n_955)
);

BUFx10_ASAP7_75t_L g956 ( 
.A(n_607),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_528),
.Y(n_957)
);

INVxp67_ASAP7_75t_SL g958 ( 
.A(n_702),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_539),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_541),
.Y(n_960)
);

INVxp33_ASAP7_75t_SL g961 ( 
.A(n_611),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_543),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_549),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_549),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_545),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_547),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_549),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_548),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_599),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_599),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_599),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_664),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_550),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_613),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_552),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_664),
.Y(n_976)
);

CKINVDCx16_ASAP7_75t_R g977 ( 
.A(n_566),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_553),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_664),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_616),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_566),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_596),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_619),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_642),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_558),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_646),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_668),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_675),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_736),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_904),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_889),
.A2(n_680),
.B1(n_678),
.B2(n_456),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_734),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_736),
.Y(n_993)
);

OA21x2_ASAP7_75t_L g994 ( 
.A1(n_759),
.A2(n_761),
.B(n_760),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_823),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_852),
.B(n_477),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_754),
.B(n_450),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_727),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_756),
.B(n_463),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_SL g1000 ( 
.A(n_767),
.B(n_596),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_823),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_882),
.B(n_647),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_840),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_840),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_765),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_823),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_943),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_766),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_899),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_988),
.B(n_500),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_783),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_784),
.B(n_524),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_786),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_943),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_943),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_795),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_797),
.B(n_615),
.Y(n_1017)
);

CKINVDCx8_ASAP7_75t_R g1018 ( 
.A(n_941),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_798),
.B(n_559),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_869),
.B(n_647),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_891),
.B(n_687),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_938),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_947),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_971),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_729),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_735),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_726),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_898),
.B(n_687),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_763),
.A2(n_465),
.B(n_521),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_800),
.B(n_562),
.Y(n_1030)
);

AND2x6_ASAP7_75t_L g1031 ( 
.A(n_776),
.B(n_503),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_899),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_SL g1033 ( 
.A1(n_789),
.A2(n_557),
.B1(n_679),
.B2(n_574),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_980),
.B(n_987),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_807),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_774),
.B(n_555),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_932),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_811),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_934),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_774),
.B(n_579),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_814),
.B(n_563),
.Y(n_1041)
);

INVx6_ASAP7_75t_L g1042 ( 
.A(n_876),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_937),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_801),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_816),
.Y(n_1045)
);

OA21x2_ASAP7_75t_L g1046 ( 
.A1(n_762),
.A2(n_581),
.B(n_569),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_740),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_751),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_944),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_950),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_951),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_820),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_983),
.B(n_590),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_831),
.B(n_612),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_952),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_957),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_984),
.B(n_624),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_876),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_963),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_870),
.B(n_655),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_822),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_832),
.B(n_583),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_738),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_964),
.Y(n_1064)
);

CKINVDCx6p67_ASAP7_75t_R g1065 ( 
.A(n_928),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_906),
.B(n_658),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_755),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_967),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_929),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_833),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_969),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_831),
.B(n_661),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_780),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_970),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_909),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_829),
.A2(n_725),
.B1(n_586),
.B2(n_588),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_972),
.Y(n_1077)
);

NOR2xp67_ASAP7_75t_L g1078 ( 
.A(n_855),
.B(n_584),
.Y(n_1078)
);

AND2x6_ASAP7_75t_L g1079 ( 
.A(n_781),
.B(n_812),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_976),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_979),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_743),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_744),
.Y(n_1083)
);

NAND2x1_ASAP7_75t_L g1084 ( 
.A(n_905),
.B(n_591),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_746),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_749),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_764),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_752),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_768),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_753),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_769),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_913),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_835),
.B(n_722),
.Y(n_1093)
);

BUFx8_ASAP7_75t_L g1094 ( 
.A(n_911),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_935),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_773),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_775),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_933),
.B(n_592),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_910),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_839),
.B(n_721),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_742),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_842),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_917),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_771),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_777),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_914),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_855),
.B(n_595),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_916),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_918),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_772),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_779),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_785),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_920),
.Y(n_1113)
);

INVx5_ASAP7_75t_L g1114 ( 
.A(n_956),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_788),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_874),
.B(n_895),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_782),
.B(n_732),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_R g1118 ( 
.A(n_737),
.B(n_598),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_845),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_790),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_924),
.Y(n_1121)
);

XNOR2x2_ASAP7_75t_R g1122 ( 
.A(n_803),
.B(n_778),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_848),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_874),
.B(n_602),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_926),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_850),
.B(n_719),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_791),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_792),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_793),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_794),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_927),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_796),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_901),
.B(n_903),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_799),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_854),
.B(n_604),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_805),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_806),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_809),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_931),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_813),
.Y(n_1140)
);

OA21x2_ASAP7_75t_L g1141 ( 
.A1(n_815),
.A2(n_610),
.B(n_609),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_817),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_818),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_819),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_858),
.B(n_614),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_824),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_825),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_867),
.B(n_617),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_879),
.B(n_939),
.Y(n_1149)
);

INVxp33_ASAP7_75t_L g1150 ( 
.A(n_802),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_895),
.B(n_621),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_826),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_827),
.Y(n_1153)
);

INVx6_ASAP7_75t_L g1154 ( 
.A(n_956),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_961),
.B(n_622),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_853),
.B(n_718),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_808),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_857),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_828),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_830),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_834),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_836),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_974),
.B(n_623),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_838),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_859),
.B(n_716),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_841),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_787),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_902),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_974),
.B(n_625),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_843),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1006),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1114),
.B(n_730),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1003),
.A2(n_731),
.B1(n_810),
.B2(n_919),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1036),
.B(n_922),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1060),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_990),
.Y(n_1176)
);

AND3x2_ASAP7_75t_L g1177 ( 
.A(n_1000),
.B(n_770),
.C(n_766),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_1079),
.Y(n_1178)
);

OAI21xp33_ASAP7_75t_L g1179 ( 
.A1(n_1040),
.A2(n_758),
.B(n_750),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1022),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1004),
.B(n_880),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1087),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1089),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1005),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1022),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1006),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1114),
.B(n_748),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1091),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1023),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1096),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1023),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1024),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1009),
.B(n_883),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1097),
.Y(n_1194)
);

INVx8_ASAP7_75t_L g1195 ( 
.A(n_1114),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1066),
.B(n_996),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1024),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1018),
.B(n_757),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1039),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1001),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1111),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_989),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1054),
.B(n_888),
.Y(n_1203)
);

AND2x2_ASAP7_75t_SL g1204 ( 
.A(n_1008),
.B(n_878),
.Y(n_1204)
);

NOR2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1065),
.B(n_739),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1032),
.B(n_893),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1007),
.Y(n_1207)
);

NAND2xp33_ASAP7_75t_L g1208 ( 
.A(n_1031),
.B(n_907),
.Y(n_1208)
);

INVxp33_ASAP7_75t_SL g1209 ( 
.A(n_1033),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1112),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1107),
.B(n_908),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1120),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1127),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1128),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1072),
.B(n_953),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1092),
.Y(n_1216)
);

NAND2xp33_ASAP7_75t_L g1217 ( 
.A(n_1031),
.B(n_912),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1039),
.Y(n_1218)
);

INVxp33_ASAP7_75t_L g1219 ( 
.A(n_1117),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1014),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1124),
.B(n_915),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1050),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1015),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_995),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_R g1225 ( 
.A(n_1008),
.B(n_745),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1129),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_995),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1130),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_992),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1132),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1169),
.B(n_923),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1136),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1137),
.Y(n_1233)
);

AND2x2_ASAP7_75t_SL g1234 ( 
.A(n_1133),
.B(n_887),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_993),
.B(n_925),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1138),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1116),
.A2(n_921),
.B1(n_948),
.B2(n_945),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1150),
.B(n_986),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1095),
.Y(n_1239)
);

NOR2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1011),
.B(n_741),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_1042),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1050),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1046),
.A2(n_958),
.B1(n_946),
.B2(n_846),
.Y(n_1243)
);

INVx2_ASAP7_75t_SL g1244 ( 
.A(n_1151),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1071),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_994),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1034),
.B(n_936),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1163),
.Y(n_1248)
);

NOR3xp33_ASAP7_75t_L g1249 ( 
.A(n_1073),
.B(n_954),
.C(n_930),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1071),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1051),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1019),
.B(n_940),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1059),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1149),
.B(n_942),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_994),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1010),
.B(n_959),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1074),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_998),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1144),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1064),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1135),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1140),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1164),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1030),
.B(n_960),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1046),
.A2(n_847),
.B1(n_851),
.B2(n_849),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1170),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1041),
.B(n_965),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1105),
.Y(n_1268)
);

BUFx10_ASAP7_75t_L g1269 ( 
.A(n_1042),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1037),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1145),
.Y(n_1271)
);

AND2x4_ASAP7_75t_SL g1272 ( 
.A(n_1027),
.B(n_804),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1148),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1062),
.B(n_966),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1043),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1064),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1101),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1068),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1101),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1068),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1013),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1105),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1049),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1115),
.Y(n_1284)
);

INVxp67_ASAP7_75t_SL g1285 ( 
.A(n_1115),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1055),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1093),
.B(n_968),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1053),
.A2(n_949),
.B1(n_975),
.B2(n_962),
.Y(n_1288)
);

INVx5_ASAP7_75t_L g1289 ( 
.A(n_1031),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1002),
.Y(n_1290)
);

NOR2xp67_ASAP7_75t_L g1291 ( 
.A(n_1052),
.B(n_973),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1026),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1100),
.B(n_978),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1134),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1146),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1056),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1152),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1153),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1126),
.B(n_985),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1081),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1156),
.B(n_856),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1134),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1099),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_991),
.B(n_986),
.Y(n_1304)
);

NOR3xp33_ASAP7_75t_L g1305 ( 
.A(n_1076),
.B(n_977),
.C(n_770),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1057),
.B(n_981),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1106),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1142),
.Y(n_1308)
);

NAND2xp33_ASAP7_75t_SL g1309 ( 
.A(n_1020),
.B(n_1157),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1058),
.A2(n_982),
.B1(n_750),
.B2(n_733),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_997),
.B(n_890),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1165),
.B(n_860),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1077),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1142),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_999),
.B(n_1012),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1141),
.A2(n_862),
.B1(n_865),
.B2(n_861),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1078),
.B(n_1021),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1108),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1174),
.B(n_1028),
.Y(n_1319)
);

NAND2xp33_ASAP7_75t_SL g1320 ( 
.A(n_1175),
.B(n_1118),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1260),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1176),
.B(n_1075),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1215),
.B(n_1168),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1238),
.B(n_1098),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1196),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1260),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1277),
.B(n_1103),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1289),
.B(n_1016),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1276),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1184),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1259),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1263),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1171),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1315),
.B(n_1155),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1279),
.B(n_1044),
.Y(n_1335)
);

INVx5_ASAP7_75t_L g1336 ( 
.A(n_1241),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1266),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1276),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1219),
.B(n_1035),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1301),
.B(n_1017),
.Y(n_1340)
);

AND2x2_ASAP7_75t_SL g1341 ( 
.A(n_1234),
.B(n_1122),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1278),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1278),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1281),
.Y(n_1344)
);

BUFx4f_ASAP7_75t_L g1345 ( 
.A(n_1195),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1280),
.Y(n_1346)
);

INVxp67_ASAP7_75t_SL g1347 ( 
.A(n_1268),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1171),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_R g1349 ( 
.A(n_1225),
.B(n_1047),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1180),
.B(n_1069),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1181),
.B(n_1038),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1312),
.B(n_1141),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1280),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1216),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1313),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1313),
.Y(n_1356)
);

NAND2x1p5_ASAP7_75t_L g1357 ( 
.A(n_1289),
.B(n_1070),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1289),
.B(n_1290),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1171),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1216),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1229),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1239),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1182),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1252),
.B(n_1045),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1183),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1180),
.B(n_821),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1268),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1189),
.B(n_837),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1239),
.Y(n_1369)
);

INVx4_ASAP7_75t_L g1370 ( 
.A(n_1268),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1292),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1179),
.B(n_1063),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1186),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1193),
.B(n_1061),
.Y(n_1374)
);

OAI221xp5_ASAP7_75t_L g1375 ( 
.A1(n_1243),
.A2(n_872),
.B1(n_873),
.B2(n_875),
.C(n_877),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1306),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1284),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1188),
.Y(n_1378)
);

NAND2x1p5_ASAP7_75t_L g1379 ( 
.A(n_1282),
.B(n_1084),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1303),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1173),
.B(n_1154),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1189),
.B(n_844),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1264),
.B(n_1102),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1206),
.B(n_1119),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1190),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1186),
.Y(n_1386)
);

CKINVDCx8_ASAP7_75t_R g1387 ( 
.A(n_1195),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1203),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1284),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_1241),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1194),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1201),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1304),
.B(n_1123),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1210),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1269),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1211),
.A2(n_1158),
.B1(n_864),
.B2(n_892),
.Y(n_1396)
);

AND2x6_ASAP7_75t_L g1397 ( 
.A(n_1246),
.B(n_866),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1212),
.Y(n_1398)
);

OA22x2_ASAP7_75t_L g1399 ( 
.A1(n_1177),
.A2(n_1237),
.B1(n_1248),
.B2(n_1244),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1242),
.B(n_863),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1267),
.B(n_1079),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1186),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1284),
.Y(n_1403)
);

AO22x2_ASAP7_75t_L g1404 ( 
.A1(n_1288),
.A2(n_728),
.B1(n_733),
.B2(n_868),
.Y(n_1404)
);

NAND2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1294),
.B(n_1084),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1213),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1221),
.B(n_1143),
.Y(n_1407)
);

OAI221xp5_ASAP7_75t_L g1408 ( 
.A1(n_1265),
.A2(n_900),
.B1(n_897),
.B2(n_871),
.C(n_881),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1214),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1274),
.B(n_1287),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1269),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1235),
.B(n_1154),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1226),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1202),
.Y(n_1414)
);

INVx4_ASAP7_75t_L g1415 ( 
.A(n_1294),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1317),
.A2(n_1079),
.B1(n_633),
.B2(n_636),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1185),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1293),
.B(n_1029),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1272),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1261),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1191),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1299),
.B(n_1255),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1240),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1208),
.A2(n_638),
.B1(n_641),
.B2(n_630),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1192),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1228),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1230),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1307),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1232),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1318),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1255),
.B(n_1160),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1197),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1251),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1253),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1321),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_SL g1436 ( 
.A(n_1330),
.B(n_1048),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1334),
.B(n_1231),
.Y(n_1437)
);

NOR2x2_ASAP7_75t_L g1438 ( 
.A(n_1354),
.B(n_1209),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1323),
.B(n_1256),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1411),
.B(n_1271),
.Y(n_1440)
);

NOR2x1_ASAP7_75t_L g1441 ( 
.A(n_1393),
.B(n_1328),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1340),
.B(n_1316),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1319),
.B(n_1204),
.Y(n_1443)
);

AND2x6_ASAP7_75t_L g1444 ( 
.A(n_1422),
.B(n_1410),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1326),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1329),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1360),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1414),
.B(n_1273),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1338),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1362),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1351),
.B(n_1311),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1403),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1352),
.A2(n_1246),
.B1(n_1233),
.B2(n_1236),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1374),
.B(n_1067),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1361),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1384),
.B(n_1342),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1344),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1371),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1339),
.B(n_1104),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1364),
.A2(n_1383),
.B1(n_1399),
.B2(n_1343),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1346),
.A2(n_1262),
.B1(n_1297),
.B2(n_1295),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1353),
.B(n_1291),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1388),
.B(n_1110),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1355),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1341),
.A2(n_1217),
.B1(n_1167),
.B2(n_1247),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1324),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1356),
.B(n_1298),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1369),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1319),
.B(n_1412),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1381),
.B(n_1254),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1327),
.B(n_1314),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1403),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1363),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_SL g1474 ( 
.A(n_1390),
.B(n_1094),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_SL g1475 ( 
.A(n_1322),
.Y(n_1475)
);

INVx5_ASAP7_75t_L g1476 ( 
.A(n_1397),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1372),
.B(n_1285),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1365),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1400),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1372),
.A2(n_1309),
.B1(n_1178),
.B2(n_1310),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1378),
.B(n_1224),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1350),
.Y(n_1482)
);

INVx5_ASAP7_75t_L g1483 ( 
.A(n_1397),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1385),
.B(n_1227),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1391),
.B(n_1270),
.Y(n_1485)
);

OAI21xp33_ASAP7_75t_L g1486 ( 
.A1(n_1325),
.A2(n_1305),
.B(n_1187),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1414),
.B(n_1314),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1331),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1392),
.A2(n_1283),
.B1(n_1286),
.B2(n_1275),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1332),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1394),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1398),
.B(n_1296),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1337),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1336),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1406),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1409),
.B(n_1245),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1336),
.B(n_1198),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1380),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1366),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1333),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1413),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1426),
.B(n_1427),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1428),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1401),
.A2(n_1178),
.B1(n_1300),
.B2(n_1257),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1429),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1368),
.Y(n_1506)
);

AND2x2_ASAP7_75t_SL g1507 ( 
.A(n_1345),
.B(n_1249),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1430),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1396),
.A2(n_747),
.B1(n_728),
.B2(n_1302),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1431),
.B(n_1200),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1433),
.B(n_1207),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1382),
.B(n_1172),
.Y(n_1512)
);

INVx5_ASAP7_75t_L g1513 ( 
.A(n_1397),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1418),
.A2(n_1223),
.B1(n_1220),
.B2(n_1308),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1376),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1455),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1458),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1439),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1443),
.B(n_1404),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1447),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1457),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1437),
.B(n_1420),
.Y(n_1522)
);

AND2x6_ASAP7_75t_L g1523 ( 
.A(n_1435),
.B(n_1335),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_L g1524 ( 
.A(n_1494),
.B(n_1205),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1456),
.B(n_1407),
.Y(n_1525)
);

NAND2x1p5_ASAP7_75t_L g1526 ( 
.A(n_1448),
.B(n_1370),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1515),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1445),
.Y(n_1528)
);

INVx2_ASAP7_75t_SL g1529 ( 
.A(n_1471),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1451),
.B(n_1434),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1500),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1446),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1500),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1479),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1442),
.A2(n_1375),
.B(n_1416),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1460),
.A2(n_1444),
.B1(n_1470),
.B2(n_1469),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1449),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1450),
.Y(n_1538)
);

AO22x1_ASAP7_75t_L g1539 ( 
.A1(n_1454),
.A2(n_1395),
.B1(n_1419),
.B2(n_1423),
.Y(n_1539)
);

BUFx12f_ASAP7_75t_L g1540 ( 
.A(n_1440),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1464),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1473),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1499),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1466),
.B(n_1349),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1444),
.B(n_1347),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1468),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1444),
.B(n_1477),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1480),
.B(n_1320),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1478),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1462),
.B(n_1415),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1438),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1448),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1506),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1482),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1502),
.B(n_1404),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1452),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1496),
.B(n_1417),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1491),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1436),
.B(n_1424),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1488),
.Y(n_1560)
);

INVx4_ASAP7_75t_L g1561 ( 
.A(n_1472),
.Y(n_1561)
);

AOI22x1_ASAP7_75t_L g1562 ( 
.A1(n_1490),
.A2(n_1405),
.B1(n_1379),
.B2(n_1357),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1493),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1453),
.A2(n_1408),
.B1(n_1358),
.B2(n_1377),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1495),
.B(n_1367),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1542),
.Y(n_1566)
);

AOI222xp33_ASAP7_75t_L g1567 ( 
.A1(n_1518),
.A2(n_1459),
.B1(n_1486),
.B2(n_1463),
.C1(n_1509),
.C2(n_1505),
.Y(n_1567)
);

INVxp67_ASAP7_75t_SL g1568 ( 
.A(n_1527),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1522),
.B(n_1465),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1516),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1549),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1528),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1530),
.B(n_1501),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_L g1574 ( 
.A(n_1521),
.B(n_1441),
.Y(n_1574)
);

AND3x1_ASAP7_75t_SL g1575 ( 
.A(n_1558),
.B(n_885),
.C(n_884),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1552),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1525),
.B(n_1467),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1536),
.A2(n_1461),
.B1(n_1483),
.B2(n_1476),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1543),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1533),
.Y(n_1580)
);

NOR2xp67_ASAP7_75t_SL g1581 ( 
.A(n_1540),
.B(n_1387),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1553),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1532),
.Y(n_1583)
);

NOR2x1p5_ASAP7_75t_L g1584 ( 
.A(n_1555),
.B(n_1512),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1537),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1534),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1518),
.B(n_1496),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1554),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1556),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1541),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1536),
.B(n_1485),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1520),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1552),
.Y(n_1593)
);

NAND2x1p5_ASAP7_75t_L g1594 ( 
.A(n_1531),
.B(n_1476),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1519),
.B(n_1492),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1548),
.B(n_1481),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1531),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1517),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1552),
.Y(n_1599)
);

CKINVDCx8_ASAP7_75t_R g1600 ( 
.A(n_1523),
.Y(n_1600)
);

CKINVDCx8_ASAP7_75t_R g1601 ( 
.A(n_1523),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1529),
.Y(n_1602)
);

AND2x6_ASAP7_75t_L g1603 ( 
.A(n_1547),
.B(n_1504),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1595),
.B(n_1570),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1572),
.Y(n_1605)
);

OA21x2_ASAP7_75t_L g1606 ( 
.A1(n_1591),
.A2(n_1547),
.B(n_1535),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1569),
.A2(n_1535),
.B1(n_1559),
.B2(n_1564),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1567),
.A2(n_1507),
.B1(n_1544),
.B2(n_1551),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1566),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1578),
.A2(n_1514),
.B(n_1545),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1572),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_SL g1612 ( 
.A1(n_1596),
.A2(n_1564),
.B(n_1562),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1587),
.B(n_1557),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1584),
.B(n_1557),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1592),
.B(n_1538),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1576),
.B(n_1561),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1582),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1579),
.B(n_1551),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1590),
.A2(n_1510),
.B(n_1550),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1585),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1577),
.B(n_1474),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1573),
.A2(n_1565),
.B1(n_1526),
.B2(n_1497),
.Y(n_1622)
);

AOI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1590),
.A2(n_1484),
.B(n_1511),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1603),
.A2(n_1489),
.B(n_1546),
.Y(n_1624)
);

OR2x6_ASAP7_75t_L g1625 ( 
.A(n_1574),
.B(n_1539),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1571),
.Y(n_1626)
);

OA21x2_ASAP7_75t_L g1627 ( 
.A1(n_1583),
.A2(n_1080),
.B(n_1077),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1568),
.Y(n_1628)
);

OAI21x1_ASAP7_75t_L g1629 ( 
.A1(n_1594),
.A2(n_1563),
.B(n_1560),
.Y(n_1629)
);

AOI22x1_ASAP7_75t_L g1630 ( 
.A1(n_1597),
.A2(n_1561),
.B1(n_1417),
.B2(n_1425),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1586),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1598),
.B(n_1498),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1575),
.A2(n_1523),
.B1(n_1503),
.B2(n_1508),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1603),
.A2(n_1483),
.B(n_1476),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1576),
.Y(n_1635)
);

OAI211xp5_ASAP7_75t_L g1636 ( 
.A1(n_1589),
.A2(n_1524),
.B(n_1487),
.C(n_894),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1603),
.A2(n_1513),
.B(n_1483),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1576),
.Y(n_1638)
);

AO31x2_ASAP7_75t_L g1639 ( 
.A1(n_1603),
.A2(n_896),
.A3(n_886),
.B(n_1250),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_SL g1640 ( 
.A1(n_1600),
.A2(n_1513),
.B(n_1475),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_SL g1641 ( 
.A1(n_1597),
.A2(n_1080),
.B(n_1109),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1593),
.Y(n_1642)
);

O2A1O1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1602),
.A2(n_1085),
.B(n_1086),
.C(n_1082),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1580),
.Y(n_1644)
);

INVx5_ASAP7_75t_L g1645 ( 
.A(n_1593),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1631),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1628),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1605),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1604),
.B(n_1593),
.Y(n_1649)
);

OAI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1607),
.A2(n_1608),
.B(n_1621),
.Y(n_1650)
);

CKINVDCx6p67_ASAP7_75t_R g1651 ( 
.A(n_1645),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1612),
.A2(n_1389),
.B(n_1121),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1625),
.A2(n_1607),
.B1(n_1633),
.B2(n_1617),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1625),
.A2(n_1601),
.B1(n_1588),
.B2(n_1513),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1625),
.A2(n_1599),
.B1(n_1425),
.B2(n_1432),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1609),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1611),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1617),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1633),
.A2(n_1599),
.B1(n_1432),
.B2(n_1421),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1632),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1623),
.A2(n_1125),
.B(n_1113),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1626),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1620),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1618),
.A2(n_1599),
.B1(n_1421),
.B2(n_1348),
.Y(n_1664)
);

INVx4_ASAP7_75t_SL g1665 ( 
.A(n_1614),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1645),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1615),
.B(n_1523),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1622),
.A2(n_1088),
.B1(n_1083),
.B2(n_1162),
.C(n_1090),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1613),
.A2(n_1218),
.B1(n_1222),
.B2(n_1199),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1645),
.B(n_1333),
.Y(n_1670)
);

INVx6_ASAP7_75t_L g1671 ( 
.A(n_1616),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1606),
.B(n_1644),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1624),
.A2(n_1199),
.B1(n_1218),
.B2(n_1222),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1606),
.B(n_1131),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_SL g1675 ( 
.A(n_1636),
.B(n_644),
.C(n_643),
.Y(n_1675)
);

OAI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1624),
.A2(n_1139),
.B1(n_1581),
.B2(n_1083),
.C(n_1088),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1640),
.A2(n_1402),
.B1(n_1386),
.B2(n_1373),
.Y(n_1677)
);

OAI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1643),
.A2(n_1143),
.B1(n_1147),
.B2(n_1159),
.C(n_1161),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1641),
.A2(n_1147),
.B1(n_1159),
.B2(n_1161),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1637),
.A2(n_1359),
.B(n_1348),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1637),
.A2(n_1166),
.B1(n_652),
.B2(n_691),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1635),
.B(n_1359),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1638),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1610),
.A2(n_1166),
.B1(n_654),
.B2(n_699),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1639),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_SL g1686 ( 
.A(n_1634),
.B(n_660),
.C(n_656),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1642),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1649),
.B(n_1639),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1650),
.A2(n_1630),
.B1(n_1616),
.B2(n_1619),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1683),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1654),
.A2(n_1627),
.B1(n_955),
.B2(n_1373),
.Y(n_1691)
);

INVxp33_ASAP7_75t_L g1692 ( 
.A(n_1658),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1653),
.B(n_1629),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1646),
.B(n_1639),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1666),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1662),
.Y(n_1696)
);

CKINVDCx8_ASAP7_75t_R g1697 ( 
.A(n_1665),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1647),
.B(n_1627),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1675),
.A2(n_1676),
.B1(n_1678),
.B2(n_1667),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1672),
.Y(n_1700)
);

NOR3xp33_ASAP7_75t_SL g1701 ( 
.A(n_1655),
.B(n_665),
.C(n_663),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_R g1702 ( 
.A(n_1651),
.B(n_1386),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1648),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1660),
.A2(n_704),
.B1(n_671),
.B2(n_672),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_R g1705 ( 
.A(n_1671),
.B(n_1402),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1687),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1657),
.B(n_1025),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1671),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1663),
.B(n_670),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1656),
.Y(n_1710)
);

INVxp33_ASAP7_75t_L g1711 ( 
.A(n_1682),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1666),
.Y(n_1712)
);

BUFx5_ASAP7_75t_L g1713 ( 
.A(n_1685),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1674),
.Y(n_1714)
);

NAND2xp33_ASAP7_75t_R g1715 ( 
.A(n_1670),
.B(n_0),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1661),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1665),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1652),
.Y(n_1718)
);

AO31x2_ASAP7_75t_L g1719 ( 
.A1(n_1659),
.A2(n_1258),
.A3(n_1),
.B(n_4),
.Y(n_1719)
);

NOR3xp33_ASAP7_75t_SL g1720 ( 
.A(n_1664),
.B(n_674),
.C(n_673),
.Y(n_1720)
);

CKINVDCx6p67_ASAP7_75t_R g1721 ( 
.A(n_1670),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1677),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1686),
.A2(n_709),
.B1(n_708),
.B2(n_707),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1680),
.Y(n_1724)
);

AND2x2_ASAP7_75t_SL g1725 ( 
.A(n_1684),
.B(n_0),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1669),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1668),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1673),
.B(n_1),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1681),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1696),
.Y(n_1730)
);

BUFx2_ASAP7_75t_SL g1731 ( 
.A(n_1717),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1703),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1710),
.Y(n_1733)
);

CKINVDCx14_ASAP7_75t_R g1734 ( 
.A(n_1690),
.Y(n_1734)
);

INVx8_ASAP7_75t_L g1735 ( 
.A(n_1708),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1706),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_5),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1692),
.B(n_1679),
.Y(n_1738)
);

NAND2x1p5_ASAP7_75t_L g1739 ( 
.A(n_1693),
.B(n_50),
.Y(n_1739)
);

INVxp67_ASAP7_75t_SL g1740 ( 
.A(n_1698),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1688),
.B(n_6),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1694),
.B(n_6),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1714),
.B(n_7),
.Y(n_1743)
);

INVx5_ASAP7_75t_L g1744 ( 
.A(n_1708),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1695),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_1695),
.Y(n_1746)
);

NAND2x1_ASAP7_75t_L g1747 ( 
.A(n_1724),
.B(n_1712),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1713),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1711),
.B(n_7),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1708),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1713),
.B(n_8),
.Y(n_1751)
);

INVx2_ASAP7_75t_SL g1752 ( 
.A(n_1705),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1707),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1718),
.B(n_13),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1722),
.B(n_1709),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1713),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1721),
.B(n_14),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1713),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1716),
.B(n_16),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1697),
.B(n_17),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1740),
.B(n_1719),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1740),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1736),
.B(n_1719),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1744),
.B(n_1702),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1746),
.B(n_1719),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1753),
.B(n_1729),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1755),
.A2(n_1725),
.B1(n_1699),
.B2(n_1727),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1746),
.B(n_1689),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1734),
.B(n_1726),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1742),
.B(n_1691),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1738),
.A2(n_1728),
.B1(n_1723),
.B2(n_1704),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1733),
.B(n_1720),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1745),
.B(n_1701),
.Y(n_1773)
);

NOR3xp33_ASAP7_75t_L g1774 ( 
.A(n_1737),
.B(n_1715),
.C(n_690),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1730),
.B(n_19),
.Y(n_1775)
);

AOI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1737),
.A2(n_1743),
.B1(n_1751),
.B2(n_1749),
.C(n_1741),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1731),
.B(n_19),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1739),
.A2(n_1759),
.B1(n_1754),
.B2(n_1760),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1743),
.B(n_21),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_SL g1780 ( 
.A1(n_1739),
.A2(n_706),
.B1(n_705),
.B2(n_701),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1732),
.B(n_21),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1750),
.B(n_22),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1752),
.A2(n_1751),
.B1(n_1744),
.B2(n_1759),
.Y(n_1783)
);

NAND3xp33_ASAP7_75t_L g1784 ( 
.A(n_1754),
.B(n_676),
.C(n_22),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1765),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1763),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1766),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1762),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1768),
.B(n_1750),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1776),
.B(n_1747),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1762),
.B(n_1748),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1783),
.B(n_1744),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1773),
.B(n_1756),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1761),
.B(n_1758),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1764),
.B(n_1757),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1767),
.A2(n_1735),
.B1(n_25),
.B2(n_26),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1782),
.B(n_1735),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1778),
.B(n_1735),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1772),
.B(n_24),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1770),
.B(n_26),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1781),
.B(n_27),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1775),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1779),
.B(n_29),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1777),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1784),
.B(n_1774),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1769),
.B(n_30),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1771),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1785),
.B(n_33),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1791),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1792),
.B(n_1780),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1788),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1793),
.B(n_1780),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1807),
.B(n_33),
.Y(n_1813)
);

OR3x2_ASAP7_75t_L g1814 ( 
.A(n_1805),
.B(n_34),
.C(n_36),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1789),
.B(n_34),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1795),
.B(n_36),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1795),
.B(n_1798),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1787),
.B(n_52),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1786),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1802),
.B(n_54),
.Y(n_1820)
);

NOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1790),
.B(n_1800),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1797),
.B(n_60),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1794),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1794),
.B(n_1801),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1797),
.B(n_61),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1804),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1799),
.B(n_62),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1803),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1803),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1806),
.B(n_63),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1796),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1796),
.B(n_64),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1793),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1793),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1792),
.B(n_75),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1826),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1826),
.Y(n_1837)
);

INVxp67_ASAP7_75t_L g1838 ( 
.A(n_1821),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1813),
.B(n_76),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1824),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1828),
.B(n_78),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1817),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1811),
.Y(n_1843)
);

OA222x2_ASAP7_75t_L g1844 ( 
.A1(n_1831),
.A2(n_80),
.B1(n_81),
.B2(n_85),
.C1(n_87),
.C2(n_90),
.Y(n_1844)
);

INVx4_ASAP7_75t_L g1845 ( 
.A(n_1816),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1829),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1817),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1833),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1808),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1814),
.A2(n_93),
.B1(n_94),
.B2(n_100),
.Y(n_1850)
);

NAND2xp33_ASAP7_75t_SL g1851 ( 
.A(n_1816),
.B(n_103),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1823),
.Y(n_1852)
);

AOI211xp5_ASAP7_75t_L g1853 ( 
.A1(n_1838),
.A2(n_1831),
.B(n_1810),
.C(n_1832),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1839),
.A2(n_1821),
.B(n_1813),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1842),
.Y(n_1855)
);

INVx2_ASAP7_75t_SL g1856 ( 
.A(n_1842),
.Y(n_1856)
);

NOR2xp67_ASAP7_75t_L g1857 ( 
.A(n_1845),
.B(n_1809),
.Y(n_1857)
);

OAI21xp33_ASAP7_75t_L g1858 ( 
.A1(n_1847),
.A2(n_1812),
.B(n_1809),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1845),
.B(n_1835),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1849),
.B(n_1834),
.Y(n_1860)
);

OAI32xp33_ASAP7_75t_L g1861 ( 
.A1(n_1836),
.A2(n_1837),
.A3(n_1840),
.B1(n_1851),
.B2(n_1846),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1848),
.B(n_1835),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1852),
.B(n_1819),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1843),
.B(n_1818),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1841),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1850),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1844),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1863),
.Y(n_1868)
);

A2O1A1Ixp33_ASAP7_75t_L g1869 ( 
.A1(n_1861),
.A2(n_1830),
.B(n_1815),
.C(n_1827),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1860),
.Y(n_1870)
);

AOI21xp33_ASAP7_75t_L g1871 ( 
.A1(n_1861),
.A2(n_1830),
.B(n_1820),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1864),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1867),
.A2(n_1866),
.B1(n_1856),
.B2(n_1859),
.Y(n_1873)
);

OAI221xp5_ASAP7_75t_L g1874 ( 
.A1(n_1853),
.A2(n_1822),
.B1(n_1825),
.B2(n_109),
.C(n_112),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1857),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1858),
.B(n_104),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1870),
.B(n_1862),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_SL g1878 ( 
.A1(n_1874),
.A2(n_1854),
.B1(n_1855),
.B2(n_1865),
.Y(n_1878)
);

NAND2xp33_ASAP7_75t_SL g1879 ( 
.A(n_1875),
.B(n_106),
.Y(n_1879)
);

AOI221x1_ASAP7_75t_SL g1880 ( 
.A1(n_1872),
.A2(n_117),
.B1(n_119),
.B2(n_122),
.C(n_126),
.Y(n_1880)
);

AOI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1873),
.A2(n_127),
.B1(n_130),
.B2(n_136),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1868),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1869),
.Y(n_1883)
);

OAI31xp33_ASAP7_75t_L g1884 ( 
.A1(n_1883),
.A2(n_1871),
.A3(n_1879),
.B(n_1876),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1878),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_1885)
);

OAI21xp5_ASAP7_75t_SL g1886 ( 
.A1(n_1881),
.A2(n_141),
.B(n_146),
.Y(n_1886)
);

O2A1O1Ixp33_ASAP7_75t_L g1887 ( 
.A1(n_1882),
.A2(n_1877),
.B(n_1880),
.C(n_149),
.Y(n_1887)
);

A2O1A1Ixp33_ASAP7_75t_L g1888 ( 
.A1(n_1883),
.A2(n_147),
.B(n_148),
.C(n_154),
.Y(n_1888)
);

AOI211x1_ASAP7_75t_SL g1889 ( 
.A1(n_1885),
.A2(n_157),
.B(n_159),
.C(n_160),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1884),
.B(n_166),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1886),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1891),
.B(n_1887),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1890),
.Y(n_1893)
);

O2A1O1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1892),
.A2(n_1888),
.B(n_1889),
.C(n_183),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1893),
.B(n_175),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1893),
.Y(n_1896)
);

AO22x1_ASAP7_75t_L g1897 ( 
.A1(n_1896),
.A2(n_179),
.B1(n_185),
.B2(n_188),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1895),
.Y(n_1898)
);

OAI322xp33_ASAP7_75t_L g1899 ( 
.A1(n_1898),
.A2(n_1894),
.A3(n_191),
.B1(n_192),
.B2(n_193),
.C1(n_197),
.C2(n_199),
.Y(n_1899)
);

AOI211xp5_ASAP7_75t_SL g1900 ( 
.A1(n_1897),
.A2(n_190),
.B(n_204),
.C(n_205),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1898),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1900),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1901),
.B(n_1899),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1900),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1902),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1904),
.Y(n_1906)
);

NOR3xp33_ASAP7_75t_L g1907 ( 
.A(n_1903),
.B(n_206),
.C(n_208),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1905),
.Y(n_1908)
);

INVx4_ASAP7_75t_L g1909 ( 
.A(n_1906),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1907),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1905),
.Y(n_1911)
);

AOI21xp33_ASAP7_75t_L g1912 ( 
.A1(n_1906),
.A2(n_211),
.B(n_212),
.Y(n_1912)
);

XNOR2x1_ASAP7_75t_L g1913 ( 
.A(n_1908),
.B(n_215),
.Y(n_1913)
);

AOI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1911),
.A2(n_216),
.B(n_224),
.Y(n_1914)
);

XNOR2xp5_ASAP7_75t_L g1915 ( 
.A(n_1910),
.B(n_403),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1909),
.B(n_225),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1912),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1908),
.Y(n_1918)
);

AND3x4_ASAP7_75t_L g1919 ( 
.A(n_1909),
.B(n_235),
.C(n_236),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1908),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1908),
.Y(n_1921)
);

XNOR2xp5_ASAP7_75t_L g1922 ( 
.A(n_1908),
.B(n_401),
.Y(n_1922)
);

CKINVDCx20_ASAP7_75t_R g1923 ( 
.A(n_1909),
.Y(n_1923)
);

XOR2xp5_ASAP7_75t_L g1924 ( 
.A(n_1908),
.B(n_241),
.Y(n_1924)
);

AOI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1920),
.A2(n_252),
.B1(n_259),
.B2(n_264),
.C(n_265),
.Y(n_1925)
);

XNOR2xp5_ASAP7_75t_L g1926 ( 
.A(n_1923),
.B(n_266),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1918),
.B(n_267),
.Y(n_1927)
);

XNOR2xp5_ASAP7_75t_L g1928 ( 
.A(n_1913),
.B(n_270),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1921),
.B(n_278),
.Y(n_1929)
);

NAND2x1p5_ASAP7_75t_L g1930 ( 
.A(n_1916),
.B(n_281),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1917),
.B(n_1914),
.Y(n_1931)
);

NOR2x1p5_ASAP7_75t_L g1932 ( 
.A(n_1919),
.B(n_283),
.Y(n_1932)
);

AO22x2_ASAP7_75t_L g1933 ( 
.A1(n_1924),
.A2(n_286),
.B1(n_287),
.B2(n_292),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1915),
.B(n_293),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1922),
.Y(n_1935)
);

INVx4_ASAP7_75t_L g1936 ( 
.A(n_1918),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1936),
.A2(n_1932),
.B1(n_1931),
.B2(n_1935),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1928),
.A2(n_400),
.B(n_299),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1933),
.Y(n_1939)
);

XOR2xp5_ASAP7_75t_L g1940 ( 
.A(n_1926),
.B(n_295),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1927),
.A2(n_305),
.B1(n_307),
.B2(n_311),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1930),
.B(n_315),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1934),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1942),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1940),
.Y(n_1945)
);

XNOR2xp5_ASAP7_75t_L g1946 ( 
.A(n_1937),
.B(n_1929),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1939),
.Y(n_1947)
);

NOR3xp33_ASAP7_75t_L g1948 ( 
.A(n_1943),
.B(n_1925),
.C(n_320),
.Y(n_1948)
);

AOI222xp33_ASAP7_75t_L g1949 ( 
.A1(n_1947),
.A2(n_1941),
.B1(n_1938),
.B2(n_322),
.C1(n_324),
.C2(n_326),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1944),
.B(n_1946),
.Y(n_1950)
);

AOI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1950),
.A2(n_1948),
.B1(n_1945),
.B2(n_1949),
.Y(n_1951)
);

AOI22x1_ASAP7_75t_L g1952 ( 
.A1(n_1949),
.A2(n_319),
.B1(n_321),
.B2(n_333),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1951),
.A2(n_334),
.B1(n_335),
.B2(n_338),
.Y(n_1953)
);

AOI211xp5_ASAP7_75t_L g1954 ( 
.A1(n_1953),
.A2(n_1952),
.B(n_346),
.C(n_347),
.Y(n_1954)
);


endmodule