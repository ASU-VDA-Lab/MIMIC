module fake_jpeg_10174_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_38),
.B(n_27),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_30),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_72),
.Y(n_85)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_24),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_62),
.B(n_28),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_22),
.B1(n_17),
.B2(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

OA21x2_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_24),
.B(n_28),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_45),
.B1(n_40),
.B2(n_69),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_81),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_40),
.B1(n_45),
.B2(n_20),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_88),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_23),
.B1(n_30),
.B2(n_32),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_30),
.B1(n_27),
.B2(n_31),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_28),
.B1(n_29),
.B2(n_18),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_18),
.B1(n_21),
.B2(n_25),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_87),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_25),
.C(n_34),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_109)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_91),
.Y(n_114)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_67),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_31),
.B1(n_32),
.B2(n_24),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_44),
.C(n_47),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_60),
.C(n_59),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_61),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_101),
.C(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_103),
.B(n_109),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_106),
.A2(n_107),
.B1(n_116),
.B2(n_121),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_50),
.B1(n_49),
.B2(n_57),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_63),
.C(n_66),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_13),
.B(n_12),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_113),
.B(n_115),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_73),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_21),
.B(n_25),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_66),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_124),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_67),
.C(n_47),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_35),
.C(n_46),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_83),
.A2(n_70),
.B1(n_54),
.B2(n_34),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_89),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_21),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_50),
.B1(n_81),
.B2(n_96),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_140),
.B1(n_149),
.B2(n_23),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_124),
.A2(n_75),
.B1(n_74),
.B2(n_97),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_147),
.B1(n_152),
.B2(n_122),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_146),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_85),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_29),
.C(n_110),
.Y(n_169)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_139),
.B(n_141),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_91),
.B1(n_83),
.B2(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_148),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_87),
.B1(n_89),
.B2(n_86),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_150),
.Y(n_182)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_101),
.A2(n_71),
.B1(n_68),
.B2(n_86),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_118),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_156),
.A2(n_115),
.B(n_120),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_157),
.B(n_33),
.Y(n_212)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_111),
.B(n_120),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_160),
.A2(n_167),
.B(n_183),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_111),
.B(n_114),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_179),
.B(n_136),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_150),
.B1(n_23),
.B2(n_19),
.Y(n_199)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_166),
.Y(n_205)
);

OAI221xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_116),
.B1(n_126),
.B2(n_34),
.C(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_105),
.B(n_86),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_105),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_169),
.C(n_170),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_68),
.C(n_110),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_174),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_119),
.B1(n_46),
.B2(n_43),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_173),
.A2(n_130),
.B1(n_154),
.B2(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_172),
.B1(n_174),
.B2(n_138),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_19),
.C(n_26),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_155),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_133),
.B(n_10),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_178),
.B(n_180),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_0),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_133),
.B(n_135),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_19),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_143),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_193),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_198),
.B1(n_207),
.B2(n_158),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_196),
.B1(n_210),
.B2(n_179),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_200),
.C(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_197),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_144),
.B(n_136),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_156),
.B(n_137),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_162),
.A2(n_143),
.B1(n_151),
.B2(n_142),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_199),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_33),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_157),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_19),
.Y(n_203)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_209),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_180),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_208),
.C(n_169),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_173),
.A2(n_23),
.B1(n_26),
.B2(n_33),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_33),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_165),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_0),
.B(n_1),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_179),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_158),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_211),
.A2(n_185),
.B1(n_175),
.B2(n_160),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_207),
.B1(n_213),
.B2(n_210),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_222),
.Y(n_248)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_202),
.B1(n_188),
.B2(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_233),
.B1(n_159),
.B2(n_23),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_227),
.B(n_237),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_177),
.C(n_161),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_232),
.Y(n_254)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_182),
.C(n_181),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_164),
.B1(n_158),
.B2(n_178),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_182),
.C(n_181),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_238),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_208),
.B(n_179),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_165),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_26),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_214),
.A2(n_196),
.B1(n_186),
.B2(n_197),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_235),
.B(n_15),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_197),
.B(n_193),
.Y(n_243)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_243),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_253),
.Y(n_266)
);

XOR2x2_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_190),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_245),
.B(n_225),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_218),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_261),
.B1(n_262),
.B2(n_215),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_219),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_258),
.Y(n_269)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_218),
.A2(n_159),
.B(n_1),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_0),
.B(n_1),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_216),
.A2(n_26),
.B1(n_8),
.B2(n_9),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_220),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_262)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_279),
.Y(n_291)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_232),
.C(n_234),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_268),
.C(n_271),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_223),
.C(n_230),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_277),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_223),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_229),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_224),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_278),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_12),
.B(n_11),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_13),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_240),
.C(n_256),
.Y(n_279)
);

OAI221xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_248),
.B1(n_249),
.B2(n_262),
.C(n_261),
.Y(n_281)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_260),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_290),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_246),
.Y(n_285)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

AOI31xp33_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_242),
.A3(n_250),
.B(n_247),
.Y(n_288)
);

AOI211xp5_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_294),
.B(n_2),
.C(n_3),
.Y(n_308)
);

NOR2x1_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_241),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_285),
.B(n_286),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_252),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_267),
.C(n_268),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_300),
.C(n_302),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_291),
.B(n_279),
.Y(n_298)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_290),
.A2(n_271),
.B(n_270),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_299),
.A2(n_301),
.B(n_310),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_12),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_0),
.C(n_2),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_9),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_294),
.Y(n_313)
);

FAx1_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_2),
.CI(n_3),
.CON(n_306),
.SN(n_306)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_4),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_287),
.B1(n_293),
.B2(n_6),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_2),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_309),
.B(n_284),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_295),
.A2(n_3),
.B(n_4),
.Y(n_310)
);

NAND3xp33_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_283),
.C(n_292),
.Y(n_312)
);

NOR2x1_ASAP7_75t_SL g326 ( 
.A(n_312),
.B(n_306),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_314),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_305),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_318),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_302),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_320),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_297),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_325),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_301),
.Y(n_325)
);

OAI21x1_ASAP7_75t_L g330 ( 
.A1(n_326),
.A2(n_317),
.B(n_5),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_316),
.A2(n_306),
.B(n_309),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_312),
.B(n_4),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_321),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_330),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_4),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_323),
.B(n_322),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_334),
.B(n_331),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_335),
.B(n_333),
.Y(n_337)
);

NAND2x1_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_6),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_7),
.B(n_320),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_7),
.B(n_320),
.Y(n_340)
);


endmodule