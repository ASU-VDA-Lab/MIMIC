module fake_jpeg_9520_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_5),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_4),
.B(n_1),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_10),
.B(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_14),
.Y(n_19)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_15),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_6),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_0),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

OAI21xp33_ASAP7_75t_SL g18 ( 
.A1(n_12),
.A2(n_9),
.B(n_6),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_13),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_24),
.B1(n_25),
.B2(n_18),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_27),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_8),
.B1(n_20),
.B2(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_8),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_30),
.A2(n_8),
.B1(n_24),
.B2(n_27),
.Y(n_31)
);

AOI322xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_29),
.A3(n_7),
.B1(n_8),
.B2(n_4),
.C1(n_3),
.C2(n_2),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_1),
.B1(n_7),
.B2(n_18),
.Y(n_33)
);


endmodule