module fake_jpeg_10905_n_29 (n_3, n_2, n_1, n_0, n_4, n_5, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_R g6 ( 
.A(n_4),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_9),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_0),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_17),
.B1(n_7),
.B2(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx4_ASAP7_75t_SL g16 ( 
.A(n_8),
.Y(n_16)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_6),
.B(n_7),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_15),
.B1(n_10),
.B2(n_17),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_16),
.B(n_20),
.C(n_24),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_8),
.C(n_4),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_18),
.B(n_2),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B(n_16),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_20),
.Y(n_28)
);

HAxp5_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_27),
.CON(n_29),
.SN(n_29)
);


endmodule