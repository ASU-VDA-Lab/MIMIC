module fake_jpeg_4745_n_265 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_43),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_18),
.B1(n_31),
.B2(n_24),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_42),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_58),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_50),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_24),
.B1(n_18),
.B2(n_31),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_52),
.A2(n_32),
.B1(n_14),
.B2(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_21),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_55),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_18),
.B1(n_24),
.B2(n_31),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_61),
.A2(n_78),
.B1(n_50),
.B2(n_52),
.Y(n_108)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_64),
.Y(n_95)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_25),
.B1(n_30),
.B2(n_20),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_76),
.B1(n_82),
.B2(n_1),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_33),
.B(n_19),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_66),
.B(n_81),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_69),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_89),
.Y(n_92)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_70),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_30),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_72),
.Y(n_119)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_77),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_37),
.A2(n_28),
.B1(n_25),
.B2(n_20),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_36),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_39),
.A2(n_28),
.B1(n_19),
.B2(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_36),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_33),
.A2(n_15),
.B1(n_26),
.B2(n_22),
.Y(n_82)
);

CKINVDCx9p33_ASAP7_75t_R g83 ( 
.A(n_35),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_36),
.B(n_22),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_87),
.Y(n_93)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_36),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_32),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_32),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_1),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_110),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_59),
.A2(n_32),
.B1(n_14),
.B2(n_5),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g141 ( 
.A(n_99),
.B(n_111),
.C(n_47),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_14),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_102),
.B(n_116),
.Y(n_136)
);

AO22x2_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_85),
.B1(n_75),
.B2(n_9),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_83),
.Y(n_143)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_59),
.A2(n_63),
.B1(n_62),
.B2(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_82),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_88),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_63),
.B1(n_73),
.B2(n_8),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_57),
.B(n_6),
.Y(n_116)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_71),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_51),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_132),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_128),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_60),
.Y(n_129)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_54),
.C(n_79),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_152),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_60),
.Y(n_131)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_90),
.C(n_68),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_79),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_134),
.B(n_139),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_69),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_137),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_48),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_140),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_118),
.B(n_121),
.C(n_113),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_145),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_147),
.B1(n_116),
.B2(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_107),
.B(n_6),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_74),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_146),
.B(n_150),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_56),
.B1(n_74),
.B2(n_10),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_96),
.A2(n_74),
.B1(n_9),
.B2(n_10),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_148),
.A2(n_151),
.B1(n_105),
.B2(n_102),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_105),
.B(n_7),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_92),
.B(n_93),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_119),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_96),
.A2(n_11),
.B1(n_12),
.B2(n_114),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_93),
.B(n_11),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_166),
.B1(n_169),
.B2(n_171),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_158),
.B(n_159),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_101),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_160),
.A2(n_161),
.B(n_163),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_112),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_94),
.B(n_101),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_142),
.A2(n_118),
.B1(n_104),
.B2(n_120),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_121),
.B1(n_143),
.B2(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_135),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_125),
.A2(n_146),
.B(n_123),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_152),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_138),
.A2(n_143),
.B1(n_149),
.B2(n_130),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_179),
.A2(n_136),
.B1(n_168),
.B2(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_186),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_196),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_133),
.Y(n_182)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_176),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_187),
.C(n_191),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_127),
.Y(n_186)
);

NAND2x1_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_141),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_148),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_188),
.B(n_189),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_139),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_145),
.C(n_151),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_136),
.C(n_179),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_198),
.C(n_173),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_166),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_194),
.B(n_164),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_173),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_160),
.B(n_169),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_155),
.B(n_172),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_163),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_204),
.C(n_198),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_171),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_175),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_212),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_195),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_183),
.A2(n_165),
.B1(n_167),
.B2(n_154),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_191),
.B(n_164),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_195),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_217),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_156),
.B1(n_167),
.B2(n_161),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_187),
.B1(n_167),
.B2(n_161),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_223),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_192),
.C(n_187),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_227),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_196),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_213),
.B(n_211),
.Y(n_238)
);

HAxp5_ASAP7_75t_SL g226 ( 
.A(n_208),
.B(n_180),
.CON(n_226),
.SN(n_226)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_229),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_228),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_172),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_237),
.B(n_238),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_220),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_215),
.B(n_210),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_206),
.B1(n_207),
.B2(n_212),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_233),
.B1(n_239),
.B2(n_235),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_237),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_246),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_235),
.B(n_221),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_243),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_232),
.A2(n_227),
.B1(n_223),
.B2(n_202),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_245),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_234),
.A2(n_220),
.B1(n_226),
.B2(n_229),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_200),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_248),
.A2(n_247),
.B(n_243),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_203),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_216),
.B1(n_201),
.B2(n_231),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_242),
.C(n_224),
.Y(n_257)
);

CKINVDCx12_ASAP7_75t_R g255 ( 
.A(n_249),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_258),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_251),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_170),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_261),
.Y(n_262)
);

AO21x1_ASAP7_75t_L g263 ( 
.A1(n_260),
.A2(n_253),
.B(n_258),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_263),
.A2(n_252),
.B(n_170),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_262),
.Y(n_265)
);


endmodule