module fake_jpeg_2329_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_40),
.Y(n_50)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_48),
.Y(n_59)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_36),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

MAJx2_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_48),
.C(n_38),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_2),
.C(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_38),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_78),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_51),
.B1(n_41),
.B2(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_77),
.Y(n_83)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_45),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_42),
.B(n_37),
.C(n_65),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_6),
.B(n_7),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_86),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_63),
.B1(n_49),
.B2(n_47),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_69),
.B1(n_15),
.B2(n_17),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_49),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_47),
.B(n_3),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_2),
.B(n_4),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_6),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_71),
.B(n_67),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_97),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVxp33_ASAP7_75t_SL g97 ( 
.A(n_84),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_99),
.B(n_83),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_4),
.B(n_5),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_103),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_7),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_8),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_87),
.C(n_81),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_97),
.Y(n_109)
);

OAI322xp33_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_25),
.A3(n_13),
.B1(n_14),
.B2(n_18),
.C1(n_22),
.C2(n_34),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_90),
.B(n_10),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_93),
.B1(n_10),
.B2(n_9),
.Y(n_117)
);

AO22x1_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_24),
.B1(n_33),
.B2(n_11),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_111),
.B1(n_106),
.B2(n_109),
.Y(n_124)
);

AOI321xp33_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_121),
.A3(n_116),
.B1(n_115),
.B2(n_112),
.C(n_32),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_123),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_120),
.B1(n_113),
.B2(n_111),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_125),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_28),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_31),
.C(n_9),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_130),
.Y(n_131)
);


endmodule