module fake_jpeg_28023_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_46),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_24),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_24),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_48),
.Y(n_77)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_64),
.Y(n_92)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_25),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_21),
.B1(n_39),
.B2(n_40),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_69),
.A2(n_76),
.B1(n_97),
.B2(n_62),
.Y(n_119)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_72),
.Y(n_106)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_21),
.B1(n_26),
.B2(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_77),
.B(n_80),
.Y(n_116)
);

BUFx2_ASAP7_75t_SL g78 ( 
.A(n_61),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_82),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

INVxp67_ASAP7_75t_SL g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_87),
.Y(n_110)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_21),
.B1(n_40),
.B2(n_39),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_62),
.B1(n_49),
.B2(n_53),
.Y(n_117)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_46),
.B(n_25),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_91),
.C(n_74),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_47),
.Y(n_91)
);

CKINVDCx12_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_45),
.B1(n_39),
.B2(n_26),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_66),
.B1(n_53),
.B2(n_49),
.Y(n_111)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_57),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_32),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_45),
.B1(n_47),
.B2(n_22),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_102),
.B(n_107),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_37),
.C(n_31),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_91),
.C(n_73),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_57),
.B1(n_62),
.B2(n_49),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_119),
.B1(n_92),
.B2(n_88),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_97),
.B1(n_95),
.B2(n_71),
.Y(n_128)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_37),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_37),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_127),
.Y(n_142)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_143),
.B1(n_108),
.B2(n_112),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_129),
.B(n_22),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_123),
.A2(n_91),
.B(n_85),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_146),
.B(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_133),
.B(n_147),
.Y(n_185)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_94),
.C(n_37),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_127),
.C(n_126),
.Y(n_157)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_44),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_155),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_104),
.B1(n_117),
.B2(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_92),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_145),
.B(n_150),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_SL g146 ( 
.A(n_124),
.B(n_31),
.C(n_22),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

MAJx3_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_44),
.C(n_41),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_44),
.B1(n_41),
.B2(n_38),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_32),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_109),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_44),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_162),
.A2(n_182),
.B1(n_141),
.B2(n_139),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_129),
.B(n_138),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_166),
.B(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_181),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_144),
.A2(n_105),
.B1(n_87),
.B2(n_122),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_165),
.A2(n_174),
.B(n_186),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_112),
.B(n_125),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_168),
.B(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_71),
.B1(n_109),
.B2(n_120),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_36),
.B1(n_33),
.B2(n_30),
.Y(n_209)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_171),
.B(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_179),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_175),
.Y(n_204)
);

OA22x2_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_22),
.B1(n_17),
.B2(n_27),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_125),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_143),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_136),
.A2(n_143),
.B(n_146),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_41),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_135),
.A2(n_29),
.B1(n_34),
.B2(n_33),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_27),
.B(n_34),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_188),
.A2(n_206),
.B(n_207),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_180),
.C(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_201),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_171),
.B(n_29),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_194),
.B(n_196),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_151),
.Y(n_202)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_212),
.B1(n_169),
.B2(n_168),
.Y(n_222)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_1),
.B(n_2),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_141),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_3),
.Y(n_240)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_173),
.A2(n_30),
.B1(n_23),
.B2(n_20),
.Y(n_212)
);

INVx11_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_157),
.B(n_17),
.Y(n_215)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_158),
.B(n_17),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_162),
.A2(n_23),
.B(n_20),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_3),
.B(n_4),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_186),
.C(n_156),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_241),
.C(n_206),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_204),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_221),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_SL g260 ( 
.A(n_222),
.B(n_238),
.C(n_243),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_223),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_156),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_199),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_182),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_166),
.B1(n_4),
.B2(n_5),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_236),
.A2(n_207),
.B1(n_198),
.B2(n_219),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_189),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_245),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_212),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_3),
.C(n_5),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_6),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_205),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_202),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_246),
.B(n_241),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_214),
.B1(n_218),
.B2(n_200),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_262),
.B1(n_240),
.B2(n_251),
.Y(n_268)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_254),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_210),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_215),
.C(n_200),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_228),
.C(n_226),
.Y(n_267)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_198),
.B(n_191),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_195),
.B(n_240),
.Y(n_276)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_191),
.B1(n_192),
.B2(n_201),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_265),
.B1(n_213),
.B2(n_210),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_193),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_266),
.B(n_197),
.Y(n_270)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_269),
.C(n_271),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_273),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_244),
.C(n_227),
.Y(n_269)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_244),
.C(n_227),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_234),
.C(n_224),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_280),
.C(n_277),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_260),
.B1(n_249),
.B2(n_251),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_257),
.A2(n_224),
.B(n_197),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_248),
.B(n_265),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_259),
.B(n_258),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_284),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_236),
.C(n_238),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_210),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_194),
.B1(n_225),
.B2(n_229),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_282),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_279),
.C(n_278),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_246),
.C(n_255),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_290),
.B(n_293),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_295),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_283),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_297),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_271),
.C(n_280),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_229),
.C(n_225),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_298),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_276),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_300),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_211),
.C(n_205),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_313),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_307),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_275),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_211),
.B1(n_9),
.B2(n_10),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_308),
.B(n_309),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_7),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_SL g312 ( 
.A(n_297),
.B(n_7),
.Y(n_312)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_10),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_293),
.C(n_285),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_320),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_302),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_321),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_306),
.A2(n_294),
.B1(n_300),
.B2(n_290),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_303),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_301),
.B(n_11),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_11),
.Y(n_325)
);

NOR2x1_ASAP7_75t_SL g323 ( 
.A(n_315),
.B(n_310),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_323),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_316),
.A2(n_311),
.B1(n_305),
.B2(n_14),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_325),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_305),
.B(n_14),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.C(n_321),
.Y(n_332)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_314),
.A2(n_13),
.B(n_15),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_330),
.B(n_331),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_326),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_329),
.B1(n_318),
.B2(n_16),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_15),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_337),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_15),
.Y(n_339)
);


endmodule