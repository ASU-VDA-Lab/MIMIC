module fake_jpeg_23677_n_305 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_305);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

BUFx2_ASAP7_75t_SL g55 ( 
.A(n_28),
.Y(n_55)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_37),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_34),
.Y(n_47)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_45),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_20),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_13),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_34),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_22),
.B1(n_16),
.B2(n_23),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_70),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2x1_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_28),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_74),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_39),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_35),
.B1(n_30),
.B2(n_16),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_73),
.B1(n_29),
.B2(n_30),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_30),
.B1(n_35),
.B2(n_16),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_40),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_56),
.B(n_34),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_72),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_75),
.B1(n_74),
.B2(n_59),
.Y(n_102)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_85),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_76),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_35),
.B1(n_30),
.B2(n_29),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_89),
.B1(n_99),
.B2(n_47),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_94),
.Y(n_122)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_35),
.B1(n_29),
.B2(n_23),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_90),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_82),
.C(n_78),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_114),
.C(n_33),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_111),
.B1(n_95),
.B2(n_43),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_109),
.B(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_66),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_33),
.C(n_65),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_77),
.B(n_19),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_38),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_110),
.B(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_65),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_123),
.B(n_125),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_91),
.B1(n_87),
.B2(n_84),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_124),
.A2(n_126),
.B1(n_147),
.B2(n_107),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_80),
.B1(n_83),
.B2(n_51),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_131),
.B(n_109),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_100),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_144),
.B1(n_96),
.B2(n_98),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_108),
.B(n_106),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_145),
.C(n_68),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_135),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_140),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_117),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_51),
.B1(n_95),
.B2(n_49),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_33),
.C(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_122),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_53),
.B1(n_60),
.B2(n_94),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_167),
.B1(n_171),
.B2(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_153),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_129),
.Y(n_184)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_159),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_119),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_13),
.B(n_18),
.Y(n_198)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_157),
.Y(n_197)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_107),
.B1(n_47),
.B2(n_109),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_100),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_143),
.B(n_135),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_133),
.C(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_118),
.B1(n_120),
.B2(n_115),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_60),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_172),
.A2(n_166),
.B1(n_157),
.B2(n_159),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_39),
.B1(n_14),
.B2(n_19),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_153),
.B(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_177),
.B(n_191),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_179),
.A2(n_194),
.B1(n_178),
.B2(n_185),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_150),
.C(n_164),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_189),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_162),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_190),
.A2(n_160),
.B(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

AOI21x1_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_13),
.B(n_18),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_18),
.B(n_63),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_122),
.B1(n_120),
.B2(n_115),
.Y(n_194)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_198),
.B(n_22),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_199),
.A2(n_212),
.B(n_24),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_168),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_186),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_203),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_164),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_210),
.C(n_214),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_64),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_207),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_63),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_39),
.C(n_48),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_194),
.B1(n_182),
.B2(n_196),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_48),
.C(n_31),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_178),
.B1(n_180),
.B2(n_187),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_27),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_219),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_181),
.B(n_27),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_221),
.B(n_232),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_230),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_208),
.A2(n_197),
.B1(n_187),
.B2(n_176),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_235),
.B1(n_218),
.B2(n_24),
.Y(n_246)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_176),
.Y(n_229)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_209),
.B(n_193),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_197),
.C(n_181),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_219),
.C(n_201),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_237),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_14),
.B(n_26),
.Y(n_234)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_26),
.B1(n_19),
.B2(n_14),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_214),
.B(n_26),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_15),
.B(n_5),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_227),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_243),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_244),
.C(n_220),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_207),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_222),
.C(n_220),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_0),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_246),
.A2(n_247),
.B1(n_253),
.B2(n_7),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_203),
.B(n_15),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_250),
.A2(n_255),
.B(n_235),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_8),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_222),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_8),
.B(n_12),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_261),
.C(n_265),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_243),
.A2(n_225),
.B(n_236),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_11),
.C(n_5),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_223),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_260),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_236),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_7),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_264),
.A2(n_266),
.B1(n_268),
.B2(n_258),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_6),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_241),
.B1(n_249),
.B2(n_254),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_1),
.C(n_2),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_1),
.C(n_2),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_9),
.B1(n_11),
.B2(n_5),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_247),
.B1(n_245),
.B2(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_277),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_21),
.B1(n_17),
.B2(n_10),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_21),
.B1(n_31),
.B2(n_4),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_3),
.C(n_4),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_279),
.B(n_3),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_2),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_257),
.Y(n_284)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_285),
.B(n_287),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_286),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_280),
.B(n_4),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_17),
.B(n_21),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_4),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_290),
.A2(n_276),
.B1(n_21),
.B2(n_31),
.Y(n_296)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_281),
.B(n_278),
.Y(n_293)
);

OA21x2_ASAP7_75t_SL g299 ( 
.A1(n_293),
.A2(n_274),
.B(n_31),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_289),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_294),
.B(n_283),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_298),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_291),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_303),
.A2(n_295),
.B1(n_299),
.B2(n_292),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_292),
.Y(n_305)
);


endmodule