module fake_jpeg_872_n_262 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_51),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_50),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_57),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_67),
.Y(n_97)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g113 ( 
.A(n_62),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_9),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_63),
.B(n_68),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_28),
.B(n_9),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_26),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_71),
.Y(n_102)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_4),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_4),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_32),
.C(n_63),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_16),
.B(n_4),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_78),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_21),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_30),
.B1(n_34),
.B2(n_42),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_17),
.B(n_5),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_24),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_65),
.Y(n_107)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_6),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_32),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_21),
.B1(n_18),
.B2(n_17),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_83),
.A2(n_85),
.B1(n_89),
.B2(n_91),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_18),
.B1(n_41),
.B2(n_33),
.Y(n_85)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_41),
.B1(n_33),
.B2(n_27),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_27),
.B1(n_23),
.B2(n_42),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_106),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_39),
.B1(n_34),
.B2(n_24),
.Y(n_106)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_49),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_118),
.Y(n_134)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_45),
.B(n_26),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_52),
.B(n_26),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_124),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_126),
.Y(n_151)
);

BUFx16f_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_32),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_99),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_135),
.C(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_75),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_132),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_131),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_86),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_75),
.C(n_50),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_70),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_144),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_121),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_150),
.Y(n_177)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_74),
.C(n_81),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_74),
.C(n_56),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_90),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_154),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_97),
.B(n_66),
.C(n_59),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_90),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_58),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_157),
.A2(n_111),
.B1(n_94),
.B2(n_92),
.Y(n_176)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_SL g172 ( 
.A(n_158),
.B(n_108),
.C(n_59),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g160 ( 
.A(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_172),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_154),
.B1(n_151),
.B2(n_135),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_176),
.B1(n_179),
.B2(n_116),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_147),
.A2(n_91),
.B(n_83),
.C(n_89),
.Y(n_163)
);

BUFx24_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_98),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_149),
.C(n_148),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_112),
.B1(n_88),
.B2(n_125),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_169),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_125),
.B1(n_122),
.B2(n_104),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_170),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_127),
.A2(n_122),
.B1(n_53),
.B2(n_104),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_127),
.A2(n_92),
.B1(n_94),
.B2(n_98),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_113),
.B1(n_95),
.B2(n_93),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_184),
.C(n_198),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_153),
.C(n_133),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_189),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_157),
.B1(n_140),
.B2(n_131),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_188),
.A2(n_167),
.B1(n_179),
.B2(n_159),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_134),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_136),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_194),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_163),
.Y(n_215)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_193),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_141),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_144),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_196),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_140),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_108),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

NOR4xp25_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_142),
.C(n_139),
.D(n_48),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_111),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_207),
.B1(n_214),
.B2(n_186),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_194),
.A2(n_180),
.B(n_163),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_163),
.B1(n_181),
.B2(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_190),
.B1(n_199),
.B2(n_196),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_177),
.B(n_168),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_191),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_230),
.C(n_211),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_221),
.B(n_204),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_226),
.Y(n_235)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_229),
.B1(n_207),
.B2(n_217),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_215),
.A2(n_190),
.B1(n_187),
.B2(n_199),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_184),
.C(n_183),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_237),
.C(n_218),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_215),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_238),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_216),
.C(n_206),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_239),
.B(n_204),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_242),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_232),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_231),
.C(n_237),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_250),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_227),
.B(n_222),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_227),
.B(n_235),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_229),
.B(n_205),
.C(n_222),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_247),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_210),
.A3(n_228),
.B1(n_208),
.B2(n_193),
.C1(n_202),
.C2(n_209),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_248),
.C(n_185),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_256),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_249),
.C(n_247),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_168),
.B(n_164),
.Y(n_260)
);

AOI32xp33_ASAP7_75t_L g261 ( 
.A1(n_260),
.A2(n_258),
.A3(n_142),
.B1(n_164),
.B2(n_95),
.Y(n_261)
);

XNOR2x2_ASAP7_75t_SL g262 ( 
.A(n_261),
.B(n_142),
.Y(n_262)
);


endmodule