module fake_jpeg_19484_n_395 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_15),
.B(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_41),
.B(n_60),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_53),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_57),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_15),
.B(n_14),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_25),
.Y(n_82)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_38),
.A2(n_39),
.B1(n_47),
.B2(n_66),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_70),
.A2(n_95),
.B1(n_99),
.B2(n_101),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_32),
.B1(n_30),
.B2(n_34),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_71),
.A2(n_86),
.B1(n_103),
.B2(n_59),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_32),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_82),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_16),
.B1(n_22),
.B2(n_34),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_87),
.B1(n_21),
.B2(n_31),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_16),
.B1(n_22),
.B2(n_34),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_43),
.A2(n_16),
.B1(n_22),
.B2(n_29),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_89),
.B(n_96),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_36),
.A2(n_64),
.B1(n_52),
.B2(n_20),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_33),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_58),
.A2(n_26),
.B1(n_18),
.B2(n_29),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_31),
.B1(n_21),
.B2(n_18),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_63),
.A2(n_17),
.B1(n_26),
.B2(n_31),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_17),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_108),
.B(n_114),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_109),
.A2(n_67),
.B1(n_104),
.B2(n_73),
.Y(n_178)
);

AOI22x1_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_55),
.B1(n_45),
.B2(n_62),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_111),
.A2(n_73),
.B1(n_93),
.B2(n_88),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_127),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_77),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_33),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_116),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_21),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_118),
.B(n_128),
.Y(n_184)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_72),
.B(n_25),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_121),
.B(n_122),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_77),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_74),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_123),
.B(n_134),
.Y(n_163)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_33),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_14),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_91),
.A2(n_25),
.B1(n_59),
.B2(n_27),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_129),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_33),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_146),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_0),
.B(n_1),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_76),
.B(n_89),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_142),
.B1(n_70),
.B2(n_92),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_99),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_135),
.B(n_136),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_81),
.B(n_1),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_139),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_96),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_75),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_140),
.B(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_2),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_3),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_92),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_75),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_78),
.Y(n_145)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_2),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_151),
.A2(n_160),
.B1(n_162),
.B2(n_185),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_153),
.A2(n_123),
.B(n_113),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_164),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_90),
.B1(n_69),
.B2(n_98),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_69),
.B1(n_98),
.B2(n_78),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_74),
.Y(n_164)
);

XNOR2x1_ASAP7_75t_SL g165 ( 
.A(n_128),
.B(n_105),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_SL g218 ( 
.A(n_165),
.B(n_167),
.C(n_93),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_104),
.B(n_106),
.C(n_76),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_183),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_100),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_182),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_110),
.B(n_93),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_173),
.A2(n_116),
.B(n_131),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_181),
.B1(n_111),
.B2(n_116),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_112),
.B(n_3),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_115),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_120),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_153),
.A2(n_132),
.B(n_130),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_186),
.A2(n_195),
.B(n_197),
.Y(n_237)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_144),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_190),
.B(n_191),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_122),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_193),
.B(n_223),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_134),
.B1(n_110),
.B2(n_114),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_208),
.B1(n_209),
.B2(n_181),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_126),
.B1(n_111),
.B2(n_107),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_198),
.B(n_202),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_156),
.B(n_118),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_203),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_201),
.A2(n_216),
.B1(n_168),
.B2(n_176),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_150),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_131),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_204),
.A2(n_218),
.B1(n_220),
.B2(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_113),
.B(n_136),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_151),
.A2(n_147),
.B1(n_145),
.B2(n_133),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_172),
.A2(n_145),
.B1(n_119),
.B2(n_142),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_155),
.B(n_4),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_210),
.B(n_211),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_152),
.B(n_4),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_124),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_68),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_117),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_117),
.C(n_143),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_184),
.C(n_148),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_163),
.A2(n_143),
.B1(n_6),
.B2(n_8),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_158),
.B(n_68),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g220 ( 
.A(n_165),
.B(n_5),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_171),
.B(n_5),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_221),
.B(n_210),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_157),
.A2(n_6),
.B(n_8),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_171),
.B(n_8),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_225),
.A2(n_233),
.B1(n_235),
.B2(n_242),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_232),
.B(n_255),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_179),
.B1(n_170),
.B2(n_185),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_189),
.A2(n_173),
.B1(n_167),
.B2(n_160),
.Y(n_235)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

INVx13_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_241),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_169),
.B1(n_183),
.B2(n_168),
.Y(n_242)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_246),
.Y(n_272)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_198),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_258),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_199),
.C(n_197),
.Y(n_276)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_249),
.Y(n_266)
);

NOR4xp25_ASAP7_75t_SL g250 ( 
.A(n_218),
.B(n_148),
.C(n_174),
.D(n_11),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_250),
.A2(n_217),
.B(n_186),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_209),
.B1(n_194),
.B2(n_214),
.Y(n_265)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_205),
.Y(n_275)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_215),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_262),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_222),
.B(n_206),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_261),
.A2(n_264),
.B(n_268),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_254),
.B(n_204),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g263 ( 
.A(n_259),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_255),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_265),
.A2(n_270),
.B1(n_274),
.B2(n_242),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_259),
.B(n_196),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_267),
.B(n_284),
.Y(n_309)
);

XNOR2x1_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_186),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_237),
.A2(n_195),
.B(n_201),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_269),
.A2(n_283),
.B(n_250),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_203),
.B1(n_192),
.B2(n_197),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_225),
.A2(n_192),
.B1(n_197),
.B2(n_207),
.Y(n_274)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_233),
.C(n_235),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_223),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_243),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_232),
.B(n_221),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_280),
.Y(n_291)
);

OAI32xp33_ASAP7_75t_L g280 ( 
.A1(n_230),
.A2(n_197),
.A3(n_211),
.B1(n_196),
.B2(n_216),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_238),
.A2(n_174),
.B(n_68),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_174),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_227),
.B(n_243),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_227),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_236),
.Y(n_288)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_289),
.B(n_313),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_298),
.Y(n_317)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_293),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_287),
.C(n_272),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_295),
.A2(n_303),
.B1(n_228),
.B2(n_226),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_247),
.Y(n_296)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_296),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_246),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_244),
.Y(n_300)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_306),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_234),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_262),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_274),
.A2(n_229),
.B1(n_257),
.B2(n_231),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_261),
.A2(n_253),
.B(n_256),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_264),
.A2(n_240),
.B(n_234),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_312),
.Y(n_314)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_308),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_280),
.A2(n_231),
.B1(n_252),
.B2(n_229),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_265),
.B1(n_279),
.B2(n_269),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_258),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_311),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_285),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_SL g313 ( 
.A1(n_268),
.A2(n_239),
.A3(n_258),
.B1(n_228),
.B2(n_226),
.C1(n_240),
.C2(n_245),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_318),
.B(n_316),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_320),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_296),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_322),
.B(n_324),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_278),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_323),
.B(n_325),
.Y(n_340)
);

OA22x2_ASAP7_75t_L g324 ( 
.A1(n_307),
.A2(n_271),
.B1(n_286),
.B2(n_282),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_273),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_291),
.A2(n_271),
.B1(n_286),
.B2(n_282),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_303),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_331),
.A2(n_291),
.B1(n_312),
.B2(n_308),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_283),
.C(n_281),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_290),
.C(n_294),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_290),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_334),
.B(n_292),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_324),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_336),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_333),
.Y(n_362)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_327),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_342),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_339),
.A2(n_295),
.B1(n_321),
.B2(n_315),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_306),
.C(n_297),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_347),
.C(n_317),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_305),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_345),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_344),
.A2(n_330),
.B1(n_326),
.B2(n_329),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_293),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_320),
.A2(n_297),
.B1(n_301),
.B2(n_309),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_349),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_323),
.C(n_319),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_315),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_324),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_351),
.B(n_357),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_334),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_362),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_355),
.B(n_347),
.C(n_340),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_335),
.A2(n_329),
.B1(n_314),
.B2(n_331),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_358),
.B(n_359),
.Y(n_365)
);

OAI22x1_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_324),
.B1(n_333),
.B2(n_299),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_361),
.A2(n_299),
.B1(n_281),
.B2(n_288),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_239),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_360),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_SL g366 ( 
.A(n_361),
.B(n_337),
.Y(n_366)
);

AOI21xp33_ASAP7_75t_L g380 ( 
.A1(n_366),
.A2(n_236),
.B(n_175),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_355),
.C(n_348),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_372),
.C(n_364),
.Y(n_376)
);

AO21x1_ASAP7_75t_L g369 ( 
.A1(n_356),
.A2(n_349),
.B(n_340),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_370),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_371),
.B(n_358),
.C(n_352),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_245),
.C(n_241),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_175),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_241),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_374),
.B(n_353),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_376),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_377),
.B(n_379),
.Y(n_383)
);

AO21x2_ASAP7_75t_L g387 ( 
.A1(n_380),
.A2(n_365),
.B(n_372),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_9),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_381),
.B(n_382),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_176),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_378),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_384),
.B(n_387),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_376),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_388),
.B(n_390),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_383),
.B(n_368),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_389),
.A2(n_386),
.B(n_387),
.Y(n_392)
);

A2O1A1O1Ixp25_ASAP7_75t_L g393 ( 
.A1(n_392),
.A2(n_382),
.B(n_369),
.C(n_11),
.D(n_10),
.Y(n_393)
);

O2A1O1Ixp33_ASAP7_75t_L g394 ( 
.A1(n_393),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_391),
.Y(n_395)
);


endmodule