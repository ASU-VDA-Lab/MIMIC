module fake_jpeg_28942_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx10_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_6),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_12),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_20),
.B(n_22),
.Y(n_23)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_7),
.A2(n_14),
.B1(n_13),
.B2(n_10),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_14),
.B1(n_13),
.B2(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_14),
.B1(n_17),
.B2(n_8),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_16),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_27),
.C(n_25),
.Y(n_36)
);

OAI22x1_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_16),
.B1(n_8),
.B2(n_20),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_32),
.B1(n_24),
.B2(n_8),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_35),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_8),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_27),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_28),
.C(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_5),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_31),
.B1(n_32),
.B2(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_36),
.C(n_39),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_4),
.B1(n_42),
.B2(n_47),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_3),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_51),
.B(n_4),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_3),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_3),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_52),
.A2(n_53),
.B(n_49),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_51),
.B2(n_53),
.Y(n_57)
);


endmodule