module real_jpeg_24830_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_113),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_1),
.A2(n_26),
.B1(n_33),
.B2(n_113),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_113),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g58 ( 
.A(n_4),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_5),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_90),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_90),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_5),
.A2(n_26),
.B1(n_33),
.B2(n_90),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_6),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_6),
.A2(n_32),
.B1(n_65),
.B2(n_66),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_6),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_6),
.A2(n_32),
.B1(n_59),
.B2(n_60),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_7),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_7),
.B(n_73),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_7),
.B(n_26),
.C(n_40),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_161),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_7),
.B(n_93),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_7),
.A2(n_25),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_10),
.A2(n_63),
.B1(n_158),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_10),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_165),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_165),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_10),
.A2(n_26),
.B1(n_33),
.B2(n_165),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_11),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_11),
.A2(n_64),
.B1(n_65),
.B2(n_154),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_154),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_154),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_13),
.A2(n_48),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_48),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_13),
.A2(n_48),
.B1(n_59),
.B2(n_60),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_14),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_14),
.A2(n_26),
.B1(n_33),
.B2(n_45),
.Y(n_144)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_15),
.Y(n_180)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_15),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_135),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_115),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_20),
.B(n_115),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.C(n_95),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_21),
.A2(n_75),
.B1(n_76),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_21),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_50),
.B2(n_74),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_22),
.A2(n_51),
.B(n_53),
.Y(n_133)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_24),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_24),
.A2(n_34),
.B1(n_51),
.B2(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_30),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_25),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_25),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_25),
.A2(n_144),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_25),
.A2(n_101),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_25),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_25),
.A2(n_226),
.B1(n_233),
.B2(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_33),
.B1(n_40),
.B2(n_42),
.Y(n_43)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g198 ( 
.A(n_27),
.Y(n_198)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_27),
.Y(n_240)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_28),
.B(n_104),
.Y(n_146)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_31),
.B(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_31),
.A2(n_146),
.B(n_224),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_33),
.B(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_34),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_44),
.B(n_46),
.Y(n_34)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_35),
.A2(n_43),
.B1(n_44),
.B2(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_35),
.A2(n_43),
.B(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_35),
.A2(n_46),
.B(n_128),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_35),
.A2(n_43),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_35),
.A2(n_43),
.B1(n_211),
.B2(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_35),
.A2(n_78),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_43),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_37),
.A2(n_38),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g252 ( 
.A(n_37),
.B(n_60),
.C(n_86),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_38),
.B(n_207),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_38),
.A2(n_85),
.B(n_251),
.C(n_252),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_43),
.A2(n_80),
.B(n_106),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_43),
.B(n_161),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_49),
.A2(n_81),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_67),
.B(n_69),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_54),
.A2(n_111),
.B(n_114),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_54),
.A2(n_56),
.B1(n_164),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_55),
.B(n_70),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_55),
.A2(n_73),
.B1(n_157),
.B2(n_163),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_55),
.A2(n_73),
.B1(n_112),
.B2(n_171),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_56),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_58),
.B1(n_63),
.B2(n_66),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_57),
.A2(n_60),
.B(n_162),
.C(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_58),
.B(n_59),
.C(n_64),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_60),
.B1(n_85),
.B2(n_86),
.Y(n_87)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g251 ( 
.A(n_60),
.B(n_161),
.CON(n_251),
.SN(n_251)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_65),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_66),
.B(n_161),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_68),
.B(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_82),
.B(n_94),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_82),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_88),
.B1(n_91),
.B2(n_93),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_83),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_83),
.A2(n_93),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_83),
.A2(n_93),
.B1(n_192),
.B2(n_251),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_89),
.B(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_84),
.A2(n_125),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_93),
.B(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_93),
.B(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_117),
.B1(n_131),
.B2(n_132),
.Y(n_116)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_95),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_107),
.C(n_110),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_96),
.A2(n_97),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_105),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_98),
.A2(n_99),
.B1(n_105),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_103),
.A2(n_179),
.B(n_198),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_105),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_107),
.B(n_110),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_133),
.Y(n_115)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_130),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_129),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g293 ( 
.A1(n_125),
.A2(n_126),
.B(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_127),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_312),
.B(n_317),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_301),
.B(n_311),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_199),
.B(n_283),
.C(n_300),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_184),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_139),
.B(n_184),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_166),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_148),
.B2(n_149),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_141),
.B(n_149),
.C(n_166),
.Y(n_284)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_143),
.B(n_147),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_156),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_153),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_155),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_186),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_161),
.B(n_162),
.Y(n_157)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_161),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_176),
.B2(n_183),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_169),
.B(n_172),
.C(n_183),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_175),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_176),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_181),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.C(n_189),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_185),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_188),
.B(n_189),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.C(n_196),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_190),
.B(n_268),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_268)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_282),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_277),
.B(n_281),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_263),
.B(n_276),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_247),
.B(n_262),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_221),
.B(n_246),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_212),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_208),
.B1(n_209),
.B2(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_219),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_214),
.B(n_217),
.C(n_219),
.Y(n_261)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_220),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_230),
.B(n_245),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_228),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_241),
.B(n_244),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_237),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_242),
.B(n_243),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_261),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_261),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_256),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_257),
.C(n_260),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_253),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_264),
.B(n_265),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_272),
.C(n_274),
.Y(n_280)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_280),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_285),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_299),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_295),
.B1(n_297),
.B2(n_298),
.Y(n_286)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_291),
.C(n_292),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_295),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_297),
.C(n_299),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_303),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_310),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_307),
.C(n_310),
.Y(n_313)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);


endmodule