module real_aes_2326_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_0), .B(n_134), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_1), .A2(n_116), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_2), .B(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_3), .B(n_124), .Y(n_180) );
INVx1_ASAP7_75t_L g121 ( .A(n_4), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_5), .B(n_124), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_6), .B(n_111), .Y(n_461) );
INVx1_ASAP7_75t_L g489 ( .A(n_7), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g786 ( .A(n_8), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_9), .Y(n_504) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_10), .A2(n_99), .B1(n_779), .B2(n_790), .C1(n_802), .C2(n_806), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_10), .A2(n_103), .B1(n_772), .B2(n_793), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_10), .Y(n_793) );
NAND2xp33_ASAP7_75t_L g161 ( .A(n_11), .B(n_128), .Y(n_161) );
INVx2_ASAP7_75t_L g113 ( .A(n_12), .Y(n_113) );
AOI221x1_ASAP7_75t_L g203 ( .A1(n_13), .A2(n_25), .B1(n_116), .B2(n_134), .C(n_204), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_14), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_15), .B(n_134), .Y(n_157) );
AO21x2_ASAP7_75t_L g154 ( .A1(n_16), .A2(n_155), .B(n_156), .Y(n_154) );
INVx1_ASAP7_75t_L g470 ( .A(n_17), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_18), .B(n_147), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_19), .B(n_124), .Y(n_123) );
AO21x1_ASAP7_75t_L g175 ( .A1(n_20), .A2(n_134), .B(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g427 ( .A(n_21), .Y(n_427) );
INVx1_ASAP7_75t_L g468 ( .A(n_22), .Y(n_468) );
INVx1_ASAP7_75t_SL g454 ( .A(n_23), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_24), .B(n_135), .Y(n_548) );
NAND2x1_ASAP7_75t_L g189 ( .A(n_26), .B(n_124), .Y(n_189) );
AOI33xp33_ASAP7_75t_L g516 ( .A1(n_27), .A2(n_52), .A3(n_444), .B1(n_451), .B2(n_517), .B3(n_518), .Y(n_516) );
NAND2x1_ASAP7_75t_L g143 ( .A(n_28), .B(n_128), .Y(n_143) );
INVx1_ASAP7_75t_L g498 ( .A(n_29), .Y(n_498) );
OR2x2_ASAP7_75t_L g112 ( .A(n_30), .B(n_84), .Y(n_112) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_30), .A2(n_84), .B(n_113), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_31), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_32), .B(n_128), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_33), .B(n_124), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_34), .B(n_128), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_35), .A2(n_116), .B(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g117 ( .A(n_36), .B(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g132 ( .A(n_36), .B(n_121), .Y(n_132) );
INVx1_ASAP7_75t_L g450 ( .A(n_36), .Y(n_450) );
OR2x6_ASAP7_75t_L g425 ( .A(n_37), .B(n_426), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_38), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_39), .B(n_134), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_40), .B(n_442), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_41), .A2(n_111), .B1(n_151), .B2(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_42), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_43), .B(n_135), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_44), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_45), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_46), .B(n_128), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_47), .B(n_155), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_48), .B(n_135), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_49), .A2(n_116), .B(n_142), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_50), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_51), .B(n_128), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_53), .B(n_135), .Y(n_528) );
INVx1_ASAP7_75t_L g120 ( .A(n_54), .Y(n_120) );
INVx1_ASAP7_75t_L g130 ( .A(n_54), .Y(n_130) );
AND2x2_ASAP7_75t_L g529 ( .A(n_55), .B(n_147), .Y(n_529) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_56), .A2(n_72), .B1(n_442), .B2(n_448), .C(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_57), .B(n_442), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_58), .B(n_124), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_59), .B(n_151), .Y(n_506) );
AOI21xp5_ASAP7_75t_SL g478 ( .A1(n_60), .A2(n_448), .B(n_479), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_61), .A2(n_116), .B(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g464 ( .A(n_62), .Y(n_464) );
AO21x1_ASAP7_75t_L g177 ( .A1(n_63), .A2(n_116), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_64), .B(n_134), .Y(n_165) );
INVx1_ASAP7_75t_L g527 ( .A(n_65), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_66), .B(n_134), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_67), .A2(n_448), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g226 ( .A(n_68), .B(n_148), .Y(n_226) );
INVx1_ASAP7_75t_L g118 ( .A(n_69), .Y(n_118) );
INVx1_ASAP7_75t_L g126 ( .A(n_69), .Y(n_126) );
AND2x2_ASAP7_75t_L g149 ( .A(n_70), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_71), .B(n_442), .Y(n_519) );
AND2x2_ASAP7_75t_L g457 ( .A(n_73), .B(n_150), .Y(n_457) );
INVx1_ASAP7_75t_L g465 ( .A(n_74), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_75), .A2(n_448), .B(n_453), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_76), .A2(n_448), .B(n_511), .C(n_547), .Y(n_546) );
AOI22xp5_ASAP7_75t_SL g770 ( .A1(n_77), .A2(n_100), .B1(n_771), .B2(n_775), .Y(n_770) );
INVx1_ASAP7_75t_L g428 ( .A(n_78), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_79), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g163 ( .A(n_80), .B(n_150), .Y(n_163) );
AND2x2_ASAP7_75t_SL g476 ( .A(n_81), .B(n_150), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_82), .A2(n_448), .B1(n_514), .B2(n_515), .Y(n_513) );
AND2x2_ASAP7_75t_L g176 ( .A(n_83), .B(n_111), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_85), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g193 ( .A(n_86), .B(n_150), .Y(n_193) );
INVx1_ASAP7_75t_L g480 ( .A(n_87), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_88), .B(n_124), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_89), .A2(n_116), .B(n_122), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_90), .B(n_128), .Y(n_205) );
AND2x2_ASAP7_75t_L g520 ( .A(n_91), .B(n_150), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_92), .B(n_124), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_93), .A2(n_496), .B(n_497), .C(n_499), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_94), .Y(n_100) );
BUFx2_ASAP7_75t_L g787 ( .A(n_95), .Y(n_787) );
BUFx2_ASAP7_75t_SL g810 ( .A(n_95), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_96), .A2(n_116), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_97), .B(n_135), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_101), .B(n_770), .Y(n_99) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OAI22xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_420), .B1(n_429), .B2(n_433), .Y(n_102) );
INVx2_ASAP7_75t_L g772 ( .A(n_103), .Y(n_772) );
OR2x6_ASAP7_75t_L g103 ( .A(n_104), .B(n_318), .Y(n_103) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_105), .B(n_230), .C(n_285), .Y(n_104) );
AOI221xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_170), .B1(n_194), .B2(n_198), .C(n_208), .Y(n_105) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_153), .Y(n_106) );
AND2x2_ASAP7_75t_SL g196 ( .A(n_107), .B(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g229 ( .A(n_107), .Y(n_229) );
AND2x2_ASAP7_75t_L g274 ( .A(n_107), .B(n_211), .Y(n_274) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_138), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g262 ( .A(n_109), .Y(n_262) );
INVx1_ASAP7_75t_L g272 ( .A(n_109), .Y(n_272) );
AO21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_114), .B(n_136), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_110), .B(n_137), .Y(n_136) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_110), .A2(n_114), .B(n_136), .Y(n_236) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_111), .A2(n_157), .B(n_158), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_111), .B(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_111), .B(n_131), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_111), .A2(n_478), .B(n_482), .Y(n_477) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AND2x2_ASAP7_75t_SL g148 ( .A(n_112), .B(n_113), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_133), .Y(n_114) );
AND2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
BUFx3_ASAP7_75t_L g446 ( .A(n_117), .Y(n_446) );
AND2x6_ASAP7_75t_L g128 ( .A(n_118), .B(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g452 ( .A(n_118), .Y(n_452) );
AND2x4_ASAP7_75t_L g448 ( .A(n_119), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x4_ASAP7_75t_L g124 ( .A(n_120), .B(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g444 ( .A(n_120), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_121), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_127), .B(n_131), .Y(n_122) );
INVxp67_ASAP7_75t_L g471 ( .A(n_124), .Y(n_471) );
AND2x4_ASAP7_75t_L g135 ( .A(n_125), .B(n_129), .Y(n_135) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVxp67_ASAP7_75t_L g469 ( .A(n_128), .Y(n_469) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_131), .A2(n_143), .B(n_144), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_131), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_131), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_131), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_131), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_131), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_131), .A2(n_223), .B(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_SL g453 ( .A1(n_131), .A2(n_454), .B(n_455), .C(n_456), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_131), .A2(n_455), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_131), .A2(n_455), .B(n_489), .C(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g514 ( .A(n_131), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_131), .A2(n_455), .B(n_527), .C(n_528), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_131), .A2(n_548), .B(n_549), .Y(n_547) );
INVx5_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g134 ( .A(n_132), .B(n_135), .Y(n_134) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_132), .Y(n_499) );
INVx1_ASAP7_75t_L g466 ( .A(n_135), .Y(n_466) );
OR2x2_ASAP7_75t_L g251 ( .A(n_138), .B(n_154), .Y(n_251) );
NAND2x1p5_ASAP7_75t_L g282 ( .A(n_138), .B(n_197), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_138), .B(n_162), .Y(n_295) );
INVx2_ASAP7_75t_L g304 ( .A(n_138), .Y(n_304) );
AND2x2_ASAP7_75t_L g325 ( .A(n_138), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g409 ( .A(n_138), .B(n_228), .Y(n_409) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g237 ( .A(n_139), .B(n_162), .Y(n_237) );
AND2x2_ASAP7_75t_L g370 ( .A(n_139), .B(n_197), .Y(n_370) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_139), .Y(n_396) );
AO21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_146), .B(n_149), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
AO21x2_ASAP7_75t_L g439 ( .A1(n_146), .A2(n_440), .B(n_457), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_147), .A2(n_165), .B(n_166), .Y(n_164) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_147), .A2(n_203), .B(n_207), .Y(n_202) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_147), .A2(n_203), .B(n_207), .Y(n_214) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g192 ( .A(n_150), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_150), .A2(n_192), .B1(n_495), .B2(n_500), .Y(n_494) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_151), .B(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx4f_ASAP7_75t_L g155 ( .A(n_152), .Y(n_155) );
AND2x4_ASAP7_75t_L g324 ( .A(n_153), .B(n_325), .Y(n_324) );
AOI321xp33_ASAP7_75t_L g338 ( .A1(n_153), .A2(n_267), .A3(n_268), .B1(n_300), .B2(n_339), .C(n_342), .Y(n_338) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_162), .Y(n_153) );
BUFx3_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
INVx2_ASAP7_75t_L g228 ( .A(n_154), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_154), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g261 ( .A(n_154), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g294 ( .A(n_154), .Y(n_294) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_155), .A2(n_487), .B(n_491), .Y(n_486) );
INVx2_ASAP7_75t_SL g511 ( .A(n_155), .Y(n_511) );
INVx5_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
NOR2x1_ASAP7_75t_SL g246 ( .A(n_162), .B(n_236), .Y(n_246) );
BUFx2_ASAP7_75t_L g341 ( .A(n_162), .Y(n_341) );
OR2x6_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
INVxp67_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_183), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g239 ( .A(n_172), .B(n_240), .Y(n_239) );
NOR4xp25_ASAP7_75t_L g342 ( .A(n_172), .B(n_336), .C(n_340), .D(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g380 ( .A(n_172), .Y(n_380) );
AND2x2_ASAP7_75t_L g414 ( .A(n_172), .B(n_354), .Y(n_414) );
BUFx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g215 ( .A(n_173), .Y(n_215) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g269 ( .A(n_174), .Y(n_269) );
OAI21x1_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_177), .B(n_181), .Y(n_174) );
INVx1_ASAP7_75t_L g182 ( .A(n_176), .Y(n_182) );
AOI33xp33_ASAP7_75t_L g410 ( .A1(n_183), .A2(n_212), .A3(n_243), .B1(n_259), .B2(n_365), .B3(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g200 ( .A(n_184), .B(n_201), .Y(n_200) );
AND2x4_ASAP7_75t_L g210 ( .A(n_184), .B(n_211), .Y(n_210) );
BUFx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g217 ( .A(n_185), .Y(n_217) );
INVxp67_ASAP7_75t_L g298 ( .A(n_185), .Y(n_298) );
AND2x2_ASAP7_75t_L g354 ( .A(n_185), .B(n_219), .Y(n_354) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_192), .B(n_193), .Y(n_185) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_186), .A2(n_192), .B(n_193), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_191), .Y(n_186) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_192), .A2(n_220), .B(n_226), .Y(n_219) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_192), .A2(n_220), .B(n_226), .Y(n_255) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_192), .A2(n_523), .B(n_529), .Y(n_522) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_192), .A2(n_523), .B(n_529), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_194), .A2(n_376), .B(n_377), .Y(n_375) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
AND2x2_ASAP7_75t_L g363 ( .A(n_195), .B(n_237), .Y(n_363) );
AND3x2_ASAP7_75t_L g365 ( .A(n_195), .B(n_249), .C(n_304), .Y(n_365) );
INVx3_ASAP7_75t_SL g317 ( .A(n_196), .Y(n_317) );
INVx4_ASAP7_75t_L g211 ( .A(n_197), .Y(n_211) );
AND2x2_ASAP7_75t_L g249 ( .A(n_197), .B(n_236), .Y(n_249) );
INVxp67_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx2_ASAP7_75t_L g243 ( .A(n_201), .Y(n_243) );
AND2x4_ASAP7_75t_L g268 ( .A(n_201), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g331 ( .A(n_201), .B(n_219), .Y(n_331) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g301 ( .A(n_202), .Y(n_301) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_202), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_R g208 ( .A1(n_209), .A2(n_212), .B(n_216), .C(n_227), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g260 ( .A(n_211), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_211), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_211), .B(n_228), .Y(n_389) );
INVx1_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g371 ( .A(n_213), .B(n_361), .Y(n_371) );
AND2x2_ASAP7_75t_SL g213 ( .A(n_214), .B(n_215), .Y(n_213) );
AND2x2_ASAP7_75t_L g218 ( .A(n_214), .B(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g240 ( .A(n_214), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g256 ( .A(n_214), .B(n_257), .Y(n_256) );
AND2x4_ASAP7_75t_L g289 ( .A(n_214), .B(n_269), .Y(n_289) );
AND2x4_ASAP7_75t_L g254 ( .A(n_215), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g278 ( .A(n_215), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g316 ( .A(n_215), .B(n_241), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
AND2x2_ASAP7_75t_L g244 ( .A(n_217), .B(n_241), .Y(n_244) );
AND2x2_ASAP7_75t_L g259 ( .A(n_217), .B(n_219), .Y(n_259) );
BUFx2_ASAP7_75t_L g315 ( .A(n_217), .Y(n_315) );
AND2x2_ASAP7_75t_L g329 ( .A(n_217), .B(n_240), .Y(n_329) );
INVx2_ASAP7_75t_L g241 ( .A(n_219), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_221), .B(n_225), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g277 ( .A1(n_227), .A2(n_278), .B1(n_280), .B2(n_284), .Y(n_277) );
INVx2_ASAP7_75t_SL g308 ( .A(n_227), .Y(n_308) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
AND2x2_ASAP7_75t_L g283 ( .A(n_228), .B(n_236), .Y(n_283) );
INVx1_ASAP7_75t_L g390 ( .A(n_229), .Y(n_390) );
NOR3xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_263), .C(n_277), .Y(n_230) );
OAI221xp5_ASAP7_75t_SL g231 ( .A1(n_232), .A2(n_238), .B1(n_242), .B2(n_245), .C(n_247), .Y(n_231) );
INVx1_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_237), .Y(n_233) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g291 ( .A(n_235), .Y(n_291) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_235), .Y(n_419) );
INVx1_ASAP7_75t_L g382 ( .A(n_237), .Y(n_382) );
AND2x2_ASAP7_75t_SL g392 ( .A(n_237), .B(n_261), .Y(n_392) );
INVxp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_241), .B(n_269), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
OR2x2_ASAP7_75t_L g275 ( .A(n_243), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g353 ( .A(n_243), .Y(n_353) );
AND2x2_ASAP7_75t_L g288 ( .A(n_244), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g334 ( .A(n_246), .B(n_294), .Y(n_334) );
AND2x2_ASAP7_75t_L g411 ( .A(n_246), .B(n_409), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_252), .B1(n_259), .B2(n_260), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g270 ( .A(n_251), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
INVx2_ASAP7_75t_L g276 ( .A(n_254), .Y(n_276) );
AND2x4_ASAP7_75t_L g300 ( .A(n_254), .B(n_301), .Y(n_300) );
OAI21xp33_ASAP7_75t_SL g330 ( .A1(n_254), .A2(n_331), .B(n_332), .Y(n_330) );
AND2x2_ASAP7_75t_L g357 ( .A(n_254), .B(n_315), .Y(n_357) );
INVx2_ASAP7_75t_L g279 ( .A(n_255), .Y(n_279) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_255), .Y(n_312) );
INVx1_ASAP7_75t_SL g336 ( .A(n_256), .Y(n_336) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx2_ASAP7_75t_L g267 ( .A(n_258), .Y(n_267) );
AND2x4_ASAP7_75t_SL g361 ( .A(n_258), .B(n_279), .Y(n_361) );
AND2x2_ASAP7_75t_L g358 ( .A(n_261), .B(n_304), .Y(n_358) );
AND2x2_ASAP7_75t_L g384 ( .A(n_261), .B(n_370), .Y(n_384) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_262), .Y(n_306) );
INVx1_ASAP7_75t_L g326 ( .A(n_262), .Y(n_326) );
OAI22xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_270), .B1(n_273), .B2(n_275), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_268), .B(n_279), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_268), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g407 ( .A(n_268), .Y(n_407) );
INVx2_ASAP7_75t_SL g332 ( .A(n_270), .Y(n_332) );
AND2x2_ASAP7_75t_L g344 ( .A(n_272), .B(n_304), .Y(n_344) );
INVx2_ASAP7_75t_L g350 ( .A(n_272), .Y(n_350) );
INVxp33_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g309 ( .A(n_275), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_278), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g400 ( .A(n_278), .Y(n_400) );
INVx1_ASAP7_75t_L g328 ( .A(n_280), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_281), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g339 ( .A(n_283), .B(n_340), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_283), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_412) );
NOR3xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_307), .C(n_310), .Y(n_285) );
OAI221xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_290), .B1(n_292), .B2(n_296), .C(n_299), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_SL g405 ( .A(n_290), .Y(n_405) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g374 ( .A(n_291), .B(n_340), .Y(n_374) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g305 ( .A(n_294), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g376 ( .A(n_296), .Y(n_376) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g373 ( .A(n_297), .Y(n_373) );
INVx1_ASAP7_75t_L g379 ( .A(n_298), .Y(n_379) );
OR2x2_ASAP7_75t_L g402 ( .A(n_298), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_SL g311 ( .A(n_301), .Y(n_311) );
AND2x2_ASAP7_75t_L g381 ( .A(n_301), .B(n_361), .Y(n_381) );
AND2x2_ASAP7_75t_SL g413 ( .A(n_301), .B(n_314), .Y(n_413) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g418 ( .A(n_304), .Y(n_418) );
INVx1_ASAP7_75t_L g368 ( .A(n_306), .Y(n_368) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B(n_313), .C(n_317), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_311), .B(n_361), .Y(n_385) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_314), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g322 ( .A(n_316), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g403 ( .A(n_316), .Y(n_403) );
NAND4xp75_ASAP7_75t_L g318 ( .A(n_319), .B(n_375), .C(n_391), .D(n_412), .Y(n_318) );
NOR3x1_ASAP7_75t_L g319 ( .A(n_320), .B(n_337), .C(n_359), .Y(n_319) );
NAND4xp75_ASAP7_75t_L g320 ( .A(n_321), .B(n_327), .C(n_330), .D(n_333), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_322), .B(n_324), .Y(n_321) );
AND2x2_ASAP7_75t_L g372 ( .A(n_323), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g397 ( .A(n_324), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_SL g386 ( .A(n_329), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_345), .Y(n_337) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_341), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_351), .B(n_355), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI322xp33_ASAP7_75t_L g377 ( .A1(n_349), .A2(n_378), .A3(n_382), .B1(n_383), .B2(n_385), .C1(n_386), .C2(n_387), .Y(n_377) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_350), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_353), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_354), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
OAI211xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B(n_364), .C(n_366), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B1(n_372), .B2(n_374), .Y(n_366) );
NOR2xp33_ASAP7_75t_SL g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B(n_381), .Y(n_378) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_384), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g394 ( .A(n_389), .B(n_395), .Y(n_394) );
O2A1O1Ixp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_398), .C(n_401), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_394), .B(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI221xp5_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_404), .B1(n_406), .B2(n_408), .C(n_410), .Y(n_401) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
CKINVDCx6p67_ASAP7_75t_R g420 ( .A(n_421), .Y(n_420) );
INVx4_ASAP7_75t_SL g773 ( .A(n_421), .Y(n_773) );
INVx3_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_423), .Y(n_422) );
AND2x6_ASAP7_75t_SL g423 ( .A(n_424), .B(n_425), .Y(n_423) );
OR2x6_ASAP7_75t_SL g431 ( .A(n_424), .B(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g778 ( .A(n_424), .B(n_425), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_424), .B(n_432), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_425), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
CKINVDCx11_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
OAI22x1_ASAP7_75t_L g771 ( .A1(n_431), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_771) );
INVx1_ASAP7_75t_L g774 ( .A(n_433), .Y(n_774) );
OR3x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_635), .C(n_706), .Y(n_433) );
NAND3x1_ASAP7_75t_SL g434 ( .A(n_435), .B(n_562), .C(n_584), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_552), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_483), .B1(n_530), .B2(n_534), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_437), .A2(n_738), .B1(n_739), .B2(n_741), .Y(n_737) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_458), .Y(n_437) );
AND2x2_ASAP7_75t_L g553 ( .A(n_438), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_438), .B(n_600), .Y(n_619) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g537 ( .A(n_439), .Y(n_537) );
AND2x2_ASAP7_75t_L g587 ( .A(n_439), .B(n_460), .Y(n_587) );
INVx1_ASAP7_75t_L g626 ( .A(n_439), .Y(n_626) );
OR2x2_ASAP7_75t_L g663 ( .A(n_439), .B(n_475), .Y(n_663) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_439), .Y(n_675) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_439), .Y(n_699) );
AND2x2_ASAP7_75t_L g756 ( .A(n_439), .B(n_583), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_447), .Y(n_440) );
INVx1_ASAP7_75t_L g507 ( .A(n_442), .Y(n_507) );
AND2x4_ASAP7_75t_L g442 ( .A(n_443), .B(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g543 ( .A(n_443), .Y(n_543) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
OR2x6_ASAP7_75t_L g455 ( .A(n_444), .B(n_452), .Y(n_455) );
INVxp33_ASAP7_75t_L g517 ( .A(n_444), .Y(n_517) );
INVx1_ASAP7_75t_L g544 ( .A(n_446), .Y(n_544) );
INVxp67_ASAP7_75t_L g505 ( .A(n_448), .Y(n_505) );
NOR2x1p5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g518 ( .A(n_451), .Y(n_518) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_455), .A2(n_464), .B1(n_465), .B2(n_466), .Y(n_463) );
INVxp67_ASAP7_75t_L g496 ( .A(n_455), .Y(n_496) );
INVx2_ASAP7_75t_L g550 ( .A(n_455), .Y(n_550) );
NOR2x1_ASAP7_75t_L g458 ( .A(n_459), .B(n_473), .Y(n_458) );
INVx1_ASAP7_75t_L g631 ( .A(n_459), .Y(n_631) );
AND2x2_ASAP7_75t_L g657 ( .A(n_459), .B(n_475), .Y(n_657) );
NAND2x1_ASAP7_75t_L g673 ( .A(n_459), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g554 ( .A(n_460), .B(n_540), .Y(n_554) );
INVx3_ASAP7_75t_L g583 ( .A(n_460), .Y(n_583) );
NOR2x1_ASAP7_75t_SL g702 ( .A(n_460), .B(n_475), .Y(n_702) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_467), .B(n_472), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_466), .B(n_498), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_470), .B2(n_471), .Y(n_467) );
NOR2x1_ASAP7_75t_L g610 ( .A(n_473), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g581 ( .A(n_474), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx4_ASAP7_75t_L g551 ( .A(n_475), .Y(n_551) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_475), .Y(n_596) );
AND2x2_ASAP7_75t_L g668 ( .A(n_475), .B(n_540), .Y(n_668) );
AND2x4_ASAP7_75t_L g685 ( .A(n_475), .B(n_629), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_475), .B(n_627), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_475), .B(n_536), .Y(n_761) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_483), .A2(n_578), .B1(n_649), .B2(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_508), .Y(n_483) );
INVx2_ASAP7_75t_L g651 ( .A(n_484), .Y(n_651) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_492), .Y(n_484) );
BUFx3_ASAP7_75t_L g641 ( .A(n_485), .Y(n_641) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_486), .B(n_510), .Y(n_533) );
INVx2_ASAP7_75t_L g557 ( .A(n_486), .Y(n_557) );
INVx1_ASAP7_75t_L g569 ( .A(n_486), .Y(n_569) );
AND2x4_ASAP7_75t_L g576 ( .A(n_486), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g593 ( .A(n_486), .B(n_493), .Y(n_593) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_486), .Y(n_607) );
INVxp67_ASAP7_75t_L g615 ( .A(n_486), .Y(n_615) );
AND2x2_ASAP7_75t_L g644 ( .A(n_492), .B(n_560), .Y(n_644) );
AND2x2_ASAP7_75t_L g660 ( .A(n_492), .B(n_561), .Y(n_660) );
NOR2xp67_ASAP7_75t_L g747 ( .A(n_492), .B(n_560), .Y(n_747) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g556 ( .A(n_493), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g567 ( .A(n_493), .Y(n_567) );
INVx1_ASAP7_75t_L g580 ( .A(n_493), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_493), .B(n_522), .Y(n_617) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_501), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_505), .B1(n_506), .B2(n_507), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g740 ( .A(n_508), .Y(n_740) );
AND2x4_ASAP7_75t_L g508 ( .A(n_509), .B(n_521), .Y(n_508) );
AND2x2_ASAP7_75t_L g614 ( .A(n_509), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g643 ( .A(n_509), .Y(n_643) );
AND2x2_ASAP7_75t_L g745 ( .A(n_509), .B(n_560), .Y(n_745) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_510), .B(n_522), .Y(n_605) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_520), .Y(n_510) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_511), .A2(n_512), .B(n_520), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_513), .B(n_519), .Y(n_512) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx3_ASAP7_75t_L g531 ( .A(n_521), .Y(n_531) );
NAND2x1p5_ASAP7_75t_L g720 ( .A(n_521), .B(n_641), .Y(n_720) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_522), .Y(n_634) );
AND2x2_ASAP7_75t_L g661 ( .A(n_522), .B(n_607), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
AND2x2_ASAP7_75t_L g575 ( .A(n_531), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g591 ( .A(n_531), .Y(n_591) );
AND2x2_ASAP7_75t_L g679 ( .A(n_531), .B(n_556), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_531), .B(n_699), .Y(n_704) );
AND2x2_ASAP7_75t_L g714 ( .A(n_531), .B(n_593), .Y(n_714) );
OR2x2_ASAP7_75t_L g751 ( .A(n_531), .B(n_651), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_532), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g711 ( .A(n_532), .B(n_567), .Y(n_711) );
AND2x2_ASAP7_75t_L g727 ( .A(n_532), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g721 ( .A(n_533), .B(n_617), .Y(n_721) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
INVx1_ASAP7_75t_L g603 ( .A(n_535), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_535), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g701 ( .A(n_535), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_535), .B(n_582), .Y(n_726) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_536), .Y(n_573) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_537), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_538), .A2(n_571), .B1(n_589), .B2(n_592), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_538), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g705 ( .A(n_538), .Y(n_705) );
AND2x4_ASAP7_75t_SL g538 ( .A(n_539), .B(n_551), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g582 ( .A(n_540), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g602 ( .A(n_540), .Y(n_602) );
INVx1_ASAP7_75t_L g629 ( .A(n_540), .Y(n_629) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_546), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .C(n_545), .Y(n_542) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_551), .Y(n_571) );
AND2x4_ASAP7_75t_L g628 ( .A(n_551), .B(n_629), .Y(n_628) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_551), .B(n_658), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
AND2x2_ASAP7_75t_L g653 ( .A(n_553), .B(n_596), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_553), .A2(n_734), .B(n_735), .Y(n_733) );
INVx2_ASAP7_75t_L g611 ( .A(n_554), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_555), .A2(n_665), .B1(n_669), .B2(n_672), .Y(n_664) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_556), .Y(n_622) );
AND2x2_ASAP7_75t_L g632 ( .A(n_556), .B(n_633), .Y(n_632) );
INVx3_ASAP7_75t_L g671 ( .A(n_556), .Y(n_671) );
NAND2x1_ASAP7_75t_SL g696 ( .A(n_556), .B(n_565), .Y(n_696) );
AND2x2_ASAP7_75t_L g592 ( .A(n_558), .B(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NOR2x1_ASAP7_75t_L g568 ( .A(n_560), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g565 ( .A(n_561), .Y(n_565) );
INVx2_ASAP7_75t_L g577 ( .A(n_561), .Y(n_577) );
AOI21xp5_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_570), .B(n_574), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_565), .B(n_759), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_566), .A2(n_655), .B1(n_659), .B2(n_662), .Y(n_654) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
BUFx2_ASAP7_75t_L g759 ( .A(n_567), .Y(n_759) );
INVx1_ASAP7_75t_SL g766 ( .A(n_567), .Y(n_766) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_568), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OA21x2_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_578), .B(n_581), .Y(n_574) );
AND2x2_ASAP7_75t_L g578 ( .A(n_576), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g620 ( .A(n_576), .B(n_616), .Y(n_620) );
AND2x2_ASAP7_75t_L g735 ( .A(n_576), .B(n_633), .Y(n_735) );
AND2x2_ASAP7_75t_L g738 ( .A(n_576), .B(n_644), .Y(n_738) );
AND2x4_ASAP7_75t_L g746 ( .A(n_576), .B(n_747), .Y(n_746) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_578), .A2(n_701), .B(n_703), .Y(n_700) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g728 ( .A(n_580), .Y(n_728) );
AND2x2_ASAP7_75t_L g744 ( .A(n_580), .B(n_745), .Y(n_744) );
INVx4_ASAP7_75t_L g658 ( .A(n_582), .Y(n_658) );
INVx1_ASAP7_75t_L g627 ( .A(n_583), .Y(n_627) );
AND2x2_ASAP7_75t_L g649 ( .A(n_583), .B(n_602), .Y(n_649) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_608), .Y(n_584) );
OAI21xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B(n_594), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g595 ( .A(n_587), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_SL g748 ( .A(n_587), .B(n_600), .Y(n_748) );
AND2x2_ASAP7_75t_L g769 ( .A(n_587), .B(n_685), .Y(n_769) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g695 ( .A(n_592), .Y(n_695) );
OAI21xp5_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_597), .B(n_604), .Y(n_594) );
OR2x6_ASAP7_75t_L g647 ( .A(n_596), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_603), .Y(n_598) );
INVx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
OR2x2_ASAP7_75t_L g670 ( .A(n_605), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g767 ( .A(n_605), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_606), .B(n_740), .Y(n_739) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_621), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_612), .B1(n_618), .B2(n_620), .Y(n_609) );
OR2x2_ASAP7_75t_L g681 ( .A(n_611), .B(n_682), .Y(n_681) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_613), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g687 ( .A(n_616), .Y(n_687) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVxp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B1(n_630), .B2(n_632), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_628), .Y(n_624) );
AND2x4_ASAP7_75t_SL g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_628), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g691 ( .A(n_631), .B(n_685), .Y(n_691) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_636), .B(n_676), .Y(n_635) );
NOR2xp67_ASAP7_75t_L g636 ( .A(n_637), .B(n_650), .Y(n_636) );
AOI21xp33_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B(n_645), .Y(n_637) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2x1p5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI22xp33_ASAP7_75t_SL g715 ( .A1(n_647), .A2(n_716), .B1(n_718), .B2(n_721), .Y(n_715) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_648), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g698 ( .A(n_649), .B(n_699), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B(n_654), .C(n_664), .Y(n_650) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp33_ASAP7_75t_SL g655 ( .A(n_656), .B(n_658), .Y(n_655) );
INVxp33_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g667 ( .A(n_658), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_659), .A2(n_679), .B1(n_680), .B2(n_683), .C(n_686), .Y(n_678) );
AND2x4_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g719 ( .A(n_660), .Y(n_719) );
INVx2_ASAP7_75t_SL g717 ( .A(n_663), .Y(n_717) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NAND2x1_ASAP7_75t_L g716 ( .A(n_667), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g713 ( .A(n_673), .Y(n_713) );
INVx1_ASAP7_75t_L g742 ( .A(n_674), .Y(n_742) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_692), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_690), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g731 ( .A(n_682), .Y(n_731) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g752 ( .A(n_685), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g757 ( .A(n_685), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVxp33_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
BUFx2_ASAP7_75t_L g710 ( .A(n_689), .Y(n_710) );
OAI21xp5_ASAP7_75t_SL g692 ( .A1(n_693), .A2(n_697), .B(n_700), .Y(n_692) );
INVxp67_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
BUFx2_ASAP7_75t_L g753 ( .A(n_699), .Y(n_753) );
AND2x2_ASAP7_75t_L g741 ( .A(n_702), .B(n_742), .Y(n_741) );
NOR2xp33_ASAP7_75t_R g703 ( .A(n_704), .B(n_705), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_722), .C(n_749), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_715), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_709), .B(n_712), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
OR2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_736), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_724), .B(n_733), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g724 ( .A1(n_725), .A2(n_727), .B1(n_729), .B2(n_730), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NOR2x1_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVxp67_ASAP7_75t_SL g734 ( .A(n_732), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_737), .B(n_743), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_746), .B(n_748), .Y(n_743) );
INVx1_ASAP7_75t_L g762 ( .A(n_746), .Y(n_762) );
AOI211xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_752), .B(n_754), .C(n_763), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_758), .B1(n_760), .B2(n_762), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_768), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVxp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
INVx3_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_782), .B(n_788), .Y(n_781) );
INVxp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g783 ( .A(n_784), .B(n_787), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
OR2x2_ASAP7_75t_SL g805 ( .A(n_785), .B(n_787), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g807 ( .A1(n_785), .A2(n_808), .B(n_811), .Y(n_807) );
BUFx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
BUFx2_ASAP7_75t_L g795 ( .A(n_789), .Y(n_795) );
BUFx3_ASAP7_75t_L g800 ( .A(n_789), .Y(n_800) );
INVxp67_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_794), .B(n_796), .Y(n_791) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g811 ( .A(n_795), .Y(n_811) );
NOR2xp33_ASAP7_75t_SL g796 ( .A(n_797), .B(n_801), .Y(n_796) );
INVx1_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
BUFx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
CKINVDCx11_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
CKINVDCx8_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
endmodule