module fake_jpeg_17829_n_360 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_360);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_31),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_24),
.B(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_24),
.A2(n_45),
.B1(n_42),
.B2(n_37),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_37),
.B1(n_29),
.B2(n_47),
.Y(n_77)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_60),
.Y(n_79)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_21),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_68),
.Y(n_102)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_37),
.B1(n_29),
.B2(n_38),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_96),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_77),
.A2(n_47),
.B1(n_33),
.B2(n_43),
.Y(n_131)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_48),
.A2(n_29),
.B1(n_34),
.B2(n_27),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_63),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

BUFx2_ASAP7_75t_SL g155 ( 
.A(n_112),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_113),
.Y(n_163)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_116),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_118),
.B(n_129),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_130),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_51),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_68),
.B1(n_92),
.B2(n_85),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_70),
.B(n_60),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_80),
.B1(n_97),
.B2(n_95),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_147),
.B1(n_148),
.B2(n_121),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_33),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_23),
.C(n_35),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_151),
.B1(n_137),
.B2(n_154),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_52),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_156),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_131),
.A2(n_78),
.B1(n_49),
.B2(n_57),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_145),
.B1(n_123),
.B2(n_64),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_92),
.B1(n_61),
.B2(n_53),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_126),
.A2(n_85),
.B1(n_40),
.B2(n_43),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_102),
.A2(n_40),
.B1(n_43),
.B2(n_33),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_69),
.B1(n_53),
.B2(n_61),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_102),
.A2(n_33),
.B1(n_43),
.B2(n_27),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_153),
.A2(n_121),
.B1(n_81),
.B2(n_76),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_76),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_104),
.A2(n_21),
.B1(n_25),
.B2(n_22),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_108),
.B(n_35),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_109),
.Y(n_177)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_173),
.B1(n_178),
.B2(n_151),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_166),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_119),
.Y(n_166)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_167),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_159),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_SL g194 ( 
.A1(n_170),
.A2(n_178),
.B(n_155),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_103),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_152),
.B1(n_156),
.B2(n_134),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_141),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_179),
.Y(n_198)
);

OAI22x1_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_64),
.B1(n_122),
.B2(n_132),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_109),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_134),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_184),
.A2(n_186),
.B1(n_195),
.B2(n_199),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_183),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_171),
.B1(n_178),
.B2(n_175),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_176),
.C(n_146),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_175),
.B(n_136),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_188),
.Y(n_212)
);

AO21x1_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_187),
.B(n_179),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_180),
.B1(n_168),
.B2(n_165),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_169),
.A2(n_157),
.B1(n_152),
.B2(n_146),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_183),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_183),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_166),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_202),
.B(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_204),
.A2(n_208),
.B(n_144),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_171),
.B1(n_176),
.B2(n_181),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_210),
.B1(n_211),
.B2(n_184),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_201),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_221),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_212),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_199),
.A2(n_163),
.B1(n_170),
.B2(n_174),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_174),
.B1(n_143),
.B2(n_144),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_149),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_214),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_149),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_218),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_200),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_156),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_137),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_163),
.C(n_113),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_189),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_167),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_223),
.B(n_225),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_150),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_187),
.B1(n_192),
.B2(n_193),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_231),
.B1(n_241),
.B2(n_249),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_192),
.B1(n_200),
.B2(n_185),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_247),
.B(n_215),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_233),
.B(n_245),
.Y(n_260)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_145),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_239),
.C(n_240),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_189),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_210),
.A2(n_185),
.B1(n_163),
.B2(n_160),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_182),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_204),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_211),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_182),
.Y(n_245)
);

XOR2x2_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_88),
.Y(n_246)
);

XOR2x2_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_214),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_142),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_207),
.A2(n_142),
.B1(n_161),
.B2(n_139),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_204),
.B(n_206),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_251),
.A2(n_258),
.B(n_265),
.Y(n_272)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_267),
.Y(n_274)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_255),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_244),
.A2(n_224),
.B1(n_220),
.B2(n_205),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_259),
.B1(n_261),
.B2(n_231),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_257),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_248),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_246),
.A2(n_220),
.B1(n_213),
.B2(n_222),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

AOI21x1_ASAP7_75t_SL g290 ( 
.A1(n_266),
.A2(n_44),
.B(n_36),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_216),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_216),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_229),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_139),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_237),
.B1(n_25),
.B2(n_26),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_88),
.C(n_172),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_229),
.C(n_230),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_247),
.B1(n_243),
.B2(n_238),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_284),
.B1(n_285),
.B2(n_288),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_252),
.A2(n_247),
.B1(n_226),
.B2(n_241),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_276),
.A2(n_290),
.B1(n_251),
.B2(n_264),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_256),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_280),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_235),
.Y(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_172),
.C(n_158),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_283),
.B(n_287),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_26),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_158),
.B1(n_111),
.B2(n_115),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_271),
.C(n_261),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_259),
.A2(n_110),
.B1(n_39),
.B2(n_34),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_250),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_290),
.B1(n_277),
.B2(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_298),
.Y(n_309)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_297),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_276),
.A2(n_255),
.B1(n_260),
.B2(n_258),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_275),
.A2(n_286),
.B1(n_281),
.B2(n_253),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_304),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_306),
.C(n_44),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_289),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_302),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_262),
.Y(n_303)
);

OAI321xp33_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_288),
.A3(n_273),
.B1(n_285),
.B2(n_279),
.C(n_8),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_250),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_278),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_264),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_253),
.B1(n_269),
.B2(n_254),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_310),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_304),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_36),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_293),
.A2(n_41),
.B1(n_39),
.B2(n_44),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_315),
.C(n_316),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_295),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_36),
.C(n_30),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_296),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_294),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_6),
.Y(n_330)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_321),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_322),
.B(n_324),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_309),
.B(n_301),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_326),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_117),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_318),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_319),
.C(n_318),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_311),
.B(n_299),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_329),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_299),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_8),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_332),
.B(n_335),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_307),
.C(n_30),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_334),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_35),
.C(n_9),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_35),
.C(n_9),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_325),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_10),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_11),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_343),
.B(n_345),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_340),
.B(n_10),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_11),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_346),
.A2(n_348),
.B(n_12),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_347),
.A2(n_12),
.B(n_13),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_35),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_350),
.Y(n_354)
);

NAND4xp25_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_338),
.C(n_337),
.D(n_14),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_351),
.B(n_342),
.C(n_14),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_353),
.A2(n_354),
.B1(n_352),
.B2(n_16),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_355),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_13),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_17),
.C(n_15),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_15),
.C(n_16),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_15),
.Y(n_360)
);


endmodule