module fake_ibex_1353_n_1930 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_357, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_317, n_340, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_366, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_320, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_324, n_78, n_20, n_69, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1930);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_357;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_366;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1930;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1883;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_1922;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_1778;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_447;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_379;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1717;
wire n_1609;
wire n_391;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_737;
wire n_606;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_395;
wire n_1786;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_981;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_974;
wire n_1036;
wire n_1831;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_388;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1806;
wire n_1599;
wire n_650;
wire n_409;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_1925;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1894;
wire n_634;
wire n_961;
wire n_991;
wire n_1349;
wire n_1223;
wire n_1331;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_403;
wire n_1353;
wire n_423;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1830;
wire n_1629;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1899;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1839;
wire n_1617;
wire n_1587;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_804;
wire n_484;
wire n_1455;
wire n_1871;
wire n_1642;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_1767;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_1928;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1892;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1635;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1757;
wire n_699;
wire n_918;
wire n_1913;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_548;
wire n_1158;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_405;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_414;
wire n_378;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1900;
wire n_519;
wire n_1843;
wire n_408;
wire n_1665;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_394;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_344),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_115),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_36),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_198),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_257),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_356),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_298),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_372),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_312),
.Y(n_386)
);

BUFx10_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_19),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_79),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_189),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_255),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_238),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_18),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_291),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_200),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_277),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_101),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_51),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_253),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_300),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_212),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_313),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_352),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_370),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_225),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_147),
.B(n_152),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_315),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_210),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_112),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_0),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_292),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_103),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_282),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_267),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_116),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_322),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_124),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_287),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_4),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_135),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_373),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_371),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_26),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_244),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_317),
.Y(n_429)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_305),
.Y(n_430)
);

BUFx8_ASAP7_75t_SL g431 ( 
.A(n_186),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_87),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_193),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_116),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_316),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_165),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_358),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_241),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_326),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_206),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_107),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_323),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_365),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_307),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_157),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_350),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_239),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_20),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_328),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_355),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_362),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_124),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_219),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_51),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_351),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_348),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_93),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_91),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_179),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_231),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_304),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_109),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_217),
.Y(n_463)
);

INVxp33_ASAP7_75t_SL g464 ( 
.A(n_233),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_186),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_180),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_178),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_324),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_203),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_28),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_211),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_301),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_163),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_154),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_235),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_101),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_295),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_311),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_341),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_319),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_173),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_246),
.Y(n_482)
);

BUFx5_ASAP7_75t_L g483 ( 
.A(n_3),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_90),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_285),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_314),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_284),
.Y(n_487)
);

BUFx10_ASAP7_75t_L g488 ( 
.A(n_197),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_150),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_72),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_53),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_374),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_64),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_50),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_122),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_64),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_182),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_225),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_243),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_333),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_320),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_331),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_229),
.Y(n_503)
);

BUFx10_ASAP7_75t_L g504 ( 
.A(n_224),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_18),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_276),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_226),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_32),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_346),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_252),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_82),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_27),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_217),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_158),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_239),
.B(n_123),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_164),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_293),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_294),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_29),
.Y(n_519)
);

CKINVDCx14_ASAP7_75t_R g520 ( 
.A(n_330),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_229),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_274),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_183),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_349),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_288),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_241),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_363),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_179),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_134),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_78),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_143),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_369),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_335),
.Y(n_533)
);

BUFx2_ASAP7_75t_SL g534 ( 
.A(n_106),
.Y(n_534)
);

BUFx5_ASAP7_75t_L g535 ( 
.A(n_102),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_302),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_347),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_193),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_68),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_244),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_63),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_54),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_126),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_214),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_59),
.Y(n_545)
);

CKINVDCx14_ASAP7_75t_R g546 ( 
.A(n_127),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_149),
.Y(n_547)
);

BUFx5_ASAP7_75t_L g548 ( 
.A(n_268),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_367),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_46),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_223),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_357),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_190),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_62),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_318),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_218),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_30),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_150),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_56),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_139),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_142),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_281),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_297),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_137),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_238),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_209),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_240),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_366),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_250),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_204),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_272),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_266),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_233),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_104),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_342),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_0),
.Y(n_576)
);

CKINVDCx14_ASAP7_75t_R g577 ( 
.A(n_290),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_308),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_216),
.Y(n_579)
);

INVxp67_ASAP7_75t_SL g580 ( 
.A(n_21),
.Y(n_580)
);

NOR2xp67_ASAP7_75t_L g581 ( 
.A(n_103),
.B(n_156),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_214),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_309),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_345),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_209),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_136),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_110),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_235),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_176),
.Y(n_589)
);

INVxp67_ASAP7_75t_SL g590 ( 
.A(n_236),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_299),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_310),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_343),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_159),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_30),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_1),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_188),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_104),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_269),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_52),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_237),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_232),
.B(n_29),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_306),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_264),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_275),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_61),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_303),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_48),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_353),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_195),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_234),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_391),
.B(n_2),
.Y(n_612)
);

AND2x6_ASAP7_75t_L g613 ( 
.A(n_446),
.B(n_477),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_540),
.B(n_2),
.Y(n_614)
);

CKINVDCx6p67_ASAP7_75t_R g615 ( 
.A(n_410),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_391),
.B(n_5),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_546),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_446),
.B(n_251),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_418),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_483),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_589),
.B(n_382),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_483),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_483),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_391),
.B(n_6),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_491),
.B(n_7),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_548),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_544),
.B(n_8),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_546),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_464),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_483),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_483),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_548),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_387),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_544),
.B(n_9),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_418),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_387),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_418),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_548),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_418),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_380),
.A2(n_256),
.B(n_254),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_535),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_535),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_478),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_535),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_535),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_422),
.B(n_10),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_535),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_422),
.B(n_11),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_535),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_535),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_548),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_387),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_380),
.A2(n_259),
.B(n_258),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_413),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_548),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_450),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_610),
.B(n_11),
.Y(n_657)
);

BUFx8_ASAP7_75t_L g658 ( 
.A(n_548),
.Y(n_658)
);

OA21x2_ASAP7_75t_L g659 ( 
.A1(n_401),
.A2(n_455),
.B(n_442),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_411),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_500),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_430),
.B(n_12),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_500),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_413),
.B(n_13),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_464),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_665)
);

AND2x2_ASAP7_75t_SL g666 ( 
.A(n_449),
.B(n_260),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_376),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_419),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_548),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_401),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_536),
.Y(n_671)
);

AND2x6_ASAP7_75t_L g672 ( 
.A(n_477),
.B(n_261),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_500),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_419),
.Y(n_674)
);

OAI21x1_ASAP7_75t_L g675 ( 
.A1(n_442),
.A2(n_263),
.B(n_262),
.Y(n_675)
);

BUFx12f_ASAP7_75t_L g676 ( 
.A(n_536),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_421),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_421),
.B(n_16),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_430),
.B(n_17),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_455),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_539),
.Y(n_681)
);

OA21x2_ASAP7_75t_L g682 ( 
.A1(n_479),
.A2(n_270),
.B(n_265),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_432),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_479),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_500),
.Y(n_685)
);

CKINVDCx8_ASAP7_75t_R g686 ( 
.A(n_517),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_432),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_539),
.Y(n_688)
);

BUFx12f_ASAP7_75t_L g689 ( 
.A(n_488),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_539),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_527),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_599),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_SL g693 ( 
.A1(n_376),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_411),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_447),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_447),
.Y(n_696)
);

OA21x2_ASAP7_75t_L g697 ( 
.A1(n_522),
.A2(n_273),
.B(n_271),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_475),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_488),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_527),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_522),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_537),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_552),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_SL g704 ( 
.A1(n_378),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_527),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_412),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_552),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_656),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_664),
.A2(n_515),
.B1(n_389),
.B2(n_393),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_SL g710 ( 
.A(n_662),
.B(n_375),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_643),
.B(n_520),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_612),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_612),
.Y(n_713)
);

NOR2x1p5_ASAP7_75t_L g714 ( 
.A(n_689),
.B(n_676),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_612),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_613),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_643),
.B(n_520),
.Y(n_717)
);

XNOR2xp5_ASAP7_75t_L g718 ( 
.A(n_628),
.B(n_378),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_619),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_612),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_620),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_616),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_621),
.B(n_412),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_671),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_636),
.B(n_475),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_689),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_671),
.B(n_476),
.Y(n_727)
);

XOR2xp5_ASAP7_75t_L g728 ( 
.A(n_692),
.B(n_375),
.Y(n_728)
);

AND3x2_ASAP7_75t_L g729 ( 
.A(n_657),
.B(n_706),
.C(n_660),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_658),
.B(n_578),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_616),
.B(n_584),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_616),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_616),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_624),
.B(n_584),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_624),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_624),
.Y(n_736)
);

OAI22xp33_ASAP7_75t_L g737 ( 
.A1(n_629),
.A2(n_665),
.B1(n_694),
.B2(n_625),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_624),
.B(n_593),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_676),
.B(n_534),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_618),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_664),
.Y(n_741)
);

BUFx4f_ASAP7_75t_L g742 ( 
.A(n_615),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_622),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_622),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_636),
.B(n_476),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_613),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_615),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_623),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_619),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_623),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_636),
.B(n_481),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_652),
.B(n_481),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_699),
.B(n_652),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_L g754 ( 
.A(n_646),
.B(n_498),
.C(n_471),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_641),
.Y(n_755)
);

XNOR2xp5_ASAP7_75t_L g756 ( 
.A(n_666),
.B(n_390),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_662),
.Y(n_757)
);

INVx5_ASAP7_75t_L g758 ( 
.A(n_618),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_652),
.B(n_407),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_652),
.B(n_451),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_627),
.B(n_593),
.Y(n_761)
);

NAND2x1p5_ASAP7_75t_L g762 ( 
.A(n_679),
.B(n_377),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_678),
.Y(n_763)
);

OR2x6_ASAP7_75t_L g764 ( 
.A(n_625),
.B(n_409),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_644),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_627),
.B(n_379),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_678),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_679),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_627),
.B(n_381),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_618),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_659),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_678),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_657),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_659),
.Y(n_774)
);

AND3x2_ASAP7_75t_L g775 ( 
.A(n_646),
.B(n_580),
.C(n_459),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_678),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_633),
.B(n_484),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_627),
.B(n_484),
.Y(n_778)
);

BUFx4f_ASAP7_75t_L g779 ( 
.A(n_666),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_648),
.B(n_579),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_686),
.Y(n_781)
);

AND2x6_ASAP7_75t_L g782 ( 
.A(n_634),
.B(n_555),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_634),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_666),
.A2(n_399),
.B1(n_402),
.B2(n_394),
.Y(n_784)
);

AND3x2_ASAP7_75t_L g785 ( 
.A(n_634),
.B(n_590),
.C(n_431),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_634),
.B(n_654),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_654),
.B(n_489),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_626),
.Y(n_788)
);

BUFx10_ASAP7_75t_L g789 ( 
.A(n_613),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_619),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_630),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_670),
.Y(n_792)
);

INVx4_ASAP7_75t_L g793 ( 
.A(n_618),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_630),
.Y(n_794)
);

BUFx10_ASAP7_75t_L g795 ( 
.A(n_613),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_631),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_631),
.B(n_383),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_686),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_668),
.B(n_674),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_642),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_668),
.B(n_456),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_619),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_642),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_645),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_674),
.B(n_489),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_645),
.B(n_385),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_614),
.B(n_577),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_632),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_647),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_677),
.B(n_388),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_635),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_683),
.B(n_392),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_683),
.B(n_577),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_647),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_649),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_687),
.B(n_493),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_687),
.B(n_586),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_635),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_638),
.Y(n_819)
);

BUFx10_ASAP7_75t_L g820 ( 
.A(n_613),
.Y(n_820)
);

OAI22xp33_ASAP7_75t_L g821 ( 
.A1(n_629),
.A2(n_665),
.B1(n_694),
.B2(n_617),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_695),
.B(n_488),
.Y(n_822)
);

AND2x2_ASAP7_75t_SL g823 ( 
.A(n_682),
.B(n_602),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_638),
.Y(n_824)
);

AND2x6_ASAP7_75t_L g825 ( 
.A(n_638),
.B(n_555),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_618),
.Y(n_826)
);

AND2x6_ASAP7_75t_L g827 ( 
.A(n_651),
.B(n_562),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_695),
.B(n_395),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_651),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_649),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_650),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_672),
.B(n_607),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_655),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_650),
.B(n_397),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_655),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_613),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_696),
.B(n_698),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_655),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_680),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_635),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_672),
.A2(n_415),
.B1(n_423),
.B2(n_408),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_684),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_701),
.Y(n_843)
);

AND2x6_ASAP7_75t_L g844 ( 
.A(n_672),
.B(n_562),
.Y(n_844)
);

NAND2xp33_ASAP7_75t_L g845 ( 
.A(n_672),
.B(n_527),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_698),
.B(n_504),
.Y(n_846)
);

XNOR2xp5_ASAP7_75t_L g847 ( 
.A(n_667),
.B(n_390),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_672),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_669),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_702),
.B(n_493),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_702),
.B(n_405),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_L g852 ( 
.A(n_844),
.B(n_672),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_731),
.A2(n_738),
.B(n_734),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_813),
.B(n_404),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_807),
.B(n_406),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_727),
.B(n_406),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_784),
.A2(n_384),
.B1(n_425),
.B2(n_414),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_789),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_724),
.B(n_416),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_822),
.B(n_416),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_784),
.A2(n_425),
.B1(n_472),
.B2(n_414),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_739),
.B(n_472),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_846),
.B(n_386),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_779),
.A2(n_709),
.B1(n_723),
.B2(n_762),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_759),
.B(n_403),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_745),
.B(n_703),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_779),
.A2(n_707),
.B1(n_703),
.B2(n_428),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_782),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_711),
.B(n_504),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_725),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_759),
.B(n_437),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_726),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_760),
.B(n_751),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_752),
.B(n_707),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_717),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_725),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_742),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_782),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_731),
.A2(n_653),
.B(n_640),
.Y(n_879)
);

AND2x6_ASAP7_75t_SL g880 ( 
.A(n_739),
.B(n_693),
.Y(n_880)
);

AND2x2_ASAP7_75t_SL g881 ( 
.A(n_742),
.B(n_682),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_757),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_753),
.B(n_417),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_725),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_763),
.A2(n_438),
.B1(n_440),
.B2(n_434),
.Y(n_885)
);

OR2x6_ASAP7_75t_L g886 ( 
.A(n_739),
.B(n_704),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_780),
.B(n_468),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_786),
.B(n_487),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_786),
.B(n_492),
.Y(n_889)
);

BUFx6f_ASAP7_75t_SL g890 ( 
.A(n_708),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_712),
.A2(n_653),
.B(n_675),
.C(n_640),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_768),
.B(n_509),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_777),
.B(n_420),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_777),
.B(n_524),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_767),
.A2(n_445),
.B1(n_448),
.B2(n_441),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_754),
.A2(n_510),
.B1(n_572),
.B2(n_506),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_714),
.B(n_704),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_747),
.B(n_504),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_799),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_817),
.B(n_563),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_767),
.A2(n_457),
.B1(n_460),
.B2(n_452),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_737),
.A2(n_510),
.B1(n_572),
.B2(n_506),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_785),
.B(n_775),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_SL g904 ( 
.A1(n_810),
.A2(n_812),
.B(n_828),
.C(n_837),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_734),
.A2(n_738),
.B(n_766),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_708),
.B(n_554),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_708),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_778),
.B(n_603),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_781),
.B(n_554),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_778),
.B(n_604),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_776),
.A2(n_467),
.B1(n_473),
.B2(n_463),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_766),
.B(n_426),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_769),
.B(n_429),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_787),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_769),
.B(n_435),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_801),
.B(n_439),
.Y(n_916)
);

XNOR2xp5_ASAP7_75t_L g917 ( 
.A(n_756),
.B(n_433),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_801),
.B(n_400),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_741),
.B(n_480),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_715),
.A2(n_575),
.B1(n_396),
.B2(n_398),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_772),
.B(n_443),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_722),
.B(n_501),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_805),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_713),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_732),
.B(n_502),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_735),
.B(n_549),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_821),
.A2(n_575),
.B1(n_424),
.B2(n_427),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_740),
.B(n_770),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_798),
.B(n_681),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_736),
.B(n_720),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_720),
.B(n_733),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_761),
.B(n_444),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_783),
.A2(n_497),
.B1(n_499),
.B2(n_490),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_816),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_733),
.A2(n_507),
.B1(n_508),
.B2(n_505),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_816),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_789),
.Y(n_937)
);

BUFx12f_ASAP7_75t_L g938 ( 
.A(n_764),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_792),
.B(n_436),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_793),
.B(n_461),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_789),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_764),
.B(n_554),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_764),
.B(n_581),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_816),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_839),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_850),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_842),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_843),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_850),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_771),
.A2(n_514),
.B1(n_516),
.B2(n_513),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_774),
.A2(n_697),
.B(n_682),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_730),
.B(n_485),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_810),
.B(n_454),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_851),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_812),
.B(n_486),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_851),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_841),
.B(n_458),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_841),
.B(n_465),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_797),
.B(n_469),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_806),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_834),
.B(n_791),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_823),
.A2(n_528),
.B1(n_529),
.B2(n_526),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_823),
.A2(n_545),
.B1(n_547),
.B2(n_538),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_834),
.B(n_474),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_794),
.B(n_518),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_796),
.B(n_482),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_800),
.B(n_494),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_758),
.B(n_525),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_803),
.B(n_503),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_804),
.B(n_532),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_825),
.A2(n_551),
.B1(n_553),
.B2(n_550),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_809),
.B(n_511),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_729),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_718),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_814),
.B(n_533),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_815),
.B(n_830),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_795),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_831),
.B(n_512),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_825),
.Y(n_979)
);

NOR3xp33_ASAP7_75t_L g980 ( 
.A(n_710),
.B(n_594),
.C(n_523),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_827),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_832),
.A2(n_559),
.B(n_560),
.C(n_558),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_788),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_827),
.B(n_519),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_827),
.A2(n_564),
.B1(n_566),
.B2(n_561),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_827),
.A2(n_573),
.B1(n_574),
.B2(n_569),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_728),
.B(n_611),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_847),
.B(n_611),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_SL g989 ( 
.A(n_826),
.B(n_433),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_827),
.A2(n_585),
.B1(n_588),
.B2(n_582),
.Y(n_990)
);

NOR2x2_ASAP7_75t_L g991 ( 
.A(n_710),
.B(n_453),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_808),
.B(n_541),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_819),
.B(n_542),
.Y(n_993)
);

INVxp67_ASAP7_75t_SL g994 ( 
.A(n_848),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_832),
.A2(n_596),
.B1(n_597),
.B2(n_595),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_716),
.B(n_521),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_716),
.B(n_568),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_824),
.B(n_543),
.Y(n_998)
);

AND2x6_ASAP7_75t_SL g999 ( 
.A(n_845),
.B(n_600),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_845),
.A2(n_565),
.B1(n_567),
.B2(n_557),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_849),
.Y(n_1001)
);

INVx8_ASAP7_75t_L g1002 ( 
.A(n_746),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_849),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_829),
.B(n_598),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_746),
.B(n_583),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_795),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_829),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_833),
.B(n_601),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_833),
.B(n_606),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_836),
.B(n_591),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_835),
.B(n_608),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_835),
.B(n_592),
.Y(n_1012)
);

INVx8_ASAP7_75t_L g1013 ( 
.A(n_820),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_838),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_721),
.B(n_605),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_719),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_721),
.B(n_462),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_909),
.B(n_882),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_868),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_899),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_872),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_1017),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_882),
.B(n_462),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_989),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_862),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_951),
.A2(n_744),
.B(n_743),
.Y(n_1026)
);

INVx5_ASAP7_75t_L g1027 ( 
.A(n_878),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_853),
.A2(n_748),
.B(n_750),
.C(n_744),
.Y(n_1028)
);

OAI22x1_ASAP7_75t_L g1029 ( 
.A1(n_902),
.A2(n_470),
.B1(n_495),
.B2(n_466),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_862),
.B(n_466),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_890),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_931),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_875),
.B(n_470),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_890),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_873),
.B(n_755),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_857),
.B(n_495),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_962),
.A2(n_496),
.B1(n_531),
.B2(n_530),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_928),
.A2(n_765),
.B(n_697),
.Y(n_1038)
);

AO22x1_ASAP7_75t_L g1039 ( 
.A1(n_907),
.A2(n_496),
.B1(n_531),
.B2(n_530),
.Y(n_1039)
);

INVx5_ASAP7_75t_L g1040 ( 
.A(n_996),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_869),
.B(n_864),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_962),
.A2(n_570),
.B1(n_587),
.B2(n_556),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_963),
.A2(n_539),
.B1(n_576),
.B2(n_681),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_924),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_870),
.Y(n_1045)
);

OAI21xp33_ASAP7_75t_SL g1046 ( 
.A1(n_963),
.A2(n_691),
.B(n_685),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_L g1047 ( 
.A(n_980),
.B(n_576),
.C(n_571),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_945),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_950),
.A2(n_690),
.B1(n_688),
.B2(n_691),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_947),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_948),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_R g1052 ( 
.A(n_974),
.B(n_31),
.Y(n_1052)
);

NOR2xp67_ASAP7_75t_L g1053 ( 
.A(n_973),
.B(n_33),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_860),
.B(n_34),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_927),
.B(n_35),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_L g1056 ( 
.A(n_938),
.B(n_36),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_877),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_876),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_988),
.B(n_37),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_884),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_930),
.A2(n_705),
.B(n_39),
.C(n_37),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_914),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_898),
.B(n_38),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_903),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_SL g1065 ( 
.A(n_987),
.B(n_38),
.C(n_39),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_906),
.B(n_896),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_942),
.B(n_40),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_867),
.A2(n_609),
.B1(n_607),
.B2(n_635),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_905),
.A2(n_609),
.B(n_637),
.C(n_635),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_920),
.B(n_41),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_1008),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_976),
.B(n_609),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_996),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_883),
.B(n_41),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_961),
.A2(n_639),
.B(n_661),
.C(n_637),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_855),
.B(n_42),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_883),
.A2(n_952),
.B1(n_958),
.B2(n_957),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_863),
.B(n_42),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_881),
.A2(n_790),
.B(n_749),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_854),
.B(n_43),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_881),
.A2(n_790),
.B(n_749),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_982),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_SL g1083 ( 
.A1(n_893),
.A2(n_802),
.B(n_811),
.C(n_790),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_929),
.B(n_44),
.Y(n_1084)
);

AND2x2_ASAP7_75t_SL g1085 ( 
.A(n_903),
.B(n_45),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_892),
.B(n_47),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_918),
.B(n_47),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_935),
.B(n_48),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_943),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_893),
.A2(n_912),
.B1(n_915),
.B2(n_913),
.Y(n_1090)
);

INVx4_ASAP7_75t_L g1091 ( 
.A(n_996),
.Y(n_1091)
);

NOR2xp67_ASAP7_75t_L g1092 ( 
.A(n_939),
.B(n_49),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_961),
.A2(n_811),
.B(n_802),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_953),
.A2(n_53),
.B(n_50),
.C(n_52),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_887),
.B(n_54),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_991),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_923),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_940),
.A2(n_840),
.B(n_818),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_880),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_866),
.A2(n_673),
.B(n_700),
.C(n_663),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_SL g1101 ( 
.A(n_886),
.B(n_673),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_886),
.B(n_55),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_916),
.B(n_56),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_966),
.B(n_57),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_960),
.A2(n_279),
.B(n_278),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_935),
.B(n_58),
.Y(n_1106)
);

AO21x1_ASAP7_75t_L g1107 ( 
.A1(n_955),
.A2(n_58),
.B(n_59),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_856),
.A2(n_283),
.B(n_280),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_934),
.B(n_60),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_994),
.A2(n_289),
.B(n_286),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_R g1111 ( 
.A(n_999),
.B(n_61),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_SL g1112 ( 
.A(n_886),
.B(n_897),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_967),
.B(n_62),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_1002),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_969),
.B(n_65),
.Y(n_1115)
);

BUFx2_ASAP7_75t_SL g1116 ( 
.A(n_979),
.Y(n_1116)
);

NOR2x1_ASAP7_75t_SL g1117 ( 
.A(n_981),
.B(n_66),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_897),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_897),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_936),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_1002),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_885),
.B(n_67),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_874),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_972),
.B(n_71),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_944),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_978),
.B(n_72),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_888),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_885),
.B(n_73),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_946),
.Y(n_1129)
);

INVx5_ASAP7_75t_L g1130 ( 
.A(n_1002),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_895),
.B(n_73),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_874),
.A2(n_932),
.B(n_913),
.C(n_915),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_943),
.B(n_74),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_900),
.A2(n_325),
.B(n_321),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_908),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_949),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_895),
.B(n_75),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_922),
.A2(n_329),
.B(n_327),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_889),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_925),
.A2(n_334),
.B(n_332),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_933),
.B(n_901),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_926),
.A2(n_338),
.B(n_337),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_917),
.B(n_76),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_901),
.B(n_76),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_911),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_919),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_894),
.B(n_80),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_955),
.A2(n_81),
.B(n_83),
.C(n_84),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_932),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_1149)
);

CKINVDCx10_ASAP7_75t_R g1150 ( 
.A(n_1000),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_1014),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_965),
.A2(n_88),
.B(n_89),
.C(n_90),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_910),
.A2(n_89),
.B(n_91),
.C(n_92),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1001),
.A2(n_364),
.B(n_361),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_859),
.Y(n_1155)
);

OR2x6_ASAP7_75t_SL g1156 ( 
.A(n_959),
.B(n_94),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_971),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_1157)
);

INVx5_ASAP7_75t_L g1158 ( 
.A(n_1013),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_992),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1003),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_964),
.B(n_95),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_921),
.B(n_96),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_965),
.B(n_970),
.Y(n_1163)
);

BUFx12f_ASAP7_75t_L g1164 ( 
.A(n_1016),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_993),
.Y(n_1165)
);

CKINVDCx11_ASAP7_75t_R g1166 ( 
.A(n_954),
.Y(n_1166)
);

OR2x6_ASAP7_75t_SL g1167 ( 
.A(n_865),
.B(n_871),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_971),
.B(n_97),
.C(n_98),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_985),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_970),
.B(n_99),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_975),
.B(n_100),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_975),
.B(n_102),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_921),
.B(n_105),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_985),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_1174)
);

INVx3_ASAP7_75t_SL g1175 ( 
.A(n_1016),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_SL g1176 ( 
.A(n_1013),
.B(n_108),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_956),
.B(n_108),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_998),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1004),
.A2(n_1009),
.B1(n_1011),
.B2(n_984),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_983),
.B(n_111),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_986),
.B(n_113),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_1013),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1015),
.B(n_114),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_990),
.B(n_117),
.Y(n_1184)
);

AO21x1_ASAP7_75t_L g1185 ( 
.A1(n_1012),
.A2(n_117),
.B(n_118),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1007),
.B(n_119),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_968),
.B(n_119),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_997),
.A2(n_120),
.B(n_121),
.C(n_122),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_997),
.A2(n_120),
.B(n_121),
.C(n_123),
.Y(n_1189)
);

AND2x6_ASAP7_75t_L g1190 ( 
.A(n_858),
.B(n_937),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1005),
.A2(n_125),
.B(n_126),
.C(n_127),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_995),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1010),
.B(n_130),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1022),
.B(n_131),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1031),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1020),
.B(n_131),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_1069),
.A2(n_132),
.A3(n_133),
.B(n_134),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1144),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1107),
.A2(n_133),
.A3(n_135),
.B(n_136),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1071),
.B(n_137),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1163),
.B(n_1006),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1185),
.A2(n_138),
.A3(n_139),
.B(n_140),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1090),
.B(n_138),
.Y(n_1203)
);

CKINVDCx11_ASAP7_75t_R g1204 ( 
.A(n_1031),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1021),
.Y(n_1205)
);

NOR2xp67_ASAP7_75t_L g1206 ( 
.A(n_1034),
.B(n_140),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1144),
.A2(n_941),
.B1(n_977),
.B2(n_143),
.Y(n_1207)
);

INVxp67_ASAP7_75t_SL g1208 ( 
.A(n_1037),
.Y(n_1208)
);

BUFx2_ASAP7_75t_R g1209 ( 
.A(n_1156),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1164),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1035),
.A2(n_941),
.B1(n_142),
.B2(n_144),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_1052),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1075),
.A2(n_141),
.A3(n_144),
.B(n_145),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1035),
.A2(n_141),
.B1(n_145),
.B2(n_146),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1175),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_1151),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1077),
.B(n_148),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1064),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1100),
.A2(n_151),
.A3(n_153),
.B(n_154),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1109),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1093),
.A2(n_153),
.B(n_155),
.Y(n_1221)
);

AOI221xp5_ASAP7_75t_L g1222 ( 
.A1(n_1042),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.C(n_158),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1028),
.A2(n_159),
.B(n_160),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1048),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1103),
.A2(n_161),
.B(n_162),
.C(n_163),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1025),
.B(n_162),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_1040),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_1040),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1068),
.A2(n_1043),
.A3(n_1072),
.B(n_1173),
.Y(n_1229)
);

AND2x6_ASAP7_75t_L g1230 ( 
.A(n_1114),
.B(n_165),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1050),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1039),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1051),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1023),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1068),
.A2(n_166),
.A3(n_167),
.B(n_168),
.Y(n_1235)
);

AO32x2_ASAP7_75t_L g1236 ( 
.A1(n_1043),
.A2(n_166),
.A3(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_1236)
);

NAND2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1130),
.B(n_169),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1072),
.A2(n_172),
.A3(n_173),
.B(n_174),
.Y(n_1238)
);

NAND3xp33_ASAP7_75t_L g1239 ( 
.A(n_1179),
.B(n_174),
.C(n_175),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1160),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1178),
.B(n_177),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_SL g1242 ( 
.A1(n_1177),
.A2(n_177),
.B(n_178),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1030),
.B(n_181),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1042),
.B(n_181),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1018),
.B(n_182),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1091),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1033),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1182),
.B(n_185),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1088),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1114),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1074),
.A2(n_1173),
.B1(n_1170),
.B2(n_1172),
.Y(n_1251)
);

AO32x2_ASAP7_75t_L g1252 ( 
.A1(n_1157),
.A2(n_190),
.A3(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1171),
.A2(n_1172),
.A3(n_1123),
.B(n_1110),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1046),
.A2(n_194),
.B(n_195),
.Y(n_1254)
);

INVx3_ASAP7_75t_SL g1255 ( 
.A(n_1085),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1036),
.B(n_196),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1066),
.B(n_199),
.Y(n_1257)
);

NAND2x2_ASAP7_75t_L g1258 ( 
.A(n_1143),
.B(n_1055),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1159),
.B(n_201),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1182),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1167),
.B(n_201),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1106),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1032),
.B(n_202),
.Y(n_1263)
);

INVx8_ASAP7_75t_L g1264 ( 
.A(n_1130),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1135),
.B(n_202),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1106),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1165),
.B(n_203),
.Y(n_1267)
);

BUFx10_ASAP7_75t_L g1268 ( 
.A(n_1177),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1127),
.B(n_1139),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1044),
.Y(n_1270)
);

OAI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1112),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1162),
.A2(n_207),
.B1(n_208),
.B2(n_210),
.Y(n_1272)
);

NOR2x1_ASAP7_75t_R g1273 ( 
.A(n_1118),
.B(n_211),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1089),
.B(n_213),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1130),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1091),
.Y(n_1276)
);

AO21x1_ASAP7_75t_L g1277 ( 
.A1(n_1154),
.A2(n_215),
.B(n_216),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1122),
.Y(n_1278)
);

OAI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1029),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_1279)
);

AOI21xp33_ASAP7_75t_L g1280 ( 
.A1(n_1193),
.A2(n_1061),
.B(n_1153),
.Y(n_1280)
);

O2A1O1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1148),
.A2(n_222),
.B(n_223),
.C(n_224),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1188),
.A2(n_227),
.A3(n_228),
.B(n_230),
.Y(n_1282)
);

NAND3x1_ASAP7_75t_L g1283 ( 
.A(n_1102),
.B(n_230),
.C(n_231),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1122),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1087),
.A2(n_232),
.B(n_234),
.C(n_236),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1062),
.B(n_237),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1128),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1128),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1131),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1027),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1131),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1097),
.B(n_242),
.Y(n_1292)
);

INVx4_ASAP7_75t_L g1293 ( 
.A(n_1027),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_SL g1294 ( 
.A(n_1176),
.B(n_245),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1145),
.A2(n_245),
.B(n_247),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1059),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1155),
.B(n_248),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1070),
.A2(n_249),
.B1(n_1096),
.B2(n_1184),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1166),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1098),
.A2(n_1080),
.B(n_1083),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1120),
.B(n_1125),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1137),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1129),
.B(n_1136),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1057),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1119),
.B(n_1024),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1057),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1189),
.A2(n_1191),
.A3(n_1152),
.B(n_1149),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1108),
.A2(n_1134),
.A3(n_1117),
.B(n_1186),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1095),
.A2(n_1104),
.B(n_1115),
.C(n_1124),
.Y(n_1309)
);

AO21x2_ASAP7_75t_L g1310 ( 
.A1(n_1180),
.A2(n_1138),
.B(n_1142),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1045),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1058),
.B(n_1060),
.Y(n_1312)
);

NAND2xp33_ASAP7_75t_SL g1313 ( 
.A(n_1019),
.B(n_1073),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1101),
.A2(n_1067),
.B1(n_1063),
.B2(n_1065),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1027),
.B(n_1121),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1140),
.A2(n_1169),
.A3(n_1157),
.B(n_1174),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1183),
.Y(n_1317)
);

BUFx4f_ASAP7_75t_SL g1318 ( 
.A(n_1133),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1113),
.A2(n_1126),
.B(n_1076),
.C(n_1054),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1150),
.Y(n_1320)
);

INVx6_ASAP7_75t_SL g1321 ( 
.A(n_1084),
.Y(n_1321)
);

NOR2xp67_ASAP7_75t_L g1322 ( 
.A(n_1099),
.B(n_1056),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1169),
.A2(n_1174),
.A3(n_1192),
.B(n_1105),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1078),
.A2(n_1161),
.B(n_1147),
.C(n_1086),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1053),
.A2(n_1168),
.B1(n_1092),
.B2(n_1181),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1111),
.Y(n_1326)
);

AO32x2_ASAP7_75t_L g1327 ( 
.A1(n_1049),
.A2(n_1094),
.A3(n_1146),
.B1(n_1082),
.B2(n_1047),
.Y(n_1327)
);

BUFx12f_ASAP7_75t_L g1328 ( 
.A(n_1187),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1116),
.Y(n_1329)
);

INVx5_ASAP7_75t_L g1330 ( 
.A(n_1190),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1190),
.A2(n_852),
.B(n_1038),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1022),
.B(n_773),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1037),
.A2(n_756),
.B1(n_902),
.B2(n_861),
.Y(n_1333)
);

OR2x6_ASAP7_75t_L g1334 ( 
.A(n_1182),
.B(n_862),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1020),
.B(n_1141),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1144),
.A2(n_779),
.B1(n_1041),
.B2(n_784),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1020),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1026),
.A2(n_879),
.B(n_891),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1164),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1034),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1175),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1020),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1020),
.B(n_1141),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1025),
.B(n_862),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1021),
.Y(n_1345)
);

AO32x2_ASAP7_75t_L g1346 ( 
.A1(n_1043),
.A2(n_1068),
.A3(n_1174),
.B1(n_1169),
.B2(n_1157),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_SL g1347 ( 
.A1(n_1085),
.A2(n_886),
.B1(n_897),
.B2(n_756),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_1034),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1020),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1025),
.B(n_862),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1041),
.A2(n_1163),
.B(n_1132),
.C(n_1103),
.Y(n_1351)
);

AOI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1079),
.A2(n_879),
.B(n_1081),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1041),
.A2(n_1163),
.B(n_1132),
.C(n_1103),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1020),
.B(n_1158),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1141),
.A2(n_779),
.B1(n_1144),
.B2(n_886),
.Y(n_1355)
);

CKINVDCx16_ASAP7_75t_R g1356 ( 
.A(n_1031),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1020),
.B(n_1141),
.Y(n_1357)
);

BUFx8_ASAP7_75t_SL g1358 ( 
.A(n_1034),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1158),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1022),
.B(n_773),
.Y(n_1360)
);

AO22x2_ASAP7_75t_L g1361 ( 
.A1(n_1037),
.A2(n_1042),
.B1(n_1144),
.B2(n_1109),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1164),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1020),
.B(n_1141),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1020),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1132),
.A2(n_904),
.B(n_1163),
.C(n_1074),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1020),
.B(n_1141),
.Y(n_1366)
);

INVx4_ASAP7_75t_L g1367 ( 
.A(n_1130),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1020),
.Y(n_1368)
);

BUFx12f_ASAP7_75t_L g1369 ( 
.A(n_1031),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1037),
.A2(n_756),
.B1(n_902),
.B2(n_861),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1141),
.A2(n_779),
.B1(n_1144),
.B2(n_886),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1020),
.B(n_1141),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1021),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1158),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1037),
.A2(n_902),
.B1(n_857),
.B2(n_861),
.Y(n_1375)
);

CKINVDCx8_ASAP7_75t_R g1376 ( 
.A(n_1034),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1164),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1041),
.A2(n_1163),
.B(n_1132),
.C(n_1103),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1158),
.B(n_1130),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1041),
.A2(n_1163),
.B(n_1132),
.C(n_1103),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1041),
.A2(n_1163),
.B(n_1132),
.C(n_1103),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1144),
.A2(n_779),
.B1(n_1041),
.B2(n_784),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1022),
.B(n_773),
.Y(n_1383)
);

AO31x2_ASAP7_75t_L g1384 ( 
.A1(n_1069),
.A2(n_891),
.A3(n_1107),
.B(n_1185),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1022),
.B(n_773),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1020),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1175),
.Y(n_1387)
);

INVx5_ASAP7_75t_SL g1388 ( 
.A(n_1114),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1026),
.A2(n_879),
.B(n_891),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1037),
.B(n_1042),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1037),
.A2(n_756),
.B1(n_902),
.B2(n_861),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1020),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1025),
.B(n_862),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1020),
.B(n_1141),
.Y(n_1394)
);

INVx6_ASAP7_75t_L g1395 ( 
.A(n_1031),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1144),
.A2(n_779),
.B1(n_1041),
.B2(n_784),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1132),
.A2(n_904),
.B(n_1163),
.C(n_1074),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1034),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1026),
.A2(n_879),
.B(n_891),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1031),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1020),
.B(n_1141),
.Y(n_1401)
);

AO21x2_ASAP7_75t_L g1402 ( 
.A1(n_1338),
.A2(n_1399),
.B(n_1389),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1269),
.B(n_1390),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1337),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1208),
.B(n_1375),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1341),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1392),
.Y(n_1407)
);

AOI21xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1255),
.A2(n_1347),
.B(n_1320),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1342),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1333),
.B(n_1370),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1264),
.Y(n_1411)
);

AO31x2_ASAP7_75t_L g1412 ( 
.A1(n_1277),
.A2(n_1251),
.A3(n_1353),
.B(n_1351),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1349),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1341),
.Y(n_1414)
);

CKINVDCx6p67_ASAP7_75t_R g1415 ( 
.A(n_1204),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1378),
.A2(n_1381),
.B(n_1380),
.Y(n_1416)
);

NAND3xp33_ASAP7_75t_L g1417 ( 
.A(n_1309),
.B(n_1324),
.C(n_1319),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1361),
.A2(n_1347),
.B1(n_1382),
.B2(n_1336),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1264),
.Y(n_1419)
);

INVx5_ASAP7_75t_L g1420 ( 
.A(n_1264),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1207),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1358),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1364),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1368),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1332),
.B(n_1360),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1386),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1361),
.B(n_1355),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1207),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1311),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1286),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1216),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1216),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1286),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1237),
.A2(n_1382),
.B(n_1336),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1371),
.A2(n_1396),
.B1(n_1198),
.B2(n_1391),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_SL g1436 ( 
.A1(n_1254),
.A2(n_1295),
.B(n_1223),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1223),
.A2(n_1254),
.B(n_1221),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1383),
.B(n_1385),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1215),
.Y(n_1439)
);

BUFx4f_ASAP7_75t_SL g1440 ( 
.A(n_1195),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1297),
.B(n_1256),
.Y(n_1441)
);

AO22x2_ASAP7_75t_L g1442 ( 
.A1(n_1396),
.A2(n_1295),
.B1(n_1239),
.B2(n_1244),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1357),
.B(n_1335),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1240),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1359),
.B(n_1374),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1330),
.B(n_1294),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1292),
.Y(n_1447)
);

AOI21xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1356),
.A2(n_1279),
.B(n_1232),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1292),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1258),
.A2(n_1350),
.B1(n_1393),
.B2(n_1344),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1310),
.A2(n_1280),
.B(n_1201),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_SL g1452 ( 
.A(n_1367),
.B(n_1330),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1224),
.Y(n_1453)
);

CKINVDCx11_ASAP7_75t_R g1454 ( 
.A(n_1376),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1233),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1196),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1241),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1354),
.B(n_1260),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1231),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1312),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1312),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1343),
.B(n_1363),
.Y(n_1462)
);

AOI21xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1261),
.A2(n_1398),
.B(n_1340),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1275),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1249),
.A2(n_1266),
.B(n_1262),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1354),
.B(n_1260),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1278),
.A2(n_1287),
.B(n_1284),
.Y(n_1467)
);

AO31x2_ASAP7_75t_L g1468 ( 
.A1(n_1288),
.A2(n_1289),
.A3(n_1291),
.B(n_1302),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1270),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1334),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1400),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1234),
.B(n_1328),
.Y(n_1472)
);

AND2x4_ASAP7_75t_SL g1473 ( 
.A(n_1334),
.B(n_1248),
.Y(n_1473)
);

NOR2x1_ASAP7_75t_SL g1474 ( 
.A(n_1330),
.B(n_1379),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1317),
.B(n_1220),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1366),
.B(n_1372),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1394),
.B(n_1401),
.Y(n_1477)
);

A2O1A1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1281),
.A2(n_1222),
.B(n_1217),
.C(n_1257),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_1348),
.Y(n_1479)
);

BUFx12f_ASAP7_75t_L g1480 ( 
.A(n_1369),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1301),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1325),
.A2(n_1203),
.B(n_1263),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1245),
.B(n_1298),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1297),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1294),
.B(n_1314),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1211),
.A2(n_1248),
.B(n_1214),
.Y(n_1486)
);

AO31x2_ASAP7_75t_L g1487 ( 
.A1(n_1211),
.A2(n_1214),
.A3(n_1272),
.B(n_1225),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1373),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1339),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1321),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1321),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1303),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1194),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1243),
.B(n_1200),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1267),
.B(n_1259),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1387),
.B(n_1205),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1265),
.B(n_1387),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1227),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1268),
.B(n_1226),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1272),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1268),
.B(n_1345),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1285),
.B(n_1247),
.C(n_1296),
.Y(n_1502)
);

NAND2x1p5_ASAP7_75t_L g1503 ( 
.A(n_1227),
.B(n_1228),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1274),
.B(n_1388),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1384),
.A2(n_1253),
.B(n_1229),
.Y(n_1505)
);

AO31x2_ASAP7_75t_L g1506 ( 
.A1(n_1384),
.A2(n_1229),
.A3(n_1253),
.B(n_1346),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_SL g1507 ( 
.A1(n_1290),
.A2(n_1293),
.B(n_1304),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1315),
.A2(n_1242),
.B(n_1228),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1388),
.B(n_1276),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1318),
.B(n_1305),
.Y(n_1510)
);

A2O1A1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1206),
.A2(n_1322),
.B(n_1346),
.C(n_1313),
.Y(n_1511)
);

NAND2x1p5_ASAP7_75t_L g1512 ( 
.A(n_1250),
.B(n_1246),
.Y(n_1512)
);

AOI222xp33_ASAP7_75t_L g1513 ( 
.A1(n_1273),
.A2(n_1326),
.B1(n_1299),
.B2(n_1212),
.C1(n_1209),
.C2(n_1271),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1308),
.A2(n_1202),
.B(n_1199),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1202),
.A2(n_1199),
.B(n_1316),
.Y(n_1515)
);

BUFx10_ASAP7_75t_L g1516 ( 
.A(n_1230),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1283),
.A2(n_1388),
.B1(n_1346),
.B2(n_1329),
.Y(n_1517)
);

AO21x2_ASAP7_75t_L g1518 ( 
.A1(n_1316),
.A2(n_1323),
.B(n_1327),
.Y(n_1518)
);

AO31x2_ASAP7_75t_L g1519 ( 
.A1(n_1199),
.A2(n_1323),
.A3(n_1282),
.B(n_1197),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1306),
.B(n_1210),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_L g1521 ( 
.A(n_1230),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1230),
.A2(n_1218),
.B1(n_1395),
.B2(n_1377),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1230),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1362),
.B(n_1307),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1252),
.A2(n_1307),
.B(n_1282),
.C(n_1236),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1213),
.A2(n_1197),
.B(n_1219),
.Y(n_1526)
);

A2O1A1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1252),
.A2(n_1236),
.B(n_1235),
.C(n_1197),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1235),
.Y(n_1528)
);

OA21x2_ASAP7_75t_L g1529 ( 
.A1(n_1213),
.A2(n_1238),
.B(n_1235),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1236),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1207),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1269),
.B(n_1037),
.Y(n_1532)
);

A2O1A1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1365),
.A2(n_1397),
.B(n_1295),
.C(n_1353),
.Y(n_1533)
);

AOI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1352),
.A2(n_1300),
.B(n_1331),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1208),
.B(n_1141),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1264),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1264),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1354),
.B(n_1260),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1207),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1337),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1341),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1375),
.B(n_1390),
.Y(n_1542)
);

AO31x2_ASAP7_75t_L g1543 ( 
.A1(n_1277),
.A2(n_1251),
.A3(n_1353),
.B(n_1351),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1361),
.A2(n_1042),
.B1(n_1037),
.B2(n_1347),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1264),
.Y(n_1545)
);

AO21x2_ASAP7_75t_L g1546 ( 
.A1(n_1338),
.A2(n_1399),
.B(n_1389),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1338),
.A2(n_1399),
.B(n_1389),
.Y(n_1547)
);

AO21x2_ASAP7_75t_L g1548 ( 
.A1(n_1338),
.A2(n_1399),
.B(n_1389),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1337),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1390),
.B(n_1332),
.Y(n_1550)
);

INVx6_ASAP7_75t_L g1551 ( 
.A(n_1264),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1361),
.A2(n_1390),
.B1(n_1085),
.B2(n_1347),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1208),
.B(n_1141),
.Y(n_1553)
);

OR2x6_ASAP7_75t_L g1554 ( 
.A(n_1264),
.B(n_1334),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1467),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1410),
.B(n_1550),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1460),
.B(n_1461),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1410),
.B(n_1532),
.Y(n_1558)
);

AO21x1_ASAP7_75t_SL g1559 ( 
.A1(n_1421),
.A2(n_1531),
.B(n_1428),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1521),
.A2(n_1446),
.B(n_1437),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1450),
.B(n_1484),
.Y(n_1561)
);

AO31x2_ASAP7_75t_L g1562 ( 
.A1(n_1525),
.A2(n_1533),
.A3(n_1527),
.B(n_1451),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1409),
.Y(n_1563)
);

INVxp67_ASAP7_75t_SL g1564 ( 
.A(n_1473),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1444),
.B(n_1418),
.Y(n_1565)
);

INVx4_ASAP7_75t_SL g1566 ( 
.A(n_1521),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1444),
.B(n_1418),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1403),
.B(n_1427),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1481),
.B(n_1492),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1413),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1420),
.B(n_1473),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1423),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1484),
.B(n_1472),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1424),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1552),
.A2(n_1542),
.B1(n_1435),
.B2(n_1544),
.Y(n_1575)
);

AOI221xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1448),
.A2(n_1408),
.B1(n_1517),
.B2(n_1483),
.C(n_1416),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1426),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1488),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1478),
.A2(n_1502),
.B(n_1482),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1420),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1488),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1425),
.B(n_1438),
.Y(n_1582)
);

INVx4_ASAP7_75t_L g1583 ( 
.A(n_1420),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1429),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1464),
.Y(n_1585)
);

INVx3_ASAP7_75t_L g1586 ( 
.A(n_1420),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1468),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1468),
.Y(n_1588)
);

AO21x2_ASAP7_75t_L g1589 ( 
.A1(n_1534),
.A2(n_1533),
.B(n_1436),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1468),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1554),
.B(n_1523),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1472),
.B(n_1441),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1496),
.Y(n_1593)
);

INVx8_ASAP7_75t_L g1594 ( 
.A(n_1554),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1431),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1551),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1552),
.B(n_1404),
.Y(n_1597)
);

BUFx4f_ASAP7_75t_SL g1598 ( 
.A(n_1480),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1551),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1407),
.B(n_1540),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1431),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1462),
.B(n_1476),
.Y(n_1602)
);

INVxp33_ASAP7_75t_L g1603 ( 
.A(n_1419),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1549),
.B(n_1459),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1536),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1536),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1432),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1469),
.B(n_1443),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1405),
.B(n_1524),
.Y(n_1609)
);

INVxp67_ASAP7_75t_SL g1610 ( 
.A(n_1464),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1551),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1453),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1439),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1417),
.A2(n_1486),
.B(n_1482),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1535),
.B(n_1553),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1455),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1516),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1430),
.B(n_1433),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1406),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1414),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1477),
.B(n_1500),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1489),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1528),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1541),
.B(n_1499),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1516),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1411),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1554),
.B(n_1523),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1447),
.B(n_1449),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1475),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1475),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_1537),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1498),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1457),
.B(n_1456),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1530),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1442),
.B(n_1412),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1442),
.B(n_1412),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1493),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1434),
.A2(n_1465),
.B(n_1478),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1503),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1442),
.B(n_1412),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1497),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1501),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1545),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1412),
.B(n_1543),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1508),
.B(n_1452),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1489),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1543),
.B(n_1518),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1428),
.A2(n_1531),
.B1(n_1539),
.B2(n_1485),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1494),
.A2(n_1495),
.B(n_1511),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1520),
.B(n_1458),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1543),
.B(n_1518),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1507),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1512),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1512),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1519),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1519),
.Y(n_1656)
);

CKINVDCx20_ASAP7_75t_R g1657 ( 
.A(n_1598),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1609),
.B(n_1402),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1645),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1555),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1635),
.B(n_1515),
.Y(n_1661)
);

AND2x2_ASAP7_75t_SL g1662 ( 
.A(n_1645),
.B(n_1539),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1635),
.B(n_1519),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1645),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1580),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1636),
.B(n_1640),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1636),
.B(n_1519),
.Y(n_1667)
);

INVxp67_ASAP7_75t_SL g1668 ( 
.A(n_1632),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1563),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_1610),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1646),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1585),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1613),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1565),
.B(n_1514),
.Y(n_1674)
);

INVxp67_ASAP7_75t_SL g1675 ( 
.A(n_1595),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1578),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1568),
.B(n_1546),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1570),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1568),
.B(n_1546),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1585),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1566),
.B(n_1548),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1572),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1574),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1580),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1634),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1602),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1558),
.B(n_1487),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1646),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1567),
.B(n_1505),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1577),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1567),
.B(n_1505),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1644),
.B(n_1505),
.Y(n_1692)
);

INVx5_ASAP7_75t_L g1693 ( 
.A(n_1583),
.Y(n_1693)
);

NOR2x1_ASAP7_75t_R g1694 ( 
.A(n_1583),
.B(n_1454),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1626),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1608),
.B(n_1487),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1608),
.B(n_1487),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1651),
.B(n_1526),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1584),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1651),
.B(n_1526),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1581),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1601),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1557),
.B(n_1487),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1612),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1566),
.B(n_1506),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_SL g1706 ( 
.A1(n_1594),
.A2(n_1470),
.B1(n_1440),
.B2(n_1474),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1616),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1600),
.Y(n_1708)
);

INVx5_ASAP7_75t_L g1709 ( 
.A(n_1586),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1594),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1557),
.B(n_1513),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1600),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1556),
.B(n_1458),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1597),
.B(n_1547),
.Y(n_1714)
);

INVx5_ASAP7_75t_L g1715 ( 
.A(n_1586),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1607),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1637),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1597),
.B(n_1529),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1604),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1639),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1604),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1592),
.B(n_1463),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1579),
.B(n_1529),
.Y(n_1723)
);

AOI21xp33_ASAP7_75t_L g1724 ( 
.A1(n_1576),
.A2(n_1485),
.B(n_1504),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1593),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1660),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1693),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1666),
.B(n_1655),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1681),
.B(n_1664),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1666),
.B(n_1655),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1708),
.B(n_1641),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1696),
.B(n_1623),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1714),
.B(n_1656),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1670),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1714),
.B(n_1656),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1712),
.B(n_1575),
.Y(n_1736)
);

INVxp67_ASAP7_75t_SL g1737 ( 
.A(n_1676),
.Y(n_1737)
);

NAND2x1_ASAP7_75t_L g1738 ( 
.A(n_1664),
.B(n_1560),
.Y(n_1738)
);

NOR2xp67_ASAP7_75t_L g1739 ( 
.A(n_1693),
.B(n_1614),
.Y(n_1739)
);

OAI21xp33_ASAP7_75t_L g1740 ( 
.A1(n_1711),
.A2(n_1561),
.B(n_1624),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1663),
.B(n_1667),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1685),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1681),
.B(n_1589),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1663),
.B(n_1587),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1667),
.B(n_1588),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1701),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1681),
.B(n_1589),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1672),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1725),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1697),
.B(n_1588),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1685),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1692),
.B(n_1590),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1672),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1692),
.B(n_1689),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1665),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1719),
.B(n_1629),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1721),
.B(n_1630),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1686),
.B(n_1618),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1722),
.A2(n_1615),
.B1(n_1571),
.B2(n_1573),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1689),
.B(n_1589),
.Y(n_1760)
);

INVxp67_ASAP7_75t_SL g1761 ( 
.A(n_1680),
.Y(n_1761)
);

INVx2_ASAP7_75t_SL g1762 ( 
.A(n_1693),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1687),
.A2(n_1713),
.B1(n_1662),
.B2(n_1571),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1691),
.B(n_1562),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1718),
.B(n_1562),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1662),
.A2(n_1638),
.B1(n_1649),
.B2(n_1559),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1677),
.B(n_1648),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1679),
.B(n_1647),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1664),
.B(n_1562),
.Y(n_1769)
);

NOR2x1_ASAP7_75t_SL g1770 ( 
.A(n_1693),
.B(n_1559),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1718),
.B(n_1562),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1706),
.A2(n_1522),
.B(n_1571),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1695),
.Y(n_1773)
);

AND2x2_ASAP7_75t_SL g1774 ( 
.A(n_1659),
.B(n_1522),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1717),
.B(n_1628),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1742),
.Y(n_1776)
);

INVx2_ASAP7_75t_SL g1777 ( 
.A(n_1755),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1734),
.B(n_1668),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1741),
.B(n_1675),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1741),
.B(n_1728),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1742),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1754),
.B(n_1661),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1726),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1755),
.Y(n_1784)
);

INVx3_ASAP7_75t_L g1785 ( 
.A(n_1743),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1754),
.B(n_1661),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1751),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1751),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1727),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1764),
.B(n_1703),
.Y(n_1790)
);

INVx4_ASAP7_75t_L g1791 ( 
.A(n_1727),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1764),
.B(n_1698),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1768),
.B(n_1679),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1768),
.B(n_1658),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1765),
.B(n_1723),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1752),
.B(n_1750),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1765),
.B(n_1700),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1771),
.B(n_1723),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1771),
.B(n_1674),
.Y(n_1799)
);

INVxp67_ASAP7_75t_L g1800 ( 
.A(n_1746),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1728),
.B(n_1702),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1743),
.B(n_1705),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1762),
.B(n_1693),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1737),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1748),
.Y(n_1805)
);

INVx2_ASAP7_75t_SL g1806 ( 
.A(n_1762),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1733),
.B(n_1674),
.Y(n_1807)
);

OAI21xp33_ASAP7_75t_L g1808 ( 
.A1(n_1795),
.A2(n_1740),
.B(n_1766),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1776),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1791),
.A2(n_1763),
.B1(n_1759),
.B2(n_1772),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1782),
.B(n_1760),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1776),
.Y(n_1812)
);

AOI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1800),
.A2(n_1749),
.B1(n_1724),
.B2(n_1673),
.C(n_1758),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1781),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1783),
.Y(n_1815)
);

AOI21xp33_ASAP7_75t_SL g1816 ( 
.A1(n_1789),
.A2(n_1422),
.B(n_1471),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1781),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1782),
.B(n_1786),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1796),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1783),
.Y(n_1820)
);

INVx3_ASAP7_75t_SL g1821 ( 
.A(n_1791),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1807),
.B(n_1732),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1795),
.B(n_1798),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1805),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1786),
.B(n_1760),
.Y(n_1825)
);

OAI221xp5_ASAP7_75t_L g1826 ( 
.A1(n_1804),
.A2(n_1773),
.B1(n_1736),
.B2(n_1688),
.C(n_1622),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1807),
.B(n_1732),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1791),
.A2(n_1774),
.B1(n_1671),
.B2(n_1715),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1783),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1787),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1787),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1788),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1784),
.Y(n_1833)
);

INVxp67_ASAP7_75t_SL g1834 ( 
.A(n_1806),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1788),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1798),
.B(n_1730),
.Y(n_1836)
);

AOI21xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1821),
.A2(n_1789),
.B(n_1777),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1808),
.B(n_1792),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1833),
.Y(n_1839)
);

OAI22xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1821),
.A2(n_1803),
.B1(n_1777),
.B2(n_1806),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1819),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1824),
.Y(n_1842)
);

NAND3xp33_ASAP7_75t_L g1843 ( 
.A(n_1813),
.B(n_1778),
.C(n_1753),
.Y(n_1843)
);

AOI321xp33_ASAP7_75t_L g1844 ( 
.A1(n_1810),
.A2(n_1779),
.A3(n_1801),
.B1(n_1769),
.B2(n_1716),
.C(n_1761),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1809),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1826),
.A2(n_1774),
.B1(n_1769),
.B2(n_1767),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1823),
.B(n_1780),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1822),
.B(n_1799),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1822),
.B(n_1799),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_SL g1850 ( 
.A1(n_1834),
.A2(n_1770),
.B1(n_1785),
.B2(n_1774),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1828),
.A2(n_1790),
.B1(n_1802),
.B2(n_1730),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1815),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1812),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_SL g1854 ( 
.A1(n_1816),
.A2(n_1606),
.B(n_1605),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1812),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1836),
.A2(n_1738),
.B(n_1739),
.Y(n_1856)
);

AOI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1827),
.A2(n_1790),
.B1(n_1802),
.B2(n_1745),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1818),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1814),
.Y(n_1859)
);

OAI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1858),
.A2(n_1785),
.B1(n_1739),
.B2(n_1793),
.Y(n_1860)
);

AOI221xp5_ASAP7_75t_L g1861 ( 
.A1(n_1838),
.A2(n_1825),
.B1(n_1811),
.B2(n_1797),
.C(n_1835),
.Y(n_1861)
);

OAI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1844),
.A2(n_1785),
.B1(n_1793),
.B2(n_1794),
.C(n_1814),
.Y(n_1862)
);

AOI211xp5_ASAP7_75t_L g1863 ( 
.A1(n_1840),
.A2(n_1694),
.B(n_1802),
.C(n_1794),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1847),
.B(n_1415),
.Y(n_1864)
);

AOI222xp33_ASAP7_75t_L g1865 ( 
.A1(n_1843),
.A2(n_1756),
.B1(n_1757),
.B2(n_1619),
.C1(n_1620),
.C2(n_1797),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1848),
.B(n_1815),
.Y(n_1866)
);

AOI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1851),
.A2(n_1802),
.B1(n_1744),
.B2(n_1745),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1842),
.Y(n_1868)
);

XNOR2x1_ASAP7_75t_L g1869 ( 
.A(n_1857),
.B(n_1582),
.Y(n_1869)
);

OAI211xp5_ASAP7_75t_L g1870 ( 
.A1(n_1837),
.A2(n_1454),
.B(n_1657),
.C(n_1479),
.Y(n_1870)
);

A2O1A1Ixp33_ASAP7_75t_L g1871 ( 
.A1(n_1854),
.A2(n_1847),
.B(n_1850),
.C(n_1856),
.Y(n_1871)
);

OAI221xp5_ASAP7_75t_L g1872 ( 
.A1(n_1846),
.A2(n_1835),
.B1(n_1832),
.B2(n_1831),
.C(n_1830),
.Y(n_1872)
);

AOI221xp5_ASAP7_75t_SL g1873 ( 
.A1(n_1846),
.A2(n_1657),
.B1(n_1479),
.B2(n_1775),
.C(n_1731),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1871),
.A2(n_1839),
.B(n_1841),
.Y(n_1874)
);

AOI211xp5_ASAP7_75t_L g1875 ( 
.A1(n_1870),
.A2(n_1510),
.B(n_1849),
.C(n_1767),
.Y(n_1875)
);

AOI221xp5_ASAP7_75t_L g1876 ( 
.A1(n_1872),
.A2(n_1859),
.B1(n_1845),
.B2(n_1853),
.C(n_1855),
.Y(n_1876)
);

NAND3xp33_ASAP7_75t_L g1877 ( 
.A(n_1873),
.B(n_1852),
.C(n_1830),
.Y(n_1877)
);

NAND4xp25_ASAP7_75t_L g1878 ( 
.A(n_1873),
.B(n_1510),
.C(n_1490),
.D(n_1491),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1863),
.A2(n_1852),
.B(n_1715),
.Y(n_1879)
);

AOI322xp5_ASAP7_75t_L g1880 ( 
.A1(n_1861),
.A2(n_1744),
.A3(n_1752),
.B1(n_1735),
.B2(n_1733),
.C1(n_1669),
.C2(n_1707),
.Y(n_1880)
);

OAI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1865),
.A2(n_1720),
.B(n_1715),
.Y(n_1881)
);

AOI221x1_ASAP7_75t_L g1882 ( 
.A1(n_1864),
.A2(n_1642),
.B1(n_1652),
.B2(n_1831),
.C(n_1817),
.Y(n_1882)
);

AOI32xp33_ASAP7_75t_L g1883 ( 
.A1(n_1869),
.A2(n_1684),
.A3(n_1665),
.B1(n_1743),
.B2(n_1747),
.Y(n_1883)
);

AOI221xp5_ASAP7_75t_L g1884 ( 
.A1(n_1862),
.A2(n_1832),
.B1(n_1817),
.B2(n_1683),
.C(n_1690),
.Y(n_1884)
);

AOI211xp5_ASAP7_75t_SL g1885 ( 
.A1(n_1860),
.A2(n_1440),
.B(n_1586),
.C(n_1605),
.Y(n_1885)
);

AOI211xp5_ASAP7_75t_SL g1886 ( 
.A1(n_1868),
.A2(n_1605),
.B(n_1606),
.C(n_1564),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1867),
.A2(n_1747),
.B1(n_1743),
.B2(n_1729),
.Y(n_1887)
);

AOI221xp5_ASAP7_75t_L g1888 ( 
.A1(n_1866),
.A2(n_1682),
.B1(n_1704),
.B2(n_1678),
.C(n_1699),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1871),
.A2(n_1709),
.B(n_1603),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1877),
.Y(n_1890)
);

INVx1_ASAP7_75t_SL g1891 ( 
.A(n_1889),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1882),
.Y(n_1892)
);

NOR4xp25_ASAP7_75t_L g1893 ( 
.A(n_1878),
.B(n_1876),
.C(n_1884),
.D(n_1883),
.Y(n_1893)
);

NAND4xp25_ASAP7_75t_L g1894 ( 
.A(n_1875),
.B(n_1591),
.C(n_1627),
.D(n_1684),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1888),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_SL g1896 ( 
.A(n_1886),
.B(n_1603),
.C(n_1445),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1887),
.B(n_1747),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1880),
.B(n_1820),
.Y(n_1898)
);

NAND3xp33_ASAP7_75t_SL g1899 ( 
.A(n_1874),
.B(n_1885),
.C(n_1881),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1879),
.B(n_1820),
.Y(n_1900)
);

NOR4xp25_ASAP7_75t_L g1901 ( 
.A(n_1890),
.B(n_1631),
.C(n_1643),
.D(n_1633),
.Y(n_1901)
);

AND4x1_ASAP7_75t_L g1902 ( 
.A(n_1893),
.B(n_1654),
.C(n_1653),
.D(n_1509),
.Y(n_1902)
);

NOR2x1_ASAP7_75t_L g1903 ( 
.A(n_1899),
.B(n_1626),
.Y(n_1903)
);

NAND4xp25_ASAP7_75t_L g1904 ( 
.A(n_1894),
.B(n_1627),
.C(n_1650),
.D(n_1621),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1892),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1898),
.B(n_1829),
.Y(n_1906)
);

NOR3xp33_ASAP7_75t_L g1907 ( 
.A(n_1896),
.B(n_1891),
.C(n_1895),
.Y(n_1907)
);

NOR3xp33_ASAP7_75t_L g1908 ( 
.A(n_1900),
.B(n_1643),
.C(n_1631),
.Y(n_1908)
);

NOR2x1_ASAP7_75t_L g1909 ( 
.A(n_1897),
.B(n_1617),
.Y(n_1909)
);

NAND3xp33_ASAP7_75t_L g1910 ( 
.A(n_1902),
.B(n_1897),
.C(n_1599),
.Y(n_1910)
);

NAND3xp33_ASAP7_75t_L g1911 ( 
.A(n_1905),
.B(n_1611),
.C(n_1596),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1906),
.B(n_1829),
.Y(n_1912)
);

NAND4xp75_ASAP7_75t_L g1913 ( 
.A(n_1903),
.B(n_1611),
.C(n_1710),
.D(n_1569),
.Y(n_1913)
);

OR4x2_ASAP7_75t_L g1914 ( 
.A(n_1907),
.B(n_1901),
.C(n_1909),
.D(n_1904),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1908),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1915),
.B(n_1910),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1911),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1914),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1912),
.Y(n_1919)
);

OAI22x1_ASAP7_75t_L g1920 ( 
.A1(n_1918),
.A2(n_1913),
.B1(n_1625),
.B2(n_1538),
.Y(n_1920)
);

XNOR2x1_ASAP7_75t_L g1921 ( 
.A(n_1916),
.B(n_1466),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1919),
.Y(n_1922)
);

BUFx2_ASAP7_75t_L g1923 ( 
.A(n_1917),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1923),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1922),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1921),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1924),
.Y(n_1927)
);

XNOR2xp5_ASAP7_75t_L g1928 ( 
.A(n_1927),
.B(n_1924),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1928),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1929),
.A2(n_1926),
.B1(n_1925),
.B2(n_1920),
.Y(n_1930)
);


endmodule