module fake_jpeg_15925_n_359 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_359);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_20),
.B(n_10),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_19),
.B(n_0),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_45),
.B(n_39),
.Y(n_61)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx2_ASAP7_75t_SL g105 ( 
.A(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_61),
.B(n_71),
.Y(n_104)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_37),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_75),
.Y(n_103)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_38),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_76),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_34),
.B1(n_26),
.B2(n_19),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_48),
.B1(n_51),
.B2(n_34),
.Y(n_91)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_97),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_53),
.B1(n_56),
.B2(n_51),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_92),
.B1(n_93),
.B2(n_101),
.Y(n_119)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_91),
.B1(n_108),
.B2(n_32),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_34),
.B1(n_44),
.B2(n_49),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_55),
.B1(n_52),
.B2(n_49),
.Y(n_93)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_55),
.B1(n_52),
.B2(n_46),
.Y(n_101)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_58),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_57),
.A2(n_30),
.B1(n_22),
.B2(n_32),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_74),
.B(n_50),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_30),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_113),
.Y(n_120)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_59),
.B1(n_57),
.B2(n_80),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_131),
.B1(n_102),
.B2(n_114),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_70),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_127),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_27),
.B(n_76),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_124),
.Y(n_151)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_129),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_59),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_35),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_125),
.B(n_126),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_35),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_78),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_142),
.B1(n_143),
.B2(n_96),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_79),
.B1(n_78),
.B2(n_66),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_132),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_89),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_138),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_38),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_36),
.B(n_37),
.C(n_23),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_100),
.B(n_22),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_99),
.Y(n_140)
);

INVxp33_ASAP7_75t_SL g149 ( 
.A(n_140),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_141),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_101),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_88),
.A2(n_79),
.B1(n_21),
.B2(n_62),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_90),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_154),
.B1(n_166),
.B2(n_134),
.Y(n_175)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_96),
.B1(n_94),
.B2(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_28),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_159),
.C(n_116),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_28),
.C(n_29),
.Y(n_159)
);

OAI22x1_ASAP7_75t_SL g160 ( 
.A1(n_117),
.A2(n_25),
.B1(n_33),
.B2(n_28),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_166),
.B1(n_124),
.B2(n_115),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_138),
.B(n_126),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_162),
.A2(n_135),
.B1(n_116),
.B2(n_123),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_164),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_128),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_120),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

AO22x2_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_94),
.B1(n_25),
.B2(n_29),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_180),
.B1(n_181),
.B2(n_191),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_166),
.B1(n_153),
.B2(n_146),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_124),
.B(n_135),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_188),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_119),
.B1(n_131),
.B2(n_140),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_192),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_155),
.A2(n_119),
.B1(n_141),
.B2(n_122),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_185),
.A2(n_166),
.B1(n_147),
.B2(n_168),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_129),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_179),
.C(n_174),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_190),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_151),
.A2(n_132),
.B(n_137),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_167),
.B(n_33),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_123),
.B(n_122),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_133),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_152),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_195),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_13),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_215),
.C(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_157),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_191),
.B1(n_182),
.B2(n_161),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_194),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_207),
.B(n_213),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_128),
.B1(n_145),
.B2(n_136),
.Y(n_240)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_159),
.C(n_154),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_150),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_220),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_218),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_184),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_0),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_169),
.C(n_149),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_175),
.B1(n_181),
.B2(n_195),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_224),
.A2(n_234),
.B1(n_240),
.B2(n_218),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_188),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_232),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_227),
.B(n_237),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_222),
.A2(n_180),
.B1(n_160),
.B2(n_190),
.Y(n_231)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_176),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_184),
.B1(n_173),
.B2(n_196),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_238),
.Y(n_257)
);

AO21x2_ASAP7_75t_SL g236 ( 
.A1(n_222),
.A2(n_163),
.B(n_161),
.Y(n_236)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_223),
.B(n_156),
.Y(n_237)
);

NAND2x1_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_128),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_145),
.C(n_136),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_244),
.C(n_205),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_171),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_210),
.A2(n_145),
.B1(n_33),
.B2(n_2),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_246),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

BUFx12_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_202),
.Y(n_252)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_198),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_219),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_254),
.B(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_198),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_243),
.C(n_233),
.Y(n_280)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_261),
.B1(n_272),
.B2(n_247),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_206),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_263),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_197),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_200),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_267),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_226),
.B(n_209),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_208),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_271),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_215),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_244),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_212),
.Y(n_271)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_247),
.B1(n_260),
.B2(n_269),
.Y(n_275)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_251),
.B(n_232),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_276),
.B(n_252),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_281),
.C(n_285),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_225),
.C(n_245),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_224),
.C(n_235),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_230),
.C(n_218),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_287),
.C(n_288),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_230),
.C(n_214),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_236),
.B(n_249),
.Y(n_289)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_260),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_290)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_264),
.A2(n_258),
.B1(n_266),
.B2(n_262),
.Y(n_291)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_29),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_257),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_299),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_255),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_302),
.C(n_281),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_283),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_307),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_271),
.C(n_266),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_282),
.B(n_261),
.Y(n_303)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_276),
.B(n_250),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_1),
.Y(n_317)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_284),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_3),
.C(n_5),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_277),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_312),
.C(n_314),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_294),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_7),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_285),
.B1(n_287),
.B2(n_278),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_288),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_318),
.C(n_7),
.Y(n_333)
);

OAI321xp33_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_292),
.A3(n_250),
.B1(n_12),
.B2(n_4),
.C(n_5),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_316),
.A2(n_14),
.B(n_5),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_321),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_11),
.Y(n_318)
);

FAx1_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_2),
.CI(n_3),
.CON(n_319),
.SN(n_319)
);

OA21x2_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_3),
.B(n_4),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_293),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_324),
.Y(n_340)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_302),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_325),
.B(n_329),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_10),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_306),
.B1(n_296),
.B2(n_297),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_331),
.C(n_333),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_310),
.A2(n_7),
.B(n_8),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_332),
.B(n_9),
.Y(n_339)
);

FAx1_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_8),
.CI(n_9),
.CON(n_334),
.SN(n_334)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_13),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_310),
.B(n_321),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_335),
.A2(n_326),
.B(n_334),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_330),
.A2(n_317),
.B1(n_10),
.B2(n_12),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_343),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_342),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_23),
.C(n_13),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_14),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_347),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_334),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_348),
.A2(n_341),
.B(n_16),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_337),
.B(n_323),
.Y(n_349)
);

O2A1O1Ixp33_ASAP7_75t_SL g351 ( 
.A1(n_349),
.A2(n_336),
.B(n_343),
.C(n_323),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_351),
.B(n_352),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_353),
.A2(n_350),
.B(n_344),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_346),
.B(n_17),
.C(n_18),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_15),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_SL g357 ( 
.A(n_356),
.B(n_17),
.C(n_23),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_17),
.Y(n_358)
);

FAx1_ASAP7_75t_SL g359 ( 
.A(n_358),
.B(n_23),
.CI(n_356),
.CON(n_359),
.SN(n_359)
);


endmodule