module fake_jpeg_22127_n_45 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_45);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_2),
.A2(n_9),
.B1(n_6),
.B2(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_14),
.B1(n_20),
.B2(n_19),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_24),
.B(n_21),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_35),
.B(n_31),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_25),
.B1(n_16),
.B2(n_7),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_33),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_39),
.B(n_33),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_45)
);


endmodule