module fake_jpeg_32181_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_28),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx11_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

INVx11_ASAP7_75t_SL g71 ( 
.A(n_30),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_20),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_0),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_66),
.Y(n_81)
);

CKINVDCx6p67_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_79),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_78),
.Y(n_90)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_65),
.Y(n_97)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_89),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_63),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_71),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_103),
.Y(n_125)
);

BUFx16f_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_67),
.B1(n_63),
.B2(n_57),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_88),
.B1(n_67),
.B2(n_59),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_104),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_68),
.B1(n_65),
.B2(n_54),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_76),
.B(n_64),
.C(n_73),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_57),
.C(n_53),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_60),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_77),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_74),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_115),
.B1(n_50),
.B2(n_15),
.Y(n_133)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_120),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_116),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_128),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_114),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_83),
.B1(n_85),
.B2(n_72),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_55),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_122),
.Y(n_130)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_121),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_56),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_0),
.C(n_1),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_76),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_19),
.A3(n_49),
.B1(n_45),
.B2(n_43),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_29),
.B(n_31),
.C(n_32),
.D(n_34),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_137),
.B1(n_142),
.B2(n_150),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_3),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_139),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_17),
.B1(n_39),
.B2(n_36),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_5),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_6),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_147),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_41),
.B1(n_14),
.B2(n_24),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_13),
.C(n_33),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_133),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_8),
.Y(n_156)
);

NAND2x1_ASAP7_75t_SL g145 ( 
.A(n_112),
.B(n_6),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_7),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_7),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_137),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_150)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_12),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_163),
.B1(n_160),
.B2(n_161),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_136),
.B(n_134),
.C(n_145),
.D(n_146),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_143),
.C(n_131),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_142),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_169),
.B(n_172),
.CI(n_171),
.CON(n_177),
.SN(n_177)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_159),
.B1(n_165),
.B2(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_176),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_177),
.B(n_166),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_174),
.B(n_175),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_177),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_179),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_176),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_181),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_179),
.Y(n_188)
);


endmodule