module fake_jpeg_17492_n_324 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_2),
.B(n_6),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_40),
.B(n_45),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_42),
.B(n_49),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_54),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_SL g49 ( 
.A(n_28),
.B(n_7),
.C(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx2_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_25),
.B(n_8),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_63),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_60),
.Y(n_93)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_0),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_69),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_25),
.B(n_8),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_9),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_73),
.B(n_83),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_20),
.B1(n_34),
.B2(n_23),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_76),
.A2(n_96),
.B1(n_101),
.B2(n_116),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_84),
.Y(n_121)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_1),
.Y(n_83)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_39),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_85),
.B(n_91),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_89),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_37),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_90),
.B(n_95),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_37),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_32),
.B1(n_33),
.B2(n_19),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_58),
.B(n_33),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_98),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_48),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_16),
.B1(n_34),
.B2(n_20),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_114),
.B1(n_118),
.B2(n_87),
.Y(n_135)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_41),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_107),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_43),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_17),
.B1(n_23),
.B2(n_14),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_42),
.B(n_29),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_55),
.A2(n_17),
.B1(n_14),
.B2(n_29),
.Y(n_116)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_64),
.B(n_27),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_27),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_46),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_27),
.B1(n_101),
.B2(n_83),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_83),
.A2(n_56),
.B1(n_3),
.B2(n_12),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_123),
.A2(n_152),
.B1(n_82),
.B2(n_79),
.Y(n_178)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_132),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_72),
.B(n_12),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_131),
.B(n_133),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_3),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_47),
.B(n_14),
.C(n_29),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_136),
.B(n_153),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_135),
.A2(n_149),
.B1(n_132),
.B2(n_150),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_83),
.A2(n_27),
.B(n_29),
.C(n_64),
.Y(n_136)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_141),
.A2(n_145),
.B1(n_129),
.B2(n_166),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_142),
.B(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_147),
.Y(n_176)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_86),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_157),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_88),
.A2(n_120),
.B1(n_110),
.B2(n_94),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_77),
.A2(n_94),
.B1(n_105),
.B2(n_79),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_74),
.B(n_76),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_154),
.B(n_89),
.Y(n_179)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_159),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_116),
.B(n_93),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_163),
.C(n_130),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_93),
.B(n_78),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_162),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_177),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_173),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_175),
.B(n_178),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_162),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_190),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_142),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_122),
.B(n_71),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_190),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_135),
.A2(n_80),
.B1(n_71),
.B2(n_89),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_193),
.B1(n_196),
.B2(n_199),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g188 ( 
.A(n_155),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_155),
.B(n_109),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_189),
.B(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_125),
.B(n_124),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_134),
.B1(n_137),
.B2(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_136),
.B(n_163),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_198),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_127),
.B1(n_158),
.B2(n_149),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_167),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_192),
.B(n_195),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_128),
.B(n_161),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_145),
.A2(n_163),
.B1(n_140),
.B2(n_148),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_129),
.A2(n_146),
.B1(n_141),
.B2(n_151),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_175),
.B(n_168),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_224),
.B(n_229),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_211),
.C(n_220),
.Y(n_246)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_193),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_209),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_210),
.B(n_233),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_194),
.C(n_203),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_215),
.A2(n_219),
.B1(n_212),
.B2(n_213),
.Y(n_249)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_176),
.A2(n_178),
.B(n_168),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_205),
.B(n_213),
.C(n_220),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_221),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_186),
.B1(n_181),
.B2(n_204),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_185),
.C(n_201),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_191),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_184),
.C(n_169),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_232),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_171),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_230),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_183),
.B(n_172),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_214),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_230),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_174),
.B(n_187),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_195),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_234),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_180),
.B(n_197),
.C(n_177),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_211),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_214),
.A2(n_180),
.B1(n_209),
.B2(n_225),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_237),
.A2(n_242),
.B1(n_249),
.B2(n_256),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_241),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_247),
.C(n_252),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_218),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_234),
.B1(n_212),
.B2(n_219),
.Y(n_242)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_233),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_250),
.A2(n_258),
.B(n_236),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_232),
.B(n_222),
.Y(n_252)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_208),
.C(n_227),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_257),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_216),
.A2(n_235),
.B1(n_228),
.B2(n_207),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_263),
.A2(n_273),
.B(n_277),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_240),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_265),
.C(n_278),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_256),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_272),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_258),
.B(n_255),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_255),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_274),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_276),
.B(n_238),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_258),
.A2(n_236),
.B(n_239),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_247),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_245),
.C(n_241),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_291),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_277),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_242),
.C(n_248),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_294),
.C(n_281),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_262),
.A2(n_238),
.B(n_260),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_276),
.B1(n_270),
.B2(n_269),
.Y(n_306)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_293),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_260),
.C(n_243),
.Y(n_294)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_271),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_295),
.A2(n_243),
.B1(n_272),
.B2(n_266),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_295),
.B1(n_293),
.B2(n_285),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_300),
.C(n_302),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_265),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_263),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_305),
.C(n_289),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_273),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_299),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_275),
.C(n_269),
.Y(n_305)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_306),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_298),
.A2(n_283),
.B(n_290),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_307),
.B(n_309),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_310),
.C(n_312),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_284),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g314 ( 
.A1(n_301),
.A2(n_292),
.B(n_295),
.C(n_283),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_302),
.C(n_305),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_316),
.A2(n_309),
.B(n_313),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g318 ( 
.A(n_317),
.B(n_300),
.CI(n_308),
.CON(n_318),
.SN(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);

NAND5xp2_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_317),
.C(n_315),
.D(n_288),
.E(n_314),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_318),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_320),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_288),
.Y(n_324)
);


endmodule