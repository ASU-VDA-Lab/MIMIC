module real_jpeg_13580_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_289, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_289;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_243;
wire n_105;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_267;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_283;
wire n_181;
wire n_85;
wire n_81;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_0),
.A2(n_37),
.B1(n_46),
.B2(n_47),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_0),
.A2(n_10),
.B(n_33),
.C(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_0),
.A2(n_37),
.B1(n_57),
.B2(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_0),
.B(n_38),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_0),
.B(n_55),
.C(n_58),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_0),
.B(n_45),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_0),
.B(n_30),
.C(n_34),
.Y(n_166)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_3),
.Y(n_99)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_41),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_6),
.A2(n_41),
.B1(n_57),
.B2(n_58),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_6),
.A2(n_41),
.B1(n_46),
.B2(n_47),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_49),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_8),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_201)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_9),
.Y(n_286)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

AO22x1_ASAP7_75t_L g45 ( 
.A1(n_10),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_15),
.B(n_285),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_12),
.B(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_27),
.B1(n_46),
.B2(n_47),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_13),
.A2(n_27),
.B1(n_57),
.B2(n_58),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_281),
.B(n_283),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_73),
.B(n_280),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_70),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_18),
.B(n_70),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_63),
.C(n_67),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_19),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.C(n_50),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_20),
.A2(n_106),
.B1(n_116),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_20),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_20),
.B(n_116),
.C(n_179),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_20),
.A2(n_82),
.B1(n_83),
.B2(n_181),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_20),
.A2(n_181),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_28),
.B1(n_36),
.B2(n_38),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_22),
.A2(n_32),
.B(n_69),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_24),
.B(n_166),
.Y(n_165)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_28),
.B(n_36),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_28),
.B(n_38),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_32),
.A2(n_68),
.B(n_69),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_32),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_43),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp33_ASAP7_75t_L g237 ( 
.A(n_36),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_SL g95 ( 
.A1(n_37),
.A2(n_43),
.B(n_46),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_37),
.B(n_102),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_37),
.B(n_61),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_39),
.A2(n_50),
.B1(n_255),
.B2(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_39),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_39)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_40),
.Y(n_257)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_47),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_50),
.A2(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_50),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_50),
.B(n_169),
.C(n_256),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_61),
.B(n_62),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_51),
.A2(n_61),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_91),
.Y(n_90)
);

AO22x1_ASAP7_75t_SL g121 ( 
.A1(n_52),
.A2(n_56),
.B1(n_89),
.B2(n_91),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_52),
.A2(n_56),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

AO22x1_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_57),
.B(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_88),
.B(n_90),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_61),
.A2(n_90),
.B(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_62),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_63),
.B(n_67),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_66),
.B1(n_84),
.B2(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_65),
.A2(n_66),
.B(n_107),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_66),
.A2(n_85),
.B(n_257),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_70),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_70),
.B(n_282),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_72),
.B(n_238),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_275),
.B(n_279),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_247),
.B(n_272),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_225),
.B(n_246),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_208),
.B(n_224),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_176),
.A3(n_203),
.B1(n_206),
.B2(n_207),
.C(n_289),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_158),
.B(n_175),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_124),
.B(n_157),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_103),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_81),
.B(n_103),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_87),
.C(n_92),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_141),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_82),
.A2(n_83),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_83),
.B(n_168),
.C(n_173),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_83),
.B(n_181),
.C(n_213),
.Y(n_245)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_87),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_87),
.A2(n_128),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_87),
.A2(n_141),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_92),
.A2(n_93),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_98),
.B(n_201),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_101),
.A2(n_102),
.B1(n_184),
.B2(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_102),
.A2(n_114),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_118),
.B2(n_119),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_104),
.B(n_121),
.C(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B1(n_116),
.B2(n_117),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_109),
.C(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_111),
.B(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_112),
.B(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_116),
.A2(n_241),
.B(n_244),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_116),
.B(n_241),
.Y(n_244)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_123),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_133),
.C(n_135),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_121),
.A2(n_123),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_121),
.B(n_200),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_151),
.B(n_156),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_137),
.B(n_150),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_132),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_135),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_135),
.B(n_147),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_164),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_142),
.B(n_149),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_183),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.B(n_148),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_160),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_163),
.C(n_167),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_169),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_191),
.C(n_196),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_168),
.A2(n_169),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_168),
.A2(n_169),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_169),
.B(n_266),
.C(n_270),
.Y(n_278)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_187),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_187),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.C(n_186),
.Y(n_177)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_178),
.B(n_182),
.CI(n_186),
.CON(n_205),
.SN(n_205)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_202),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_197),
.B2(n_198),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_198),
.C(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_205),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_223),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_223),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_212),
.C(n_217),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_218),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_220),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_222),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_222),
.A2(n_231),
.B(n_236),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_227),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_245),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_239),
.B2(n_240),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_239),
.C(n_245),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_244),
.A2(n_251),
.B1(n_252),
.B2(n_259),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_244),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_262),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_261),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_261),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_260),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_259),
.C(n_260),
.Y(n_271)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_256),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_271),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_271),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_270),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_278),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);


endmodule