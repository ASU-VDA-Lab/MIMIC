module fake_jpeg_22839_n_219 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_37),
.Y(n_59)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_21),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

CKINVDCx9p33_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

NAND4xp25_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_28),
.C(n_18),
.D(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_19),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_31),
.B(n_30),
.C(n_29),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_25),
.B1(n_19),
.B2(n_23),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_64),
.B1(n_16),
.B2(n_17),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_55),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_60),
.B(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_62),
.B(n_21),
.Y(n_101)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_67),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_24),
.B1(n_27),
.B2(n_26),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_50),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_20),
.B1(n_16),
.B2(n_17),
.Y(n_91)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_79),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_77),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_1),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_27),
.C(n_26),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_66),
.Y(n_104)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_85),
.Y(n_107)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NAND2x1_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_21),
.Y(n_111)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_96),
.Y(n_124)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_24),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_46),
.A2(n_30),
.B1(n_29),
.B2(n_31),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_99),
.B1(n_63),
.B2(n_58),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_47),
.A2(n_20),
.B1(n_30),
.B2(n_31),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_103),
.B(n_104),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_118),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_66),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_75),
.B(n_78),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_128),
.B1(n_86),
.B2(n_74),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_72),
.A3(n_73),
.B1(n_51),
.B2(n_56),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_70),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_79),
.Y(n_137)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_122),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_83),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_127),
.Y(n_146)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_73),
.B1(n_72),
.B2(n_55),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_121),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_133),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_55),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_140),
.C(n_141),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_119),
.B1(n_115),
.B2(n_108),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_139),
.B1(n_128),
.B2(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_148),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_95),
.B1(n_86),
.B2(n_49),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_97),
.C(n_102),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_55),
.C(n_81),
.Y(n_141)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_147),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_106),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_94),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_150),
.B(n_3),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_115),
.B1(n_107),
.B2(n_113),
.Y(n_154)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_2),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_3),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_74),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_15),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_156),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_158),
.B1(n_160),
.B2(n_164),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_155),
.B(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_136),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_126),
.B1(n_117),
.B2(n_109),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_124),
.B1(n_127),
.B2(n_112),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_162),
.B(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_14),
.B1(n_11),
.B2(n_8),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_140),
.C(n_135),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_169),
.C(n_171),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_130),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_178),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_132),
.C(n_141),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_166),
.A2(n_133),
.B1(n_148),
.B2(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_153),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_175),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_156),
.B(n_142),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_144),
.B1(n_129),
.B2(n_8),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

BUFx4f_ASAP7_75t_SL g183 ( 
.A(n_181),
.Y(n_183)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_177),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_162),
.C(n_161),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_168),
.C(n_176),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_167),
.B(n_165),
.C(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_191),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_152),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_192),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_194),
.A2(n_201),
.B(n_189),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_183),
.B(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_196),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_177),
.C(n_15),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_191),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_199),
.A2(n_184),
.B1(n_188),
.B2(n_187),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_197),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_188),
.B(n_187),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_201),
.B(n_196),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_210),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

AOI31xp67_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_197),
.A3(n_14),
.B(n_5),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_204),
.B(n_203),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_213),
.B(n_205),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_207),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_216),
.C(n_3),
.Y(n_217)
);

AOI321xp33_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_124),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_218),
.A2(n_4),
.B(n_6),
.Y(n_219)
);


endmodule