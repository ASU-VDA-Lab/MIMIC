module fake_jpeg_18785_n_233 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_14),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_33),
.B1(n_19),
.B2(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_30),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_33),
.B1(n_19),
.B2(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_59),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_26),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_32),
.B1(n_29),
.B2(n_20),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_57),
.A2(n_60),
.B1(n_0),
.B2(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_32),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_29),
.B1(n_17),
.B2(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_26),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_67),
.B(n_74),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_70),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_24),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_91),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_27),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_27),
.B(n_22),
.C(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_79),
.Y(n_115)
);

INVx2_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_21),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_45),
.B(n_13),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_13),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_84),
.Y(n_123)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_28),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_51),
.B(n_41),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_99),
.B(n_10),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_28),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_98),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_66),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_114),
.B1(n_118),
.B2(n_124),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_66),
.A2(n_3),
.B(n_4),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_126),
.B(n_12),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_64),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_76),
.B1(n_88),
.B2(n_83),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_64),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_73),
.A2(n_10),
.B(n_11),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_69),
.B(n_70),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_142),
.B(n_143),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_68),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_128),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_74),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_131),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_67),
.B1(n_65),
.B2(n_99),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_69),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_119),
.C(n_116),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_136),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_135),
.B(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_89),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_71),
.B1(n_84),
.B2(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_82),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_114),
.B1(n_102),
.B2(n_124),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_72),
.Y(n_142)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_104),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_93),
.Y(n_146)
);

OAI22x1_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_98),
.B1(n_92),
.B2(n_85),
.Y(n_147)
);

OAI321xp33_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_113),
.A3(n_109),
.B1(n_121),
.B2(n_123),
.C(n_122),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_87),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_87),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_118),
.Y(n_156)
);

OAI21x1_ASAP7_75t_SL g184 ( 
.A1(n_154),
.A2(n_106),
.B(n_110),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_142),
.B(n_149),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_139),
.C(n_140),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_120),
.B(n_116),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_146),
.B(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_164),
.B(n_151),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_133),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_145),
.Y(n_174)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_131),
.B1(n_137),
.B2(n_141),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_177),
.B1(n_184),
.B2(n_160),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_139),
.B1(n_140),
.B2(n_129),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_143),
.B(n_127),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_152),
.B(n_163),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_162),
.C(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_166),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_185),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_106),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_188),
.C(n_194),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_198),
.B(n_176),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_158),
.C(n_151),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_189),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_150),
.B1(n_165),
.B2(n_161),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_168),
.B1(n_172),
.B2(n_159),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_160),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_152),
.B(n_150),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_202),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_184),
.B1(n_175),
.B2(n_173),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_179),
.C(n_177),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_205),
.C(n_187),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_196),
.A2(n_178),
.B1(n_182),
.B2(n_173),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_204),
.A2(n_207),
.B1(n_208),
.B2(n_197),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_178),
.C(n_180),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_193),
.A2(n_176),
.B1(n_185),
.B2(n_121),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_213),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_200),
.B(n_110),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_209),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_192),
.B(n_191),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_217),
.C(n_108),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_205),
.C(n_202),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_219),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_201),
.B1(n_206),
.B2(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_212),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_221),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_217),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_227),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_223),
.A2(n_211),
.B(n_108),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_107),
.B(n_105),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_228),
.B(n_107),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_230),
.Y(n_233)
);


endmodule