module fake_jpeg_2932_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx2_ASAP7_75t_SL g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_9),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_29),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_11),
.A2(n_20),
.B1(n_16),
.B2(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_11),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_4),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_10),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_12),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_27),
.Y(n_46)
);

OAI32xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_32),
.A3(n_31),
.B1(n_24),
.B2(n_29),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_49),
.C(n_33),
.Y(n_52)
);

AND2x6_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_8),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_28),
.B1(n_21),
.B2(n_15),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_50),
.A2(n_51),
.B1(n_35),
.B2(n_36),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_19),
.B1(n_8),
.B2(n_9),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_37),
.C(n_42),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_37),
.C(n_42),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_48),
.B1(n_47),
.B2(n_50),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_54),
.B1(n_44),
.B2(n_49),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_63),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_60),
.C(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_58),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_61),
.B(n_62),
.Y(n_66)
);

AOI21x1_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_67),
.B(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_44),
.B(n_42),
.Y(n_70)
);

BUFx24_ASAP7_75t_SL g71 ( 
.A(n_70),
.Y(n_71)
);


endmodule