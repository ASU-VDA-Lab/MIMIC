module real_aes_689_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_297;
wire n_383;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_0), .A2(n_53), .B1(n_122), .B2(n_124), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_1), .B(n_211), .Y(n_294) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_2), .A2(n_52), .B1(n_89), .B2(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g176 ( .A(n_3), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_4), .B(n_196), .Y(n_195) );
NAND2xp33_ASAP7_75t_SL g279 ( .A(n_5), .B(n_202), .Y(n_279) );
INVx1_ASAP7_75t_L g270 ( .A(n_6), .Y(n_270) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_7), .A2(n_16), .B1(n_89), .B2(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g190 ( .A(n_8), .B(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g192 ( .A(n_9), .Y(n_192) );
AOI221x1_ASAP7_75t_L g273 ( .A1(n_10), .A2(n_204), .B1(n_274), .B2(n_276), .C(n_278), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g84 ( .A1(n_11), .A2(n_40), .B1(n_85), .B2(n_102), .Y(n_84) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_12), .B(n_196), .Y(n_260) );
OAI22xp5_ASAP7_75t_SL g158 ( .A1(n_13), .A2(n_159), .B1(n_160), .B2(n_163), .Y(n_158) );
INVx1_ASAP7_75t_L g163 ( .A(n_13), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_13), .A2(n_204), .B(n_209), .Y(n_203) );
AOI221xp5_ASAP7_75t_SL g284 ( .A1(n_14), .A2(n_27), .B1(n_196), .B2(n_204), .C(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_15), .B(n_211), .Y(n_210) );
OAI221xp5_ASAP7_75t_L g168 ( .A1(n_16), .A2(n_52), .B1(n_56), .B2(n_169), .C(n_171), .Y(n_168) );
OR2x2_ASAP7_75t_L g193 ( .A(n_17), .B(n_69), .Y(n_193) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_17), .A2(n_69), .B(n_192), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_18), .B(n_213), .Y(n_264) );
INVxp67_ASAP7_75t_L g272 ( .A(n_19), .Y(n_272) );
AND2x2_ASAP7_75t_L g235 ( .A(n_20), .B(n_225), .Y(n_235) );
INVx3_ASAP7_75t_L g89 ( .A(n_21), .Y(n_89) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_22), .A2(n_204), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_23), .B(n_213), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g160 ( .A1(n_24), .A2(n_42), .B1(n_161), .B2(n_162), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_24), .Y(n_161) );
INVx1_ASAP7_75t_SL g90 ( .A(n_25), .Y(n_90) );
INVx1_ASAP7_75t_L g178 ( .A(n_26), .Y(n_178) );
AND2x2_ASAP7_75t_L g202 ( .A(n_26), .B(n_176), .Y(n_202) );
AND2x2_ASAP7_75t_L g205 ( .A(n_26), .B(n_206), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_28), .A2(n_80), .B1(n_81), .B2(n_154), .Y(n_79) );
INVx1_ASAP7_75t_L g154 ( .A(n_28), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_29), .A2(n_61), .B1(n_204), .B2(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_30), .B(n_211), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_31), .A2(n_57), .B1(n_134), .B2(n_138), .Y(n_133) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_32), .A2(n_56), .B1(n_89), .B2(n_94), .Y(n_93) );
AND2x2_ASAP7_75t_L g297 ( .A(n_33), .B(n_225), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_34), .B(n_225), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g106 ( .A1(n_35), .A2(n_55), .B1(n_107), .B2(n_111), .Y(n_106) );
INVx1_ASAP7_75t_L g199 ( .A(n_36), .Y(n_199) );
INVx1_ASAP7_75t_L g208 ( .A(n_36), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_37), .A2(n_70), .B1(n_148), .B2(n_151), .Y(n_147) );
INVx1_ASAP7_75t_L g91 ( .A(n_38), .Y(n_91) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_39), .B(n_196), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g114 ( .A1(n_41), .A2(n_66), .B1(n_115), .B2(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g162 ( .A(n_42), .Y(n_162) );
AND2x2_ASAP7_75t_L g226 ( .A(n_43), .B(n_225), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_44), .B(n_213), .Y(n_295) );
XOR2x2_ASAP7_75t_L g502 ( .A(n_45), .B(n_81), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_46), .B(n_211), .Y(n_222) );
AND2x2_ASAP7_75t_SL g265 ( .A(n_47), .B(n_191), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_48), .A2(n_204), .B(n_231), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_48), .A2(n_80), .B1(n_81), .B2(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_48), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_49), .B(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_SL g255 ( .A(n_50), .B(n_242), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_51), .A2(n_63), .B1(n_141), .B2(n_145), .Y(n_140) );
INVxp33_ASAP7_75t_L g173 ( .A(n_52), .Y(n_173) );
INVx1_ASAP7_75t_L g201 ( .A(n_54), .Y(n_201) );
INVx1_ASAP7_75t_L g206 ( .A(n_54), .Y(n_206) );
INVxp67_ASAP7_75t_L g172 ( .A(n_56), .Y(n_172) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_58), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_59), .B(n_196), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_60), .A2(n_62), .B1(n_196), .B2(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_64), .B(n_211), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_65), .B(n_211), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_67), .A2(n_204), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_68), .B(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_71), .B(n_213), .Y(n_221) );
INVxp67_ASAP7_75t_L g275 ( .A(n_72), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_73), .B(n_196), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_74), .B(n_213), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_75), .A2(n_204), .B(n_262), .Y(n_261) );
BUFx2_ASAP7_75t_SL g170 ( .A(n_76), .Y(n_170) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_165), .B1(n_179), .B2(n_491), .C(n_492), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_155), .Y(n_78) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVxp33_ASAP7_75t_SL g81 ( .A(n_82), .Y(n_81) );
NOR2x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_127), .Y(n_82) );
NAND4xp25_ASAP7_75t_L g83 ( .A(n_84), .B(n_106), .C(n_114), .D(n_121), .Y(n_83) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_95), .Y(n_85) );
AND2x2_ASAP7_75t_L g139 ( .A(n_86), .B(n_112), .Y(n_139) );
AND2x2_ASAP7_75t_L g150 ( .A(n_86), .B(n_120), .Y(n_150) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
INVx2_ASAP7_75t_L g104 ( .A(n_87), .Y(n_104) );
AND2x2_ASAP7_75t_L g132 ( .A(n_87), .B(n_93), .Y(n_132) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_87), .Y(n_153) );
OAI22x1_ASAP7_75t_L g87 ( .A1(n_88), .A2(n_89), .B1(n_90), .B2(n_91), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g94 ( .A(n_89), .Y(n_94) );
INVx2_ASAP7_75t_L g98 ( .A(n_89), .Y(n_98) );
INVx1_ASAP7_75t_L g101 ( .A(n_89), .Y(n_101) );
AND2x4_ASAP7_75t_L g103 ( .A(n_92), .B(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
AND2x2_ASAP7_75t_L g110 ( .A(n_93), .B(n_104), .Y(n_110) );
BUFx2_ASAP7_75t_L g126 ( .A(n_93), .Y(n_126) );
AND2x6_ASAP7_75t_L g109 ( .A(n_95), .B(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_L g117 ( .A(n_95), .B(n_103), .Y(n_117) );
AND2x2_ASAP7_75t_L g131 ( .A(n_95), .B(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g95 ( .A(n_96), .B(n_99), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g105 ( .A(n_97), .B(n_100), .Y(n_105) );
INVx1_ASAP7_75t_L g113 ( .A(n_97), .Y(n_113) );
AND2x4_ASAP7_75t_L g120 ( .A(n_97), .B(n_99), .Y(n_120) );
INVxp67_ASAP7_75t_L g144 ( .A(n_99), .Y(n_144) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g112 ( .A(n_100), .B(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g102 ( .A(n_103), .B(n_105), .Y(n_102) );
AND2x6_ASAP7_75t_L g111 ( .A(n_103), .B(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g119 ( .A(n_103), .B(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g125 ( .A(n_105), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g152 ( .A(n_105), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g123 ( .A(n_110), .B(n_112), .Y(n_123) );
AND2x4_ASAP7_75t_L g146 ( .A(n_110), .B(n_120), .Y(n_146) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_113), .Y(n_137) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx8_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND4xp25_ASAP7_75t_SL g127 ( .A(n_128), .B(n_133), .C(n_140), .D(n_147), .Y(n_127) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx6_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g135 ( .A(n_132), .B(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g143 ( .A(n_132), .B(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx6_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx12f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B1(n_158), .B2(n_164), .Y(n_155) );
INVx1_ASAP7_75t_L g164 ( .A(n_156), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_158), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_167), .Y(n_166) );
AND3x1_ASAP7_75t_SL g167 ( .A(n_168), .B(n_174), .C(n_177), .Y(n_167) );
INVxp67_ASAP7_75t_L g500 ( .A(n_168), .Y(n_500) );
CKINVDCx8_ASAP7_75t_R g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_174), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_174), .A2(n_508), .B(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g247 ( .A(n_175), .B(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_SL g505 ( .A(n_175), .B(n_177), .Y(n_505) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g207 ( .A(n_176), .B(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_177), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2x1p5_ASAP7_75t_L g252 ( .A(n_178), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_413), .Y(n_182) );
NOR3xp33_ASAP7_75t_SL g183 ( .A(n_184), .B(n_337), .C(n_387), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_185), .B(n_317), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_256), .B(n_298), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_236), .Y(n_187) );
INVx1_ASAP7_75t_SL g423 ( .A(n_188), .Y(n_423) );
AOI32xp33_ASAP7_75t_L g454 ( .A1(n_188), .A2(n_436), .A3(n_455), .B1(n_456), .B2(n_457), .Y(n_454) );
AND2x2_ASAP7_75t_L g456 ( .A(n_188), .B(n_313), .Y(n_456) );
AND2x4_ASAP7_75t_SL g188 ( .A(n_189), .B(n_216), .Y(n_188) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_189), .Y(n_237) );
INVx5_ASAP7_75t_L g316 ( .A(n_189), .Y(n_316) );
OR2x2_ASAP7_75t_L g323 ( .A(n_189), .B(n_315), .Y(n_323) );
INVx2_ASAP7_75t_L g328 ( .A(n_189), .Y(n_328) );
AND2x2_ASAP7_75t_L g340 ( .A(n_189), .B(n_217), .Y(n_340) );
AND2x2_ASAP7_75t_L g345 ( .A(n_189), .B(n_227), .Y(n_345) );
OR2x2_ASAP7_75t_L g352 ( .A(n_189), .B(n_239), .Y(n_352) );
AND2x4_ASAP7_75t_L g361 ( .A(n_189), .B(n_228), .Y(n_361) );
O2A1O1Ixp33_ASAP7_75t_SL g403 ( .A1(n_189), .A2(n_319), .B(n_354), .C(n_392), .Y(n_403) );
OR2x6_ASAP7_75t_L g189 ( .A(n_190), .B(n_194), .Y(n_189) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_191), .Y(n_225) );
AND2x2_ASAP7_75t_SL g191 ( .A(n_192), .B(n_193), .Y(n_191) );
AND2x4_ASAP7_75t_L g215 ( .A(n_192), .B(n_193), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_203), .B(n_215), .Y(n_194) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_202), .Y(n_196) );
INVx1_ASAP7_75t_L g280 ( .A(n_197), .Y(n_280) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_200), .Y(n_197) );
AND2x6_ASAP7_75t_L g211 ( .A(n_198), .B(n_206), .Y(n_211) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x4_ASAP7_75t_L g213 ( .A(n_200), .B(n_208), .Y(n_213) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx5_ASAP7_75t_L g214 ( .A(n_202), .Y(n_214) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_204), .Y(n_491) );
AND2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_207), .Y(n_204) );
BUFx3_ASAP7_75t_L g249 ( .A(n_205), .Y(n_249) );
INVx2_ASAP7_75t_L g254 ( .A(n_206), .Y(n_254) );
AND2x4_ASAP7_75t_L g251 ( .A(n_207), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g248 ( .A(n_208), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_212), .B(n_214), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_214), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_214), .A2(n_232), .B(n_233), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_214), .A2(n_263), .B(n_264), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_214), .A2(n_286), .B(n_287), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_214), .A2(n_294), .B(n_295), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_215), .B(n_270), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_215), .B(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_215), .B(n_275), .Y(n_274) );
NOR3xp33_ASAP7_75t_L g278 ( .A(n_215), .B(n_279), .C(n_280), .Y(n_278) );
INVx3_ASAP7_75t_SL g353 ( .A(n_216), .Y(n_353) );
AND2x2_ASAP7_75t_L g399 ( .A(n_216), .B(n_316), .Y(n_399) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_227), .Y(n_216) );
AND2x2_ASAP7_75t_L g238 ( .A(n_217), .B(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g330 ( .A(n_217), .B(n_228), .Y(n_330) );
AND2x2_ASAP7_75t_L g334 ( .A(n_217), .B(n_313), .Y(n_334) );
INVx1_ASAP7_75t_L g360 ( .A(n_217), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_217), .B(n_228), .Y(n_382) );
INVx2_ASAP7_75t_L g386 ( .A(n_217), .Y(n_386) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_217), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_217), .B(n_316), .Y(n_463) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_224), .B(n_226), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_223), .Y(n_218) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_224), .A2(n_229), .B(n_235), .Y(n_228) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_224), .A2(n_229), .B(n_235), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_225), .Y(n_224) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_225), .A2(n_284), .B(n_288), .Y(n_283) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g397 ( .A(n_228), .B(n_239), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_234), .Y(n_229) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx1_ASAP7_75t_L g407 ( .A(n_237), .Y(n_407) );
NAND2xp33_ASAP7_75t_SL g432 ( .A(n_237), .B(n_324), .Y(n_432) );
AND2x2_ASAP7_75t_L g474 ( .A(n_238), .B(n_316), .Y(n_474) );
AND2x2_ASAP7_75t_L g385 ( .A(n_239), .B(n_386), .Y(n_385) );
BUFx2_ASAP7_75t_L g448 ( .A(n_239), .Y(n_448) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
AOI21x1_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_244), .B(n_255), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_242), .A2(n_260), .B(n_261), .Y(n_259) );
BUFx4f_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx3_ASAP7_75t_L g277 ( .A(n_243), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_250), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_246), .A2(n_251), .B1(n_269), .B2(n_271), .Y(n_268) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
INVx1_ASAP7_75t_L g510 ( .A(n_247), .Y(n_510) );
INVx1_ASAP7_75t_L g509 ( .A(n_249), .Y(n_509) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_256), .A2(n_339), .B1(n_441), .B2(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_281), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_257), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_257), .B(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g257 ( .A(n_258), .B(n_266), .Y(n_257) );
INVx2_ASAP7_75t_L g304 ( .A(n_258), .Y(n_304) );
OR2x2_ASAP7_75t_L g308 ( .A(n_258), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_258), .B(n_321), .Y(n_326) );
AND2x4_ASAP7_75t_SL g336 ( .A(n_258), .B(n_267), .Y(n_336) );
OR2x2_ASAP7_75t_L g343 ( .A(n_258), .B(n_283), .Y(n_343) );
OR2x2_ASAP7_75t_L g355 ( .A(n_258), .B(n_267), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_258), .B(n_283), .Y(n_369) );
INVx1_ASAP7_75t_L g374 ( .A(n_258), .Y(n_374) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_258), .Y(n_392) );
AND2x2_ASAP7_75t_L g455 ( .A(n_258), .B(n_375), .Y(n_455) );
INVx2_ASAP7_75t_L g459 ( .A(n_258), .Y(n_459) );
OR2x2_ASAP7_75t_L g466 ( .A(n_258), .B(n_356), .Y(n_466) );
OR2x2_ASAP7_75t_L g488 ( .A(n_258), .B(n_489), .Y(n_488) );
OR2x6_ASAP7_75t_L g258 ( .A(n_259), .B(n_265), .Y(n_258) );
AND2x2_ASAP7_75t_L g305 ( .A(n_266), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_266), .B(n_289), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_266), .B(n_365), .Y(n_427) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g324 ( .A(n_267), .Y(n_324) );
AND2x4_ASAP7_75t_L g375 ( .A(n_267), .B(n_376), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_267), .B(n_320), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_267), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_267), .B(n_309), .Y(n_468) );
AND2x4_ASAP7_75t_L g267 ( .A(n_268), .B(n_273), .Y(n_267) );
INVx4_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI21x1_ASAP7_75t_L g290 ( .A1(n_277), .A2(n_291), .B(n_297), .Y(n_290) );
AND2x2_ASAP7_75t_L g335 ( .A(n_281), .B(n_336), .Y(n_335) );
AO221x1_ASAP7_75t_L g409 ( .A1(n_281), .A2(n_324), .B1(n_355), .B2(n_410), .C(n_411), .Y(n_409) );
OAI322xp33_ASAP7_75t_L g461 ( .A1(n_281), .A2(n_381), .A3(n_462), .B1(n_464), .B2(n_465), .C1(n_466), .C2(n_467), .Y(n_461) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_289), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx3_ASAP7_75t_L g303 ( .A(n_283), .Y(n_303) );
INVx2_ASAP7_75t_L g309 ( .A(n_283), .Y(n_309) );
AND2x2_ASAP7_75t_L g321 ( .A(n_283), .B(n_289), .Y(n_321) );
INVx1_ASAP7_75t_L g366 ( .A(n_283), .Y(n_366) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_283), .Y(n_422) );
INVx1_ASAP7_75t_L g306 ( .A(n_289), .Y(n_306) );
OR2x2_ASAP7_75t_L g356 ( .A(n_289), .B(n_309), .Y(n_356) );
INVx2_ASAP7_75t_L g376 ( .A(n_289), .Y(n_376) );
INVx1_ASAP7_75t_L g429 ( .A(n_289), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_289), .B(n_459), .Y(n_458) );
INVx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_296), .Y(n_291) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI21xp33_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_307), .B(n_310), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_300), .A2(n_339), .B1(n_341), .B2(n_345), .C(n_346), .Y(n_338) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .Y(n_301) );
NOR2x1p5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g425 ( .A(n_304), .Y(n_425) );
INVx1_ASAP7_75t_SL g344 ( .A(n_305), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_305), .A2(n_450), .B(n_452), .Y(n_449) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_306), .Y(n_349) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_309), .Y(n_412) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
OAI211xp5_ASAP7_75t_L g387 ( .A1(n_312), .A2(n_388), .B(n_393), .C(n_404), .Y(n_387) );
OR2x2_ASAP7_75t_L g477 ( .A(n_312), .B(n_382), .Y(n_477) );
AND2x2_ASAP7_75t_L g479 ( .A(n_312), .B(n_345), .Y(n_479) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g319 ( .A(n_313), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g381 ( .A(n_313), .B(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g419 ( .A(n_313), .B(n_386), .Y(n_419) );
OA33x2_ASAP7_75t_L g426 ( .A1(n_313), .A2(n_343), .A3(n_427), .B1(n_428), .B2(n_430), .B3(n_432), .Y(n_426) );
OR2x2_ASAP7_75t_L g437 ( .A(n_313), .B(n_422), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_313), .B(n_361), .Y(n_451) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g339 ( .A(n_315), .B(n_340), .Y(n_339) );
AOI22xp33_ASAP7_75t_SL g388 ( .A1(n_315), .A2(n_345), .B1(n_389), .B2(n_390), .Y(n_388) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_316), .B(n_396), .C(n_429), .Y(n_428) );
AOI322xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_322), .A3(n_324), .B1(n_325), .B2(n_327), .C1(n_331), .C2(n_335), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g424 ( .A(n_320), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
A2O1A1Ixp33_ASAP7_75t_L g379 ( .A1(n_321), .A2(n_336), .B(n_380), .C(n_383), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_322), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
NAND4xp25_ASAP7_75t_SL g443 ( .A(n_323), .B(n_352), .C(n_444), .D(n_446), .Y(n_443) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx2_ASAP7_75t_L g333 ( .A(n_328), .Y(n_333) );
OR2x2_ASAP7_75t_L g378 ( .A(n_328), .B(n_330), .Y(n_378) );
AND2x2_ASAP7_75t_L g447 ( .A(n_329), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g452 ( .A(n_333), .B(n_447), .Y(n_452) );
BUFx2_ASAP7_75t_L g445 ( .A(n_334), .Y(n_445) );
INVx1_ASAP7_75t_SL g475 ( .A(n_335), .Y(n_475) );
AND2x4_ASAP7_75t_L g411 ( .A(n_336), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g464 ( .A(n_336), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_357), .C(n_379), .Y(n_337) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_SL g401 ( .A(n_343), .Y(n_401) );
OAI211xp5_ASAP7_75t_L g469 ( .A1(n_343), .A2(n_470), .B(n_471), .C(n_480), .Y(n_469) );
OR2x2_ASAP7_75t_L g391 ( .A(n_344), .B(n_392), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_350), .B1(n_353), .B2(n_354), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_348), .B(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_351), .B(n_408), .Y(n_490) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g465 ( .A(n_352), .B(n_353), .Y(n_465) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g410 ( .A(n_356), .Y(n_410) );
AOI222xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_362), .B1(n_367), .B2(n_371), .C1(n_372), .C2(n_377), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_360), .Y(n_371) );
AND2x2_ASAP7_75t_L g418 ( .A(n_361), .B(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_361), .A2(n_434), .B1(n_439), .B2(n_443), .Y(n_433) );
INVx2_ASAP7_75t_SL g486 ( .A(n_361), .Y(n_486) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g442 ( .A(n_366), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_366), .B(n_429), .Y(n_489) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g402 ( .A(n_370), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_372), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g440 ( .A(n_374), .Y(n_440) );
AND2x2_ASAP7_75t_SL g441 ( .A(n_375), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g483 ( .A(n_375), .B(n_412), .Y(n_483) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g408 ( .A(n_382), .Y(n_408) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g487 ( .A(n_385), .Y(n_487) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_386), .Y(n_431) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_398), .B(n_400), .C(n_403), .Y(n_393) );
AND2x2_ASAP7_75t_SL g394 ( .A(n_395), .B(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g438 ( .A(n_400), .Y(n_438) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_409), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_407), .B(n_408), .Y(n_406) );
NOR3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_453), .C(n_469), .Y(n_413) );
NAND3xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_433), .C(n_449), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .B1(n_423), .B2(n_424), .C(n_426), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_435), .B(n_438), .Y(n_434) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g462 ( .A(n_448), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g470 ( .A(n_452), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_460), .Y(n_453) );
INVx2_ASAP7_75t_L g476 ( .A(n_455), .Y(n_476) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g467 ( .A(n_458), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI221xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_475), .B1(n_476), .B2(n_477), .C(n_478), .Y(n_472) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B1(n_488), .B2(n_490), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
OAI222xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B1(n_495), .B2(n_501), .C1(n_503), .C2(n_506), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
INVxp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
endmodule