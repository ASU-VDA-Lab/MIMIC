module fake_jpeg_13936_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_21),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_27),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_65),
.Y(n_77)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_20),
.B(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_1),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_80),
.B1(n_45),
.B2(n_77),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_54),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_55),
.B1(n_44),
.B2(n_53),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_52),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_92),
.Y(n_103)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_6),
.Y(n_107)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_98),
.Y(n_99)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_3),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_23),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_95),
.C(n_7),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_40),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_49),
.C(n_22),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_25),
.Y(n_96)
);

NOR2x1_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_97),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_2),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_101),
.Y(n_125)
);

NOR2xp67_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_4),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_5),
.Y(n_105)
);

AO22x1_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_114),
.B1(n_115),
.B2(n_15),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_5),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_111),
.B(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_6),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_7),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_8),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_8),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_121),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_96),
.B1(n_89),
.B2(n_83),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_108),
.B1(n_30),
.B2(n_31),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_10),
.B(n_12),
.C(n_14),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_111),
.C(n_113),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_107),
.B(n_103),
.C(n_104),
.D(n_99),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_127),
.A2(n_117),
.B1(n_124),
.B2(n_125),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_122),
.B1(n_118),
.B2(n_120),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_128),
.Y(n_137)
);

AOI322xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_128),
.A3(n_130),
.B1(n_134),
.B2(n_131),
.C1(n_127),
.C2(n_28),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_SL g139 ( 
.A(n_138),
.B(n_32),
.C(n_33),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_34),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_38),
.Y(n_141)
);


endmodule