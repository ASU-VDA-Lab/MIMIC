module fake_jpeg_22725_n_86 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_11),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_2),
.B(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_3),
.B(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_65)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_51),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_41),
.C(n_25),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_47),
.B(n_50),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

HAxp5_ASAP7_75t_SL g50 ( 
.A(n_30),
.B(n_40),
.CON(n_50),
.SN(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_28),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_23),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_36),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_68),
.Y(n_73)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_53),
.B(n_58),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.C(n_71),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_57),
.C(n_58),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_79),
.B(n_78),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_56),
.C(n_59),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_49),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_82),
.B(n_47),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_65),
.C(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_66),
.Y(n_86)
);


endmodule