module fake_jpeg_17314_n_262 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_44),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_32),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx12f_ASAP7_75t_SL g42 ( 
.A(n_18),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_29),
.B1(n_21),
.B2(n_18),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_44),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_59),
.Y(n_102)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_26),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_17),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_69),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_1),
.B(n_2),
.Y(n_95)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_71),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_21),
.B1(n_18),
.B2(n_33),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_25),
.B1(n_19),
.B2(n_23),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_33),
.Y(n_69)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx6f_ASAP7_75t_SL g83 ( 
.A(n_73),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_75),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_18),
.B(n_34),
.C(n_19),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_SL g118 ( 
.A(n_76),
.B(n_28),
.C(n_35),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_21),
.B1(n_41),
.B2(n_45),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_87),
.B1(n_96),
.B2(n_71),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_78),
.B(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_91),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_45),
.B1(n_41),
.B2(n_33),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_86),
.B1(n_88),
.B2(n_93),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_36),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_56),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_30),
.B1(n_24),
.B2(n_25),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_23),
.B1(n_20),
.B2(n_30),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_20),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_30),
.B1(n_24),
.B2(n_35),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_103),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_95),
.A2(n_60),
.B1(n_58),
.B2(n_73),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_24),
.B1(n_32),
.B2(n_35),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_24),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_72),
.Y(n_116)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_106),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_126),
.B(n_105),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_121),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_116),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_117),
.B(n_122),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_102),
.C(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_134),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_28),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_13),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_123),
.B(n_102),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_133),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_2),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_111),
.B1(n_121),
.B2(n_115),
.Y(n_157)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_85),
.A2(n_43),
.A3(n_36),
.B1(n_31),
.B2(n_32),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_92),
.B(n_89),
.Y(n_149)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_132),
.Y(n_135)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_43),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_136),
.A2(n_149),
.B(n_110),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_77),
.B1(n_84),
.B2(n_80),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_142),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_84),
.B1(n_85),
.B2(n_96),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_95),
.B1(n_84),
.B2(n_99),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_99),
.B1(n_82),
.B2(n_76),
.Y(n_142)
);

OR2x6_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_78),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_144),
.A2(n_126),
.B(n_116),
.C(n_112),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_143),
.Y(n_185)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_87),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_160),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_82),
.B1(n_81),
.B2(n_107),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_158),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_14),
.B(n_15),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_28),
.B1(n_8),
.B2(n_9),
.Y(n_186)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_94),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_4),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_108),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_162),
.B(n_112),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_174),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_170),
.B(n_146),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_168),
.B(n_169),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_137),
.A2(n_138),
.B(n_159),
.C(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_130),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_125),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_173),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_125),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_31),
.C(n_120),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_139),
.C(n_142),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_120),
.B1(n_133),
.B2(n_5),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_152),
.B1(n_158),
.B2(n_153),
.Y(n_203)
);

AO22x1_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_28),
.B1(n_31),
.B2(n_5),
.Y(n_178)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_151),
.B(n_3),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_180),
.B(n_185),
.Y(n_205)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_155),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_182),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_7),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_186),
.A2(n_144),
.B1(n_8),
.B2(n_10),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_144),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_SL g211 ( 
.A(n_188),
.B(n_165),
.C(n_178),
.Y(n_211)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_193),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_198),
.B1(n_165),
.B2(n_168),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_146),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_170),
.B(n_165),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_175),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_183),
.B(n_140),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_184),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_176),
.B(n_150),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_187),
.A2(n_140),
.B1(n_154),
.B2(n_135),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_163),
.B1(n_164),
.B2(n_182),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_209),
.C(n_219),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_166),
.C(n_179),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_218),
.Y(n_227)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_223),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_188),
.A2(n_187),
.B(n_191),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_215),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_191),
.A2(n_207),
.B1(n_201),
.B2(n_189),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_216),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_170),
.B(n_179),
.C(n_178),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_217),
.A2(n_222),
.B(n_221),
.C(n_211),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_170),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_209),
.B(n_194),
.CI(n_196),
.CON(n_226),
.SN(n_226)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_235),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_228),
.A2(n_205),
.B1(n_204),
.B2(n_28),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_199),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_234),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_198),
.C(n_206),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_218),
.C(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_216),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_232),
.B(n_219),
.CI(n_206),
.CON(n_237),
.SN(n_237)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_241),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_199),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_239),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_195),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_217),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_192),
.C(n_217),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_245),
.A2(n_228),
.B1(n_227),
.B2(n_11),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_234),
.A3(n_228),
.B1(n_229),
.B2(n_227),
.C1(n_233),
.C2(n_15),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_241),
.B1(n_244),
.B2(n_16),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_237),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_240),
.A2(n_228),
.B(n_13),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_251),
.B(n_7),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_242),
.A2(n_16),
.B(n_10),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_252),
.B(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_243),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_254),
.B(n_255),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_7),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_11),
.B1(n_12),
.B2(n_220),
.Y(n_258)
);

AO21x1_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_12),
.B(n_257),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_259),
.Y(n_262)
);


endmodule