module fake_jpeg_31983_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_12),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_26),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_0),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_0),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_81),
.Y(n_91)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_53),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_58),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_93),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_73),
.B1(n_62),
.B2(n_54),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_92),
.B1(n_98),
.B2(n_53),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_62),
.B1(n_54),
.B2(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_70),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_96),
.B(n_1),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_65),
.C(n_60),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_68),
.C(n_69),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_61),
.B1(n_58),
.B2(n_55),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_114),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_1),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_108),
.Y(n_124)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_110),
.B1(n_113),
.B2(n_4),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_8),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_53),
.B1(n_64),
.B2(n_71),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_64),
.B1(n_71),
.B2(n_25),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_71),
.B(n_2),
.C(n_3),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_117),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_2),
.B(n_3),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_131),
.B1(n_14),
.B2(n_17),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_29),
.A3(n_47),
.B1(n_43),
.B2(n_42),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_130),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_4),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_6),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_7),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_129),
.B(n_48),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_8),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_128),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_9),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_9),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_19),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_136),
.B(n_144),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_140),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_22),
.C(n_23),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_142),
.C(n_119),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_32),
.C(n_33),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_40),
.B1(n_35),
.B2(n_36),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_145),
.B1(n_149),
.B2(n_128),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_116),
.Y(n_144)
);

NAND2x1p5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_39),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_126),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_148),
.Y(n_150)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_142),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_154),
.B(n_135),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_155),
.A2(n_124),
.B1(n_145),
.B2(n_141),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_159),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_157),
.B(n_158),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_138),
.C(n_150),
.Y(n_158)
);

NOR2x1_ASAP7_75t_R g162 ( 
.A(n_160),
.B(n_154),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_161),
.B(n_135),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_161),
.B(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_152),
.B(n_147),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_153),
.Y(n_168)
);


endmodule