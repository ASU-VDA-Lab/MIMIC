module real_jpeg_24675_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_0),
.B(n_15),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_0),
.B(n_29),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_0),
.B(n_38),
.Y(n_152)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_2),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_2),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_2),
.B(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_2),
.B(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_2),
.B(n_87),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_3),
.B(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_3),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_3),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_3),
.B(n_118),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_6),
.B(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_6),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_6),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_6),
.B(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_6),
.B(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_6),
.B(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_7),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_7),
.B(n_29),
.Y(n_133)
);

INVx8_ASAP7_75t_SL g119 ( 
.A(n_8),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_9),
.B(n_15),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_11),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_11),
.B(n_29),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_11),
.B(n_38),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_11),
.B(n_35),
.Y(n_151)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_12),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_13),
.B(n_29),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_13),
.B(n_38),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_13),
.B(n_35),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_13),
.B(n_73),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_99),
.C(n_100),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.C(n_79),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_55),
.C(n_56),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_40),
.C(n_45),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_34),
.C(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_31),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.C(n_50),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_48),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_68),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_61),
.C(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_67),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_77),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_76),
.C(n_77),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_90),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_82),
.C(n_90),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_85),
.C(n_86),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_93),
.C(n_94),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_98),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_115),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_116),
.C(n_122),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_111),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_110),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_110),
.C(n_111),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_104),
.Y(n_109)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_109),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_111),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_113),
.CI(n_114),
.CON(n_111),
.SN(n_111)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_113),
.C(n_114),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.CI(n_121),
.CON(n_116),
.SN(n_116)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_140),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_131),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.CI(n_134),
.CON(n_131),
.SN(n_131)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_147),
.B1(n_153),
.B2(n_154),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_143),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_145),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_147),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);


endmodule