module fake_netlist_1_973_n_703 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_703);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_703;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_27), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_11), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_2), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_18), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_46), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_39), .Y(n_84) );
NOR2xp33_ASAP7_75t_L g85 ( .A(n_20), .B(n_23), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_78), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_37), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_19), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_11), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_44), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_43), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_50), .Y(n_92) );
CKINVDCx14_ASAP7_75t_R g93 ( .A(n_72), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_77), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_30), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_56), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_63), .Y(n_97) );
BUFx3_ASAP7_75t_L g98 ( .A(n_68), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_2), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_65), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_45), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_1), .Y(n_102) );
OR2x2_ASAP7_75t_L g103 ( .A(n_7), .B(n_76), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_34), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_19), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_31), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_7), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_64), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_28), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_48), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_47), .Y(n_111) );
BUFx5_ASAP7_75t_L g112 ( .A(n_17), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_3), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_16), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_35), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_1), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_8), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_12), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_60), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_52), .Y(n_121) );
BUFx8_ASAP7_75t_SL g122 ( .A(n_18), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_51), .Y(n_123) );
INVxp33_ASAP7_75t_L g124 ( .A(n_66), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_14), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_112), .Y(n_126) );
OAI21x1_ASAP7_75t_L g127 ( .A1(n_90), .A2(n_33), .B(n_74), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_112), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_98), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_98), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_90), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_112), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_112), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_104), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_112), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_123), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_112), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_123), .B(n_32), .Y(n_138) );
INVx4_ASAP7_75t_L g139 ( .A(n_112), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_79), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_112), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
OR2x6_ASAP7_75t_L g144 ( .A(n_103), .B(n_29), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_86), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_122), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_94), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_124), .B(n_0), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_95), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_97), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_101), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_106), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_109), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_113), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_82), .B(n_0), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_116), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_88), .B(n_3), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_125), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_125), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_92), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_103), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_80), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_111), .B(n_91), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_89), .B(n_4), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_99), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_102), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_162), .B(n_87), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_163), .B(n_114), .Y(n_171) );
NOR2x1p5_ASAP7_75t_L g172 ( .A(n_146), .B(n_107), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_163), .B(n_107), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_159), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_134), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_131), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_131), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_131), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_129), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_131), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_162), .B(n_87), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_134), .B(n_108), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_129), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_159), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_159), .B(n_85), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_163), .B(n_93), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_129), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_159), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_159), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_134), .B(n_91), .Y(n_193) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_148), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_163), .A2(n_119), .B1(n_115), .B2(n_89), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_136), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_163), .B(n_118), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_160), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_129), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_160), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_161), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_165), .B(n_108), .Y(n_202) );
OAI21xp33_ASAP7_75t_L g203 ( .A1(n_142), .A2(n_121), .B(n_100), .Y(n_203) );
OAI21xp33_ASAP7_75t_L g204 ( .A1(n_142), .A2(n_110), .B(n_118), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_148), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_136), .Y(n_206) );
INVx4_ASAP7_75t_L g207 ( .A(n_144), .Y(n_207) );
INVx8_ASAP7_75t_L g208 ( .A(n_144), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_144), .Y(n_209) );
INVx4_ASAP7_75t_SL g210 ( .A(n_138), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_148), .B(n_105), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_136), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_165), .B(n_120), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_145), .B(n_120), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_144), .A2(n_117), .B1(n_81), .B2(n_6), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_136), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_145), .B(n_147), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_144), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_144), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_147), .B(n_117), .Y(n_220) );
INVxp67_ASAP7_75t_L g221 ( .A(n_156), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_136), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_136), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_173), .B(n_168), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_215), .A2(n_156), .B1(n_153), .B2(n_154), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_208), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_208), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_176), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_208), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_189), .B(n_153), .Y(n_230) );
NOR2x1p5_ASAP7_75t_L g231 ( .A(n_220), .B(n_146), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_197), .Y(n_232) );
INVxp67_ASAP7_75t_L g233 ( .A(n_214), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_182), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_189), .B(n_154), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_208), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_191), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_191), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_197), .B(n_156), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_207), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_194), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_207), .A2(n_138), .B1(n_152), .B2(n_150), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_182), .Y(n_243) );
NOR2xp67_ASAP7_75t_L g244 ( .A(n_221), .B(n_150), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_205), .B(n_166), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_211), .B(n_171), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_171), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_199), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_198), .A2(n_168), .B(n_161), .C(n_166), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_171), .B(n_152), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_199), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_185), .B(n_164), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_207), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_200), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_201), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_191), .Y(n_256) );
INVx4_ASAP7_75t_L g257 ( .A(n_209), .Y(n_257) );
HB1xp67_ASAP7_75t_SL g258 ( .A(n_220), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_169), .B(n_152), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_174), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_209), .B(n_164), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_209), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_181), .Y(n_263) );
AOI211xp5_ASAP7_75t_L g264 ( .A1(n_220), .A2(n_164), .B(n_155), .C(n_157), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_187), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_192), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_193), .B(n_150), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_211), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_184), .B(n_152), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_202), .B(n_150), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_217), .B(n_150), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_204), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_188), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_181), .Y(n_274) );
NOR2xp67_ASAP7_75t_L g275 ( .A(n_213), .B(n_155), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_203), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_188), .B(n_151), .Y(n_277) );
INVx5_ASAP7_75t_L g278 ( .A(n_218), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_188), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_188), .Y(n_280) );
INVx3_ASAP7_75t_SL g281 ( .A(n_218), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_181), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_188), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_218), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_195), .B(n_157), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_188), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_226), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_238), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_233), .A2(n_219), .B1(n_172), .B2(n_81), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_225), .A2(n_219), .B1(n_138), .B2(n_151), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_228), .Y(n_291) );
INVx6_ASAP7_75t_L g292 ( .A(n_227), .Y(n_292) );
INVx4_ASAP7_75t_L g293 ( .A(n_227), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_238), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_226), .B(n_219), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_256), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_246), .B(n_210), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_237), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_227), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_246), .B(n_210), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_230), .A2(n_127), .B(n_223), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_257), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_228), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_237), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_257), .Y(n_305) );
INVx4_ASAP7_75t_L g306 ( .A(n_227), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_239), .B(n_210), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_258), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_227), .Y(n_309) );
INVx5_ASAP7_75t_L g310 ( .A(n_229), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_237), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_265), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_257), .Y(n_313) );
BUFx8_ASAP7_75t_L g314 ( .A(n_239), .Y(n_314) );
OR2x6_ASAP7_75t_SL g315 ( .A(n_245), .B(n_210), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_239), .B(n_149), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_235), .A2(n_127), .B(n_222), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_234), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_231), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_229), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_268), .A2(n_138), .B1(n_155), .B2(n_157), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_275), .A2(n_138), .B1(n_149), .B2(n_151), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_234), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_243), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_229), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_232), .B(n_139), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_244), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_253), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_224), .B(n_139), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_253), .Y(n_330) );
INVx5_ASAP7_75t_L g331 ( .A(n_229), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_243), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_229), .A2(n_149), .B1(n_158), .B2(n_139), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_241), .A2(n_285), .B1(n_264), .B2(n_247), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_248), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_236), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_236), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_248), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_261), .A2(n_138), .B1(n_133), .B2(n_126), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_236), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_301), .A2(n_259), .B(n_269), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_287), .B(n_245), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_317), .A2(n_277), .B(n_242), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_288), .Y(n_344) );
INVx6_ASAP7_75t_L g345 ( .A(n_310), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_290), .A2(n_236), .B1(n_250), .B2(n_280), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_325), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_290), .A2(n_236), .B1(n_273), .B2(n_280), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_288), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_314), .A2(n_273), .B1(n_283), .B2(n_286), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_294), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_287), .B(n_249), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_334), .B(n_252), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_314), .A2(n_267), .B1(n_278), .B2(n_261), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_303), .B(n_271), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_312), .Y(n_356) );
NOR2xp67_ASAP7_75t_L g357 ( .A(n_310), .B(n_278), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_294), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_312), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_314), .Y(n_360) );
AOI222xp33_ASAP7_75t_L g361 ( .A1(n_291), .A2(n_255), .B1(n_254), .B2(n_260), .C1(n_266), .C2(n_265), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_329), .B(n_261), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_310), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_325), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_329), .B(n_281), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_310), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_296), .Y(n_367) );
INVxp33_ASAP7_75t_L g368 ( .A(n_289), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_296), .A2(n_270), .B(n_279), .Y(n_369) );
CKINVDCx16_ASAP7_75t_R g370 ( .A(n_315), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g371 ( .A1(n_308), .A2(n_278), .B1(n_253), .B2(n_284), .Y(n_371) );
NOR2xp67_ASAP7_75t_L g372 ( .A(n_310), .B(n_278), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_310), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_291), .A2(n_281), .B1(n_278), .B2(n_284), .Y(n_374) );
AO22x1_ASAP7_75t_L g375 ( .A1(n_331), .A2(n_138), .B1(n_272), .B2(n_253), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_368), .A2(n_327), .B1(n_319), .B2(n_316), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_359), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_361), .A2(n_295), .B1(n_319), .B2(n_321), .Y(n_378) );
AOI21x1_ASAP7_75t_L g379 ( .A1(n_375), .A2(n_170), .B(n_190), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_361), .A2(n_295), .B1(n_276), .B2(n_322), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_355), .A2(n_339), .B1(n_307), .B2(n_333), .C(n_311), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_370), .A2(n_315), .B1(n_295), .B2(n_331), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_342), .B(n_326), .Y(n_383) );
OAI211xp5_ASAP7_75t_L g384 ( .A1(n_352), .A2(n_158), .B(n_167), .C(n_326), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_359), .B(n_331), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_360), .A2(n_299), .B1(n_336), .B2(n_311), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_359), .B(n_331), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_341), .A2(n_335), .B(n_338), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_358), .Y(n_389) );
OAI21xp5_ASAP7_75t_L g390 ( .A1(n_353), .A2(n_127), .B(n_338), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_342), .B(n_331), .Y(n_391) );
AOI222xp33_ASAP7_75t_L g392 ( .A1(n_360), .A2(n_158), .B1(n_138), .B2(n_304), .C1(n_299), .C2(n_336), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_365), .A2(n_304), .B1(n_302), .B2(n_305), .Y(n_393) );
AOI22xp33_ASAP7_75t_SL g394 ( .A1(n_370), .A2(n_331), .B1(n_302), .B2(n_305), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_356), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_365), .A2(n_305), .B1(n_313), .B2(n_302), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_355), .A2(n_126), .B1(n_133), .B2(n_139), .C(n_135), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_356), .B(n_293), .Y(n_398) );
OAI21x1_ASAP7_75t_L g399 ( .A1(n_343), .A2(n_330), .B(n_328), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_358), .Y(n_400) );
AND2x4_ASAP7_75t_SL g401 ( .A(n_358), .B(n_293), .Y(n_401) );
BUFx4f_ASAP7_75t_SL g402 ( .A(n_373), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_345), .A2(n_373), .B1(n_363), .B2(n_366), .Y(n_403) );
CKINVDCx11_ASAP7_75t_R g404 ( .A(n_344), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_378), .A2(n_354), .B1(n_362), .B2(n_367), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_376), .A2(n_350), .B1(n_367), .B2(n_371), .C(n_369), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_378), .A2(n_362), .B1(n_344), .B2(n_349), .Y(n_407) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_404), .B(n_167), .C(n_143), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_400), .B(n_349), .Y(n_409) );
AO21x2_ASAP7_75t_L g410 ( .A1(n_399), .A2(n_346), .B(n_351), .Y(n_410) );
INVx2_ASAP7_75t_SL g411 ( .A(n_401), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_382), .A2(n_351), .B1(n_138), .B2(n_366), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_383), .A2(n_167), .B1(n_136), .B2(n_140), .C(n_143), .Y(n_413) );
OA21x2_ASAP7_75t_L g414 ( .A1(n_399), .A2(n_170), .B(n_186), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_380), .A2(n_363), .B1(n_357), .B2(n_372), .C(n_167), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_385), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_380), .A2(n_345), .B1(n_348), .B2(n_372), .Y(n_417) );
AOI222xp33_ASAP7_75t_L g418 ( .A1(n_382), .A2(n_138), .B1(n_357), .B2(n_375), .C1(n_167), .C2(n_140), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_392), .B(n_167), .C(n_143), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_400), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_377), .B(n_389), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_386), .A2(n_167), .B1(n_313), .B2(n_320), .C(n_337), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_377), .B(n_364), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_385), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_395), .A2(n_143), .B1(n_140), .B2(n_133), .C(n_126), .Y(n_425) );
NAND2x1p5_ASAP7_75t_L g426 ( .A(n_387), .B(n_364), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_377), .B(n_364), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_391), .A2(n_345), .B1(n_293), .B2(n_306), .Y(n_428) );
AOI33xp33_ASAP7_75t_L g429 ( .A1(n_395), .A2(n_141), .A3(n_135), .B1(n_128), .B2(n_132), .B3(n_137), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_393), .A2(n_313), .B1(n_320), .B2(n_337), .C(n_298), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_402), .A2(n_345), .B1(n_374), .B2(n_306), .Y(n_431) );
AND2x4_ASAP7_75t_SL g432 ( .A(n_387), .B(n_306), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_389), .B(n_398), .Y(n_433) );
OAI221xp5_ASAP7_75t_SL g434 ( .A1(n_384), .A2(n_298), .B1(n_126), .B2(n_133), .C(n_141), .Y(n_434) );
OAI33xp33_ASAP7_75t_L g435 ( .A1(n_389), .A2(n_183), .A3(n_223), .B1(n_222), .B2(n_212), .B3(n_206), .Y(n_435) );
OAI21xp33_ASAP7_75t_L g436 ( .A1(n_392), .A2(n_133), .B(n_126), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_396), .A2(n_140), .B1(n_143), .B2(n_330), .C(n_328), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_432), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_433), .B(n_398), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_421), .Y(n_440) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_407), .A2(n_390), .B1(n_401), .B2(n_381), .C1(n_140), .C2(n_143), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_420), .B(n_401), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_421), .Y(n_443) );
OAI21xp33_ASAP7_75t_L g444 ( .A1(n_408), .A2(n_143), .B(n_140), .Y(n_444) );
AND3x2_ASAP7_75t_L g445 ( .A(n_416), .B(n_390), .C(n_394), .Y(n_445) );
AOI211xp5_ASAP7_75t_L g446 ( .A1(n_415), .A2(n_140), .B(n_130), .C(n_129), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_420), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_409), .B(n_403), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_433), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_432), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_409), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_424), .B(n_364), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_423), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_406), .A2(n_139), .B1(n_397), .B2(n_137), .C(n_132), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_423), .B(n_347), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_411), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_411), .B(n_4), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_405), .B(n_388), .Y(n_458) );
OAI33xp33_ASAP7_75t_L g459 ( .A1(n_417), .A2(n_132), .A3(n_137), .B1(n_128), .B2(n_183), .B3(n_180), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_427), .B(n_5), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_427), .B(n_5), .Y(n_461) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_419), .A2(n_347), .B1(n_292), .B2(n_340), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_435), .A2(n_347), .B(n_325), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_422), .A2(n_309), .B1(n_129), .B2(n_130), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_426), .B(n_6), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_426), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_414), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_434), .B(n_128), .C(n_379), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_426), .B(n_347), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_429), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_429), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_410), .B(n_8), .Y(n_472) );
NAND3xp33_ASAP7_75t_SL g473 ( .A(n_418), .B(n_9), .C(n_10), .Y(n_473) );
NAND3xp33_ASAP7_75t_SL g474 ( .A(n_412), .B(n_9), .C(n_10), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_430), .Y(n_475) );
NAND2xp33_ASAP7_75t_R g476 ( .A(n_414), .B(n_379), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_410), .B(n_347), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_431), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_428), .B(n_12), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_410), .B(n_13), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_414), .B(n_13), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_437), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_413), .B(n_340), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_425), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_447), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_443), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_451), .B(n_14), .Y(n_487) );
OAI31xp33_ASAP7_75t_L g488 ( .A1(n_438), .A2(n_436), .A3(n_300), .B(n_297), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_440), .B(n_130), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_443), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_449), .B(n_15), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_440), .B(n_130), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_440), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_467), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_453), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_449), .B(n_130), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_467), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_450), .B(n_15), .Y(n_498) );
BUFx2_ASAP7_75t_L g499 ( .A(n_450), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_472), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_477), .B(n_130), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_465), .A2(n_292), .B1(n_340), .B2(n_325), .Y(n_502) );
OAI31xp33_ASAP7_75t_L g503 ( .A1(n_465), .A2(n_300), .A3(n_297), .B(n_309), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_472), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_455), .B(n_130), .Y(n_505) );
BUFx2_ASAP7_75t_SL g506 ( .A(n_442), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_480), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_477), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_474), .B(n_186), .C(n_190), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_457), .B(n_16), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_439), .B(n_17), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_442), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_481), .Y(n_513) );
INVxp33_ASAP7_75t_L g514 ( .A(n_442), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_446), .A2(n_340), .B(n_325), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_481), .Y(n_516) );
INVxp67_ASAP7_75t_SL g517 ( .A(n_439), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_455), .B(n_21), .Y(n_518) );
NAND2x1p5_ASAP7_75t_L g519 ( .A(n_456), .B(n_340), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_448), .B(n_22), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_448), .B(n_24), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_458), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_478), .B(n_335), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_456), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_456), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_452), .B(n_25), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_452), .B(n_26), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_460), .Y(n_528) );
AOI211xp5_ASAP7_75t_L g529 ( .A1(n_473), .A2(n_180), .B(n_177), .C(n_178), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_475), .A2(n_330), .B1(n_328), .B2(n_292), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_461), .B(n_332), .Y(n_531) );
NOR3xp33_ASAP7_75t_L g532 ( .A(n_479), .B(n_178), .C(n_175), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_469), .B(n_36), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_469), .B(n_38), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_470), .A2(n_471), .B1(n_482), .B2(n_441), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_466), .B(n_40), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_463), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_483), .Y(n_538) );
OAI31xp33_ASAP7_75t_L g539 ( .A1(n_444), .A2(n_300), .A3(n_297), .B(n_179), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_483), .B(n_41), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_445), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_483), .B(n_42), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_517), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_506), .B(n_462), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_508), .B(n_464), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_486), .B(n_464), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_485), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_506), .B(n_484), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_495), .B(n_468), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_493), .B(n_49), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_512), .B(n_53), .Y(n_551) );
NOR2x1_ASAP7_75t_R g552 ( .A(n_499), .B(n_292), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_485), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_498), .A2(n_454), .B(n_459), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_508), .B(n_196), .Y(n_555) );
NAND2xp33_ASAP7_75t_L g556 ( .A(n_540), .B(n_476), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_495), .B(n_175), .Y(n_557) );
NOR2x1_ASAP7_75t_L g558 ( .A(n_499), .B(n_476), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_486), .Y(n_559) );
XNOR2xp5_ASAP7_75t_L g560 ( .A(n_541), .B(n_54), .Y(n_560) );
OAI211xp5_ASAP7_75t_L g561 ( .A1(n_541), .A2(n_206), .B(n_212), .C(n_179), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_490), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_522), .B(n_196), .C(n_216), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_490), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_507), .B(n_177), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_507), .B(n_332), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_528), .B(n_324), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_514), .B(n_55), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_500), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_522), .B(n_324), .Y(n_570) );
AND2x2_ASAP7_75t_SL g571 ( .A(n_540), .B(n_284), .Y(n_571) );
NAND2xp33_ASAP7_75t_SL g572 ( .A(n_520), .B(n_284), .Y(n_572) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_511), .B(n_323), .C(n_318), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_505), .B(n_57), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_538), .B(n_284), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_494), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_500), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_504), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_504), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_513), .B(n_323), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_513), .B(n_318), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_505), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_493), .B(n_58), .Y(n_583) );
AND2x4_ASAP7_75t_L g584 ( .A(n_538), .B(n_59), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_487), .B(n_61), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_516), .B(n_62), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_516), .B(n_67), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_518), .Y(n_588) );
OAI31xp33_ASAP7_75t_SL g589 ( .A1(n_510), .A2(n_69), .A3(n_70), .B(n_73), .Y(n_589) );
NOR3xp33_ASAP7_75t_L g590 ( .A(n_491), .B(n_240), .C(n_251), .Y(n_590) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_542), .B(n_262), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_535), .A2(n_181), .B1(n_196), .B2(n_216), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_496), .Y(n_593) );
INVx2_ASAP7_75t_SL g594 ( .A(n_489), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_501), .B(n_75), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_501), .B(n_181), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_501), .B(n_196), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_496), .B(n_196), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_543), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_547), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_572), .A2(n_515), .B(n_542), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_569), .B(n_525), .Y(n_602) );
AOI32xp33_ASAP7_75t_L g603 ( .A1(n_556), .A2(n_521), .A3(n_520), .B1(n_527), .B2(n_526), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_553), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_577), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_578), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_588), .B(n_525), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_552), .Y(n_608) );
AO21x1_ASAP7_75t_L g609 ( .A1(n_572), .A2(n_533), .B(n_519), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_571), .A2(n_521), .B1(n_533), .B2(n_527), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_579), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_549), .B(n_524), .Y(n_612) );
XNOR2xp5_ASAP7_75t_L g613 ( .A(n_560), .B(n_518), .Y(n_613) );
NOR2x1_ASAP7_75t_L g614 ( .A(n_558), .B(n_533), .Y(n_614) );
AOI211xp5_ASAP7_75t_L g615 ( .A1(n_556), .A2(n_488), .B(n_503), .C(n_526), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_582), .B(n_524), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_595), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_559), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_571), .B(n_519), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_562), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_564), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_596), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_593), .B(n_492), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_563), .Y(n_624) );
NOR2xp67_ASAP7_75t_L g625 ( .A(n_544), .B(n_494), .Y(n_625) );
OAI222xp33_ASAP7_75t_L g626 ( .A1(n_591), .A2(n_519), .B1(n_489), .B2(n_534), .C1(n_502), .C2(n_492), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_594), .B(n_497), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_576), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_548), .B(n_523), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_594), .B(n_497), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_576), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_546), .B(n_523), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_550), .B(n_537), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_555), .Y(n_634) );
XNOR2xp5_ASAP7_75t_L g635 ( .A(n_574), .B(n_534), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_566), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_570), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_545), .B(n_537), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_545), .B(n_531), .Y(n_639) );
XOR2xp5_ASAP7_75t_L g640 ( .A(n_587), .B(n_536), .Y(n_640) );
AOI311xp33_ASAP7_75t_L g641 ( .A1(n_573), .A2(n_532), .A3(n_529), .B(n_509), .C(n_530), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_581), .Y(n_642) );
AOI22x1_ASAP7_75t_L g643 ( .A1(n_568), .A2(n_536), .B1(n_539), .B2(n_253), .Y(n_643) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_575), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_580), .B(n_216), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_573), .A2(n_590), .B1(n_554), .B2(n_592), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g647 ( .A(n_551), .Y(n_647) );
OAI22xp5_ASAP7_75t_SL g648 ( .A1(n_592), .A2(n_262), .B1(n_240), .B2(n_216), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_575), .B(n_216), .Y(n_649) );
INVxp67_ASAP7_75t_SL g650 ( .A(n_555), .Y(n_650) );
OA21x2_ASAP7_75t_L g651 ( .A1(n_567), .A2(n_263), .B(n_274), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_557), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_565), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g654 ( .A1(n_584), .A2(n_597), .B1(n_583), .B2(n_550), .Y(n_654) );
OAI22xp5_ASAP7_75t_SL g655 ( .A1(n_585), .A2(n_262), .B1(n_251), .B2(n_263), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_586), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_550), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_584), .B(n_262), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_583), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_598), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_584), .B(n_262), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_583), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_589), .A2(n_274), .B1(n_282), .B2(n_585), .C(n_590), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_561), .Y(n_664) );
BUFx8_ASAP7_75t_L g665 ( .A(n_664), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_608), .A2(n_615), .B1(n_603), .B2(n_635), .Y(n_666) );
NOR2xp67_ASAP7_75t_SL g667 ( .A(n_619), .B(n_601), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_612), .A2(n_625), .B1(n_629), .B2(n_617), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_599), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_630), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_606), .Y(n_671) );
NOR2xp67_ASAP7_75t_L g672 ( .A(n_608), .B(n_624), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_612), .A2(n_629), .B1(n_646), .B2(n_610), .Y(n_673) );
XOR2xp5_ASAP7_75t_L g674 ( .A(n_613), .B(n_640), .Y(n_674) );
NAND4xp25_ASAP7_75t_L g675 ( .A(n_641), .B(n_614), .C(n_652), .D(n_619), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g676 ( .A1(n_654), .A2(n_622), .B1(n_650), .B2(n_644), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_605), .Y(n_677) );
AOI21xp33_ASAP7_75t_SL g678 ( .A1(n_654), .A2(n_643), .B(n_647), .Y(n_678) );
OAI21xp5_ASAP7_75t_SL g679 ( .A1(n_626), .A2(n_624), .B(n_663), .Y(n_679) );
AOI211xp5_ASAP7_75t_L g680 ( .A1(n_672), .A2(n_609), .B(n_655), .C(n_653), .Y(n_680) );
AOI322xp5_ASAP7_75t_L g681 ( .A1(n_676), .A2(n_673), .A3(n_670), .B1(n_668), .B2(n_669), .C1(n_666), .C2(n_665), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_679), .A2(n_644), .B(n_633), .C(n_660), .Y(n_682) );
OAI211xp5_ASAP7_75t_L g683 ( .A1(n_678), .A2(n_660), .B(n_650), .C(n_639), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_675), .A2(n_611), .B1(n_602), .B2(n_636), .C(n_604), .Y(n_684) );
AOI211xp5_ASAP7_75t_L g685 ( .A1(n_667), .A2(n_648), .B(n_637), .C(n_656), .Y(n_685) );
AOI211xp5_ASAP7_75t_L g686 ( .A1(n_665), .A2(n_632), .B(n_642), .C(n_602), .Y(n_686) );
NAND4xp25_ASAP7_75t_SL g687 ( .A(n_674), .B(n_607), .C(n_657), .D(n_662), .Y(n_687) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_671), .B(n_651), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_681), .B(n_677), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_688), .Y(n_690) );
AOI211xp5_ASAP7_75t_SL g691 ( .A1(n_683), .A2(n_638), .B(n_645), .C(n_659), .Y(n_691) );
NAND3x1_ASAP7_75t_L g692 ( .A(n_684), .B(n_627), .C(n_658), .Y(n_692) );
NAND3xp33_ASAP7_75t_SL g693 ( .A(n_680), .B(n_661), .C(n_649), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_689), .A2(n_682), .B1(n_687), .B2(n_685), .C(n_686), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_690), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_691), .A2(n_600), .B1(n_616), .B2(n_621), .C(n_618), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_695), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_694), .A2(n_693), .B(n_692), .Y(n_698) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_697), .Y(n_699) );
OAI21xp5_ASAP7_75t_L g700 ( .A1(n_698), .A2(n_696), .B(n_633), .Y(n_700) );
OR2x2_ASAP7_75t_L g701 ( .A(n_699), .B(n_620), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_701), .A2(n_700), .B1(n_623), .B2(n_634), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_702), .A2(n_628), .B1(n_631), .B2(n_651), .C(n_282), .Y(n_703) );
endmodule