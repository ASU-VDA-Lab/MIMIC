module real_jpeg_23325_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_2),
.B(n_142),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_2),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_2),
.B(n_60),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_2),
.B(n_38),
.C(n_79),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_2),
.A2(n_61),
.B1(n_65),
.B2(n_209),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_2),
.B(n_123),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_2),
.A2(n_38),
.B1(n_40),
.B2(n_209),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_2),
.B(n_26),
.C(n_43),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_2),
.A2(n_25),
.B(n_270),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g64 ( 
.A(n_4),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_5),
.A2(n_56),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_5),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_5),
.A2(n_61),
.B1(n_65),
.B2(n_107),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_5),
.A2(n_38),
.B1(n_40),
.B2(n_107),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_5),
.A2(n_26),
.B1(n_32),
.B2(n_107),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_6),
.A2(n_61),
.B1(n_65),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_6),
.A2(n_38),
.B1(n_40),
.B2(n_83),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_6),
.A2(n_54),
.B1(n_57),
.B2(n_83),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_6),
.A2(n_26),
.B1(n_32),
.B2(n_83),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_54),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_8),
.A2(n_61),
.B1(n_65),
.B2(n_70),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_8),
.A2(n_38),
.B1(n_40),
.B2(n_70),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_8),
.A2(n_26),
.B1(n_32),
.B2(n_70),
.Y(n_240)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_37),
.B1(n_61),
.B2(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_10),
.A2(n_37),
.B1(n_71),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_10),
.A2(n_26),
.B1(n_32),
.B2(n_37),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_11),
.A2(n_38),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_26),
.B1(n_32),
.B2(n_47),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_11),
.A2(n_47),
.B1(n_61),
.B2(n_65),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_11),
.A2(n_47),
.B1(n_159),
.B2(n_338),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_12),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_12),
.A2(n_58),
.B1(n_61),
.B2(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_12),
.A2(n_38),
.B1(n_40),
.B2(n_58),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_12),
.A2(n_26),
.B1(n_32),
.B2(n_58),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_14),
.A2(n_71),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_14),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_14),
.A2(n_61),
.B1(n_65),
.B2(n_158),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_14),
.A2(n_38),
.B1(n_40),
.B2(n_158),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_14),
.A2(n_26),
.B1(n_32),
.B2(n_158),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_15),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_15),
.A2(n_33),
.B1(n_38),
.B2(n_40),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_15),
.A2(n_33),
.B1(n_61),
.B2(n_65),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_15),
.A2(n_33),
.B1(n_159),
.B2(n_338),
.Y(n_347)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_16),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_343),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_329),
.B(n_342),
.Y(n_18)
);

OAI31xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_133),
.A3(n_148),
.B(n_326),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_21),
.B(n_112),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.C(n_90),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_22),
.A2(n_74),
.B1(n_75),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_22),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_23),
.A2(n_24),
.B(n_51),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_24),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_24),
.A2(n_34),
.B1(n_35),
.B2(n_50),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_31),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_25),
.A2(n_31),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_25),
.A2(n_28),
.B1(n_95),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_25),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_25),
.A2(n_27),
.B1(n_183),
.B2(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_25),
.B(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_25),
.A2(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_45)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_27),
.Y(n_283)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_29),
.B(n_271),
.Y(n_270)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_30),
.B(n_209),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_32),
.B(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_41),
.B1(n_46),
.B2(n_48),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_36),
.A2(n_41),
.B1(n_48),
.B2(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_38),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_38),
.A2(n_40),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_38),
.B(n_277),
.Y(n_276)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_41),
.A2(n_48),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_41),
.B(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_41),
.A2(n_48),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_45),
.A2(n_86),
.B1(n_101),
.B2(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_45),
.A2(n_169),
.B(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_45),
.A2(n_205),
.B(n_243),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_45),
.B(n_209),
.Y(n_289)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_48),
.B(n_206),
.Y(n_258)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_59),
.B(n_67),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_53),
.A2(n_59),
.B1(n_109),
.B2(n_131),
.Y(n_130)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_56),
.B1(n_63),
.B2(n_66),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g184 ( 
.A1(n_55),
.A2(n_63),
.A3(n_65),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_69),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_59),
.A2(n_109),
.B1(n_131),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_59),
.A2(n_67),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_60),
.A2(n_72),
.B1(n_106),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_60),
.A2(n_72),
.B1(n_336),
.B2(n_337),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_60),
.A2(n_72),
.B1(n_337),
.B2(n_347),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_65),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_61),
.B(n_66),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_61),
.B(n_233),
.Y(n_232)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_71),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_72),
.A2(n_111),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_85),
.B(n_89),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_85),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_84),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_77),
.A2(n_78),
.B1(n_125),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_77),
.A2(n_176),
.B(n_178),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g246 ( 
.A1(n_77),
.A2(n_178),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_78),
.A2(n_103),
.B(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_78),
.A2(n_162),
.B(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_86),
.A2(n_257),
.B(n_258),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_86),
.A2(n_258),
.B(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_88),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_90),
.A2(n_91),
.B1(n_321),
.B2(n_323),
.Y(n_320)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.C(n_104),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_92),
.A2(n_93),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_94),
.A2(n_98),
.B1(n_99),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_94),
.Y(n_171)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_97),
.A2(n_167),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_102),
.B(n_104),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B(n_110),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_115),
.C(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_130),
.B2(n_132),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_127),
.C(n_130),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_122),
.A2(n_123),
.B1(n_177),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_122),
.A2(n_123),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_123),
.B(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_127),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_127),
.B(n_140),
.C(n_145),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_130),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_132),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_130),
.B(n_136),
.C(n_139),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_134),
.A2(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_147),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_135),
.B(n_147),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_141),
.Y(n_336)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_146),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_319),
.B(n_325),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_194),
.B(n_318),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_187),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_151),
.B(n_187),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_170),
.C(n_172),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_152),
.A2(n_153),
.B1(n_170),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_164),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_160),
.B2(n_161),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_160),
.C(n_164),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_159),
.Y(n_338)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_168),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_170),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_172),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_179),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_175),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_179),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_184),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_181),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_189),
.B(n_190),
.C(n_193),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_225),
.B(n_312),
.C(n_317),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_219),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_219),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_211),
.C(n_212),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_197),
.A2(n_198),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_203),
.C(n_207),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_202),
.Y(n_214)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_211),
.B(n_212),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.C(n_217),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_220),
.B(n_223),
.C(n_224),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_306),
.B(n_311),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_259),
.B(n_305),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_248),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_230),
.B(n_248),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_241),
.C(n_245),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_231),
.B(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_234),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B(n_239),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_238),
.A2(n_282),
.B(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_241),
.A2(n_245),
.B1(n_246),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_241),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_244),
.Y(n_257)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_249),
.B(n_255),
.C(n_256),
.Y(n_310)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_299),
.B(n_304),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_278),
.B(n_298),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_272),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_272),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_268),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_267),
.C(n_268),
.Y(n_303)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_269),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_276),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_287),
.B(n_297),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_285),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_285),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_292),
.B(n_296),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_290),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_303),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_310),
.Y(n_311)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_324),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_324),
.Y(n_325)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_331),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_341),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_335),
.B1(n_339),
.B2(n_340),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_333),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_339),
.C(n_341),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_349),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_348),
.Y(n_349)
);


endmodule