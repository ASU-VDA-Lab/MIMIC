module fake_jpeg_26021_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_7),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_47),
.Y(n_60)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_54),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_34),
.C(n_25),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_34),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_21),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_68),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_74),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_38),
.B1(n_44),
.B2(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_71),
.A2(n_22),
.B1(n_19),
.B2(n_30),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_25),
.B1(n_36),
.B2(n_26),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_80),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_36),
.B1(n_24),
.B2(n_26),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_96),
.B1(n_97),
.B2(n_20),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_29),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_29),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_41),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_64),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_56),
.B(n_27),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_48),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_59),
.C(n_58),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_36),
.B(n_30),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_20),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_40),
.B1(n_38),
.B2(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_43),
.B1(n_62),
.B2(n_32),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_38),
.B1(n_44),
.B2(n_46),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_103),
.B1(n_88),
.B2(n_83),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_98),
.B(n_82),
.C(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_90),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_46),
.B1(n_37),
.B2(n_22),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

AO22x1_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_37),
.B1(n_23),
.B2(n_22),
.Y(n_108)
);

AO22x1_ASAP7_75t_SL g151 ( 
.A1(n_108),
.A2(n_115),
.B1(n_59),
.B2(n_58),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_18),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_116),
.C(n_118),
.Y(n_140)
);

NAND2xp33_ASAP7_75t_R g148 ( 
.A(n_112),
.B(n_119),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_124),
.B1(n_87),
.B2(n_93),
.Y(n_146)
);

AO22x2_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_37),
.B1(n_43),
.B2(n_59),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

OR2x4_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_43),
.Y(n_119)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_73),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_73),
.Y(n_125)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_137),
.B1(n_151),
.B2(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_129),
.A2(n_153),
.B(n_27),
.Y(n_180)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_130),
.B(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_126),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_79),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_136),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_134),
.B(n_143),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_99),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_135),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_78),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_83),
.B1(n_81),
.B2(n_74),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_138),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_78),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_147),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_79),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_89),
.B(n_97),
.Y(n_153)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_77),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_112),
.B(n_102),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_156),
.A2(n_157),
.B(n_174),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_108),
.B(n_104),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_161),
.B(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_147),
.B1(n_145),
.B2(n_151),
.Y(n_201)
);

AO22x1_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_108),
.B1(n_101),
.B2(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_170),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_106),
.B1(n_120),
.B2(n_117),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_169),
.A2(n_175),
.B1(n_182),
.B2(n_154),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_179),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_91),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_176),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_18),
.B(n_19),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_106),
.B1(n_125),
.B2(n_105),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_43),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_180),
.Y(n_204)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_183),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_105),
.B1(n_92),
.B2(n_70),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_187),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_211),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_134),
.C(n_133),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_195),
.B(n_203),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_132),
.B1(n_151),
.B2(n_127),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_199),
.B1(n_201),
.B2(n_212),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_130),
.Y(n_198)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_174),
.B(n_129),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_141),
.B1(n_138),
.B2(n_154),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_205),
.A2(n_210),
.B1(n_175),
.B2(n_159),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_168),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_206),
.B(n_207),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_158),
.B(n_28),
.Y(n_207)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_208),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_92),
.B1(n_70),
.B2(n_28),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_163),
.A2(n_77),
.B1(n_58),
.B2(n_57),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_160),
.A2(n_0),
.B(n_1),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_180),
.B(n_156),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_160),
.A2(n_77),
.B1(n_57),
.B2(n_31),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_161),
.B1(n_166),
.B2(n_68),
.Y(n_240)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_56),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_222),
.A2(n_224),
.B(n_226),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_193),
.A2(n_200),
.B(n_211),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_157),
.B(n_186),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_173),
.C(n_176),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_205),
.C(n_209),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_204),
.A2(n_186),
.B(n_178),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_231),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_236),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_178),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_243),
.Y(n_265)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_216),
.B(n_166),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_244),
.Y(n_256)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

NOR4xp25_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_184),
.C(n_165),
.D(n_159),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_238),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_199),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_221),
.B1(n_218),
.B2(n_241),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_32),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_32),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_257),
.Y(n_274)
);

INVxp33_ASAP7_75t_SL g247 ( 
.A(n_223),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_218),
.C(n_209),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_259),
.C(n_264),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_251),
.B1(n_266),
.B2(n_220),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_221),
.A2(n_217),
.B1(n_197),
.B2(n_212),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_258),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_203),
.C(n_215),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_223),
.Y(n_261)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_207),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_228),
.A2(n_210),
.B1(n_197),
.B2(n_202),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_243),
.C(n_226),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_240),
.A2(n_214),
.B1(n_208),
.B2(n_191),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_255),
.A2(n_225),
.B1(n_239),
.B2(n_231),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_31),
.B1(n_8),
.B2(n_15),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_270),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_222),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_275),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_225),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_242),
.C(n_220),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_281),
.C(n_246),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_252),
.A2(n_242),
.B(n_219),
.Y(n_277)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_214),
.C(n_191),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_283),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_10),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_266),
.B1(n_261),
.B2(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_260),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_287),
.B(n_292),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_294),
.Y(n_304)
);

AO22x1_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_260),
.B1(n_251),
.B2(n_256),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_293),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_265),
.C(n_256),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_268),
.C(n_274),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_10),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_11),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_271),
.B(n_261),
.Y(n_294)
);

NOR3xp33_ASAP7_75t_SL g295 ( 
.A(n_283),
.B(n_8),
.C(n_15),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_296),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_267),
.B1(n_278),
.B2(n_281),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_268),
.C(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_300),
.B(n_309),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_310),
.C(n_289),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_35),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_307),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_35),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_286),
.A2(n_6),
.B(n_13),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_35),
.B(n_20),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_5),
.C(n_12),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_291),
.C(n_290),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_284),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_318),
.C(n_319),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_295),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_304),
.Y(n_319)
);

AOI21x1_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_13),
.B(n_8),
.Y(n_320)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_308),
.B(n_6),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_324),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_304),
.C(n_306),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_299),
.B1(n_307),
.B2(n_6),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_316),
.C(n_312),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_314),
.A2(n_0),
.B(n_1),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_4),
.Y(n_330)
);

AO21x1_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_0),
.B(n_1),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_328),
.B1(n_1),
.B2(n_2),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_329),
.B(n_322),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_322),
.C(n_323),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_0),
.C(n_2),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_2),
.C(n_3),
.Y(n_336)
);

AO22x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_3),
.B1(n_4),
.B2(n_247),
.Y(n_337)
);


endmodule