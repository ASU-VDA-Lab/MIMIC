module fake_jpeg_24150_n_260 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_245;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_114;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_9),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_40),
.B1(n_27),
.B2(n_19),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_16),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_16),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_43),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_19),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_27),
.B1(n_43),
.B2(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_50),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_22),
.B1(n_31),
.B2(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_30),
.B1(n_36),
.B2(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_20),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_23),
.B1(n_22),
.B2(n_31),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_30),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_40),
.B1(n_23),
.B2(n_37),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_67),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_58),
.Y(n_92)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_28),
.B1(n_32),
.B2(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_39),
.B1(n_32),
.B2(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_29),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_69),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_85),
.B(n_36),
.C(n_33),
.Y(n_98)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_83),
.Y(n_109)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_22),
.B1(n_31),
.B2(n_30),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_82),
.B1(n_84),
.B2(n_5),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_88),
.Y(n_100)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_87),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_55),
.B1(n_48),
.B2(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_44),
.B(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_95),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_56),
.B(n_60),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_103),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_85),
.B(n_79),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_63),
.B1(n_58),
.B2(n_75),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_87),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_1),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_5),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_76),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_111),
.B1(n_72),
.B2(n_59),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_120),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_88),
.C(n_75),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_124),
.C(n_135),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_109),
.B(n_101),
.Y(n_151)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_57),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_121),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_132),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_123),
.A2(n_138),
.B1(n_119),
.B2(n_118),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_70),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_68),
.B(n_66),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_128),
.B(n_134),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_92),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_94),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_97),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_130),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_137),
.B1(n_100),
.B2(n_108),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_6),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_78),
.C(n_71),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_140),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_64),
.B1(n_7),
.B2(n_10),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_96),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_96),
.B(n_11),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_112),
.C(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_142),
.B(n_146),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_145),
.A2(n_151),
.B1(n_157),
.B2(n_166),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_150),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_98),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_155),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_161),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_101),
.B1(n_111),
.B2(n_106),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_94),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_139),
.C(n_117),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_185),
.C(n_186),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_124),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_171),
.A2(n_150),
.B(n_156),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_141),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_175),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_134),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_174),
.B(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_122),
.A3(n_120),
.B1(n_134),
.B2(n_126),
.C1(n_137),
.C2(n_93),
.Y(n_178)
);

BUFx4f_ASAP7_75t_SL g182 ( 
.A(n_163),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_144),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_183),
.A2(n_149),
.B1(n_141),
.B2(n_152),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_93),
.B1(n_106),
.B2(n_113),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_184),
.A2(n_147),
.B1(n_157),
.B2(n_161),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_93),
.C(n_106),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_105),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_142),
.B(n_143),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_191),
.B(n_198),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_197),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_188),
.B1(n_184),
.B2(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_176),
.B(n_148),
.CI(n_167),
.CON(n_199),
.SN(n_199)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_203),
.B(n_204),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_151),
.C(n_159),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_185),
.C(n_169),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_153),
.B(n_13),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_105),
.Y(n_204)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_217),
.C(n_196),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_212),
.A2(n_193),
.B1(n_181),
.B2(n_201),
.Y(n_232)
);

BUFx12_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_175),
.B1(n_168),
.B2(n_173),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_199),
.B1(n_193),
.B2(n_205),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_181),
.C(n_171),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_171),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_206),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_177),
.C(n_183),
.Y(n_220)
);

OAI321xp33_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_193),
.A3(n_203),
.B1(n_199),
.B2(n_205),
.C(n_168),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_230),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_195),
.B1(n_192),
.B2(n_190),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_224),
.A2(n_212),
.B1(n_218),
.B2(n_211),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_SL g226 ( 
.A(n_219),
.B(n_182),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_216),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_201),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_227),
.Y(n_239)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_206),
.C(n_197),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_232),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_214),
.B1(n_216),
.B2(n_209),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_237),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_224),
.B(n_222),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_230),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_245),
.B(n_239),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_240),
.A2(n_223),
.B(n_229),
.Y(n_244)
);

AOI21x1_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_235),
.B(n_236),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_180),
.B(n_213),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_233),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_247),
.C(n_180),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_248),
.A2(n_249),
.B(n_251),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_114),
.C(n_14),
.Y(n_255)
);

NOR2x1_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_208),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_251),
.A2(n_243),
.B(n_114),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_255),
.Y(n_257)
);

AOI221xp5_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_252),
.B1(n_114),
.B2(n_15),
.C(n_14),
.Y(n_256)
);

INVxp33_ASAP7_75t_SL g258 ( 
.A(n_256),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_257),
.B(n_14),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_12),
.B(n_15),
.Y(n_260)
);


endmodule