module fake_jpeg_172_n_550 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_550);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_550;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_441;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_47),
.B(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_25),
.B(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_51),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_54),
.B(n_89),
.Y(n_141)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_56),
.Y(n_145)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g163 ( 
.A(n_57),
.Y(n_163)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_60),
.Y(n_154)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_26),
.A2(n_44),
.B(n_46),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_88),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_18),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_86),
.Y(n_104)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_14),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_15),
.B(n_0),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_22),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_96),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_15),
.B(n_20),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_94),
.B(n_95),
.Y(n_156)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

BUFx12f_ASAP7_75t_SL g96 ( 
.A(n_18),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_97),
.Y(n_153)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_99),
.Y(n_159)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_30),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_101),
.B(n_102),
.Y(n_147)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_39),
.B1(n_44),
.B2(n_28),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_109),
.A2(n_137),
.B1(n_166),
.B2(n_87),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_110),
.B(n_123),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_20),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_115),
.B(n_116),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_42),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_42),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_19),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_125),
.B(n_136),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_69),
.B(n_27),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_51),
.A2(n_44),
.B1(n_28),
.B2(n_14),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_27),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_138),
.B(n_142),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_93),
.A2(n_98),
.B1(n_55),
.B2(n_77),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_151),
.B1(n_153),
.B2(n_35),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_56),
.B(n_45),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_45),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_150),
.B(n_157),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_49),
.A2(n_14),
.B1(n_46),
.B2(n_22),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_64),
.B(n_23),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_59),
.B(n_23),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g207 ( 
.A1(n_160),
.A2(n_52),
.B(n_18),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_63),
.B(n_34),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_164),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_61),
.A2(n_44),
.B1(n_28),
.B2(n_34),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_106),
.A2(n_101),
.B1(n_97),
.B2(n_66),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_169),
.A2(n_176),
.B1(n_147),
.B2(n_144),
.Y(n_227)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_34),
.B1(n_35),
.B2(n_30),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_171),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_74),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_172),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_180),
.Y(n_221)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_175),
.Y(n_226)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_38),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_201),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_114),
.B(n_65),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_179),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_114),
.B(n_72),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_103),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_182),
.A2(n_184),
.B1(n_208),
.B2(n_209),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_121),
.Y(n_183)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_107),
.A2(n_35),
.B1(n_84),
.B2(n_82),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_186),
.A2(n_199),
.B1(n_205),
.B2(n_206),
.Y(n_224)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_190),
.B(n_191),
.Y(n_240)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_200),
.Y(n_245)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

BUFx8_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_196),
.Y(n_231)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

CKINVDCx12_ASAP7_75t_R g252 ( 
.A(n_197),
.Y(n_252)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_198),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_151),
.A2(n_80),
.B1(n_78),
.B2(n_73),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_46),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_203),
.Y(n_247)
);

BUFx4f_ASAP7_75t_SL g203 ( 
.A(n_105),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_207),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_137),
.A2(n_40),
.B(n_22),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_131),
.A2(n_70),
.B1(n_68),
.B2(n_18),
.Y(n_206)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

INVx3_ASAP7_75t_SL g209 ( 
.A(n_163),
.Y(n_209)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_108),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_213),
.A2(n_216),
.B1(n_145),
.B2(n_134),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_105),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_215),
.Y(n_236)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_120),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_144),
.B1(n_152),
.B2(n_162),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_217),
.A2(n_228),
.B1(n_237),
.B2(n_209),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_119),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_179),
.C(n_172),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_227),
.A2(n_230),
.B1(n_234),
.B2(n_235),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_162),
.B1(n_152),
.B2(n_155),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_176),
.A2(n_164),
.B1(n_166),
.B2(n_122),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_L g234 ( 
.A1(n_173),
.A2(n_163),
.B1(n_131),
.B2(n_139),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_180),
.A2(n_122),
.B1(n_139),
.B2(n_132),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_132),
.B1(n_155),
.B2(n_167),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_178),
.B(n_129),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_251),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_180),
.A2(n_135),
.B1(n_124),
.B2(n_127),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_184),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_246),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_179),
.A2(n_145),
.B1(n_128),
.B2(n_118),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_172),
.B(n_118),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_256),
.B(n_259),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_257),
.A2(n_261),
.B1(n_271),
.B2(n_275),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_177),
.B(n_181),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_258),
.A2(n_270),
.B(n_249),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_168),
.C(n_174),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_223),
.B(n_194),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_260),
.B(n_269),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_254),
.A2(n_171),
.B1(n_182),
.B2(n_127),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_210),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_263),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_200),
.C(n_188),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_264),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_267),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_187),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_277),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_183),
.Y(n_269)
);

NAND2xp67_ASAP7_75t_L g270 ( 
.A(n_221),
.B(n_112),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_224),
.A2(n_227),
.B1(n_222),
.B2(n_244),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_135),
.B1(n_167),
.B2(n_124),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_273),
.B1(n_228),
.B2(n_220),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_183),
.B1(n_185),
.B2(n_170),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_224),
.A2(n_211),
.B1(n_213),
.B2(n_215),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_203),
.C(n_208),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_203),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_217),
.A2(n_192),
.B1(n_154),
.B2(n_202),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_242),
.A2(n_237),
.B1(n_238),
.B2(n_230),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_253),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_239),
.Y(n_279)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_229),
.Y(n_280)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_233),
.Y(n_281)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_243),
.B(n_193),
.CI(n_133),
.CON(n_284),
.SN(n_284)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_284),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_226),
.Y(n_285)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_293),
.A2(n_314),
.B(n_279),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_266),
.B(n_236),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_297),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_295),
.A2(n_303),
.B1(n_311),
.B2(n_257),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_236),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_240),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_302),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_310),
.C(n_239),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_233),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_282),
.A2(n_257),
.B1(n_265),
.B2(n_271),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_307),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_308),
.Y(n_331)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_309),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_259),
.B(n_231),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_282),
.A2(n_246),
.B1(n_220),
.B2(n_241),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_283),
.A2(n_247),
.B(n_241),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_269),
.Y(n_315)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_269),
.Y(n_316)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_276),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_259),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_255),
.B(n_258),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_318),
.A2(n_329),
.B(n_339),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_289),
.B(n_260),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_343),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_320),
.A2(n_292),
.B(n_298),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_299),
.A2(n_257),
.B1(n_278),
.B2(n_269),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_322),
.A2(n_332),
.B1(n_348),
.B2(n_316),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_326),
.A2(n_330),
.B1(n_334),
.B2(n_338),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_256),
.C(n_263),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_335),
.C(n_336),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_SL g329 ( 
.A(n_312),
.B(n_262),
.C(n_256),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_303),
.A2(n_275),
.B1(n_261),
.B2(n_264),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_299),
.A2(n_272),
.B1(n_284),
.B2(n_270),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_313),
.B(n_308),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_346),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_247),
.C(n_231),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_310),
.B(n_270),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_232),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_306),
.C(n_304),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_314),
.A2(n_279),
.B(n_239),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_305),
.A2(n_284),
.B1(n_285),
.B2(n_239),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_340),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_295),
.A2(n_284),
.B(n_239),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_341),
.A2(n_292),
.B(n_252),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_296),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_342),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_296),
.B(n_225),
.Y(n_343)
);

NAND3xp33_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_252),
.C(n_248),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_344),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_290),
.B(n_232),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_299),
.A2(n_305),
.B1(n_287),
.B2(n_291),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_290),
.B(n_225),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_349),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_297),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_351),
.B(n_362),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_326),
.A2(n_287),
.B1(n_291),
.B2(n_286),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_354),
.A2(n_359),
.B1(n_361),
.B2(n_383),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_323),
.Y(n_355)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_355),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_348),
.A2(n_311),
.B1(n_315),
.B2(n_286),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_294),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_309),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_381),
.C(n_356),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_320),
.A2(n_301),
.B(n_293),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_365),
.A2(n_376),
.B(n_373),
.Y(n_391)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_321),
.Y(n_366)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_332),
.A2(n_300),
.B1(n_302),
.B2(n_288),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_367),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_322),
.A2(n_307),
.B1(n_293),
.B2(n_304),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_368),
.A2(n_373),
.B(n_377),
.Y(n_398)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_323),
.Y(n_371)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_381),
.Y(n_414)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_345),
.Y(n_374)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_324),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_328),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_318),
.A2(n_292),
.B(n_298),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_339),
.A2(n_342),
.B(n_347),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_379),
.A2(n_382),
.B(n_341),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_324),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_380),
.B(n_357),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_337),
.B(n_277),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_347),
.A2(n_285),
.B(n_248),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_330),
.A2(n_226),
.B1(n_248),
.B2(n_225),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_331),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_384),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_356),
.B(n_331),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_396),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_345),
.Y(n_386)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_386),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_388),
.B(n_408),
.Y(n_434)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_389),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_374),
.Y(n_390)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_390),
.Y(n_420)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_370),
.B(n_336),
.C(n_346),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_412),
.C(n_353),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_352),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_395),
.A2(n_406),
.B1(n_411),
.B2(n_369),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_362),
.B(n_328),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_218),
.Y(n_397)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_397),
.Y(n_427)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_399),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_325),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_401),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_404),
.B(n_410),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_351),
.B(n_218),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_405),
.B(n_407),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_379),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_360),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_355),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_360),
.B(n_226),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_366),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_370),
.B(n_329),
.C(n_350),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_197),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_415),
.B(n_436),
.Y(n_442)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_417),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_393),
.A2(n_378),
.B1(n_367),
.B2(n_359),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_419),
.A2(n_429),
.B1(n_437),
.B2(n_441),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_392),
.B(n_353),
.C(n_377),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_422),
.C(n_428),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_388),
.B(n_414),
.C(n_402),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_363),
.C(n_376),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_393),
.A2(n_378),
.B1(n_350),
.B2(n_361),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_413),
.A2(n_368),
.B1(n_365),
.B2(n_354),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_430),
.A2(n_432),
.B1(n_411),
.B2(n_409),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_406),
.A2(n_371),
.B1(n_325),
.B2(n_382),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_383),
.C(n_175),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_390),
.C(n_404),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_398),
.A2(n_190),
.B1(n_198),
.B2(n_216),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_385),
.B(n_204),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_439),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_SL g439 ( 
.A(n_391),
.B(n_133),
.C(n_161),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_389),
.A2(n_40),
.B1(n_128),
.B2(n_112),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_424),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_444),
.B(n_2),
.Y(n_476)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_420),
.Y(n_445)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_445),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_446),
.B(n_219),
.C(n_18),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_398),
.C(n_396),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_448),
.B(n_450),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_434),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_423),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_387),
.C(n_403),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_416),
.A2(n_408),
.B1(n_401),
.B2(n_387),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_453),
.A2(n_219),
.B1(n_161),
.B2(n_133),
.Y(n_477)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_426),
.Y(n_454)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_454),
.Y(n_469)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_431),
.Y(n_455)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_403),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_457),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_421),
.B(n_390),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_416),
.Y(n_458)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_458),
.Y(n_475)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_459),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_440),
.A2(n_409),
.B(n_400),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_460),
.A2(n_461),
.B(n_464),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_440),
.A2(n_435),
.B(n_430),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_462),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_400),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_463),
.B(n_2),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_437),
.A2(n_420),
.B(n_418),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_459),
.A2(n_425),
.B1(n_427),
.B2(n_394),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_466),
.A2(n_468),
.B1(n_472),
.B2(n_474),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_447),
.A2(n_394),
.B1(n_439),
.B2(n_438),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_461),
.A2(n_415),
.B1(n_433),
.B2(n_423),
.Y(n_472)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_473),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_451),
.A2(n_40),
.B1(n_130),
.B2(n_161),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_477),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_482),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_219),
.C(n_18),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_483),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_456),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_443),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_484),
.B(n_448),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_443),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_487),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_446),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_488),
.B(n_502),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_470),
.A2(n_445),
.B1(n_460),
.B2(n_453),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_489),
.A2(n_493),
.B1(n_496),
.B2(n_467),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_470),
.A2(n_452),
.B1(n_463),
.B2(n_442),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_466),
.B(n_442),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_499),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_485),
.A2(n_452),
.B1(n_52),
.B2(n_33),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_485),
.A2(n_33),
.B(n_3),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_497),
.A2(n_501),
.B(n_469),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_475),
.B(n_2),
.Y(n_498)
);

NOR3xp33_ASAP7_75t_SL g517 ( 
.A(n_498),
.B(n_5),
.C(n_6),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_472),
.B(n_473),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_471),
.B(n_3),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_500),
.B(n_4),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_467),
.A2(n_33),
.B(n_5),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_4),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_486),
.A2(n_480),
.B(n_475),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_504),
.A2(n_510),
.B(n_491),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_505),
.B(n_515),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_481),
.C(n_478),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_508),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_512),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_492),
.A2(n_471),
.B(n_469),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_499),
.B(n_468),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_498),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_516),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_495),
.B(n_477),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_490),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_517),
.B(n_518),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_6),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_502),
.Y(n_520)
);

AOI21xp33_ASAP7_75t_L g535 ( 
.A1(n_520),
.A2(n_523),
.B(n_8),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_494),
.C(n_491),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_524),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_494),
.C(n_7),
.Y(n_524)
);

NOR2x1_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_6),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_526),
.A2(n_517),
.B(n_518),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_6),
.Y(n_529)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_529),
.Y(n_537)
);

AO21x1_ASAP7_75t_L g540 ( 
.A1(n_530),
.A2(n_528),
.B(n_526),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_507),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_531),
.A2(n_532),
.B(n_535),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_519),
.B(n_7),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_522),
.B(n_8),
.C(n_9),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_534),
.B(n_11),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_8),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_536),
.A2(n_9),
.B(n_10),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_533),
.B(n_520),
.C(n_525),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_538),
.A2(n_540),
.B(n_11),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_541),
.B(n_542),
.C(n_537),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_543),
.B(n_544),
.C(n_545),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_539),
.A2(n_11),
.B(n_12),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_12),
.Y(n_547)
);

AO21x1_ASAP7_75t_L g548 ( 
.A1(n_547),
.A2(n_12),
.B(n_13),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_SL g549 ( 
.A(n_548),
.B(n_12),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_12),
.B(n_13),
.Y(n_550)
);


endmodule