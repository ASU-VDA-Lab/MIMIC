module fake_jpeg_13317_n_309 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_10),
.B(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_48),
.B(n_63),
.Y(n_143)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_74),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_13),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_68),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_71),
.B(n_80),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_76),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_86),
.Y(n_100)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_78),
.B(n_84),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_31),
.B(n_1),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_26),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_82),
.A2(n_6),
.B1(n_8),
.B2(n_12),
.Y(n_133)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_31),
.B(n_2),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_42),
.B(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_88),
.Y(n_108)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_90),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_42),
.B(n_3),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_35),
.B(n_24),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_94),
.Y(n_131)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_24),
.B1(n_41),
.B2(n_36),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_44),
.B1(n_25),
.B2(n_29),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_95),
.A2(n_101),
.B1(n_107),
.B2(n_137),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_44),
.B1(n_25),
.B2(n_29),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_23),
.B1(n_41),
.B2(n_36),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_19),
.C(n_23),
.Y(n_116)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_116),
.B(n_117),
.CI(n_139),
.CON(n_178),
.SN(n_178)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_33),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_124),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_33),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_134),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_43),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_43),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_128),
.B(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_55),
.B(n_6),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_101),
.B1(n_144),
.B2(n_95),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_61),
.B(n_6),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_59),
.A2(n_73),
.B1(n_68),
.B2(n_58),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_52),
.B(n_75),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_74),
.Y(n_148)
);

AO22x1_ASAP7_75t_SL g142 ( 
.A1(n_65),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_140),
.B1(n_137),
.B2(n_58),
.Y(n_182)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_57),
.B1(n_74),
.B2(n_132),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_184),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_105),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_154),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_98),
.A2(n_57),
.B1(n_135),
.B2(n_115),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_151),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_152),
.B(n_168),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_118),
.B1(n_144),
.B2(n_127),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_153),
.A2(n_156),
.B1(n_169),
.B2(n_182),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_100),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_99),
.A2(n_141),
.B1(n_119),
.B2(n_135),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_122),
.B(n_140),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_162),
.C(n_184),
.Y(n_200)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

INVx6_ASAP7_75t_SL g159 ( 
.A(n_112),
.Y(n_159)
);

NAND2x1_ASAP7_75t_SL g208 ( 
.A(n_159),
.B(n_177),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_102),
.A2(n_107),
.B(n_97),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_166),
.B(n_162),
.Y(n_185)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_99),
.B(n_114),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_108),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_164),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_119),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_173),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_113),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_137),
.A2(n_103),
.B1(n_109),
.B2(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_109),
.Y(n_173)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_113),
.B(n_111),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_176),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_111),
.B(n_129),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_183),
.Y(n_193)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_130),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_120),
.B(n_121),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_185),
.A2(n_171),
.B(n_158),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_184),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_179),
.C(n_180),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_166),
.A2(n_160),
.B(n_169),
.C(n_172),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_207),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_205),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_206),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_167),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_208),
.Y(n_227)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_157),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

NAND2x1_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_178),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_223),
.B(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_178),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_222),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_152),
.B1(n_173),
.B2(n_165),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_199),
.B1(n_196),
.B2(n_186),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_189),
.B(n_165),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_185),
.A2(n_145),
.B(n_163),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_R g224 ( 
.A(n_195),
.B(n_161),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_224),
.B(n_229),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_164),
.B(n_170),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_205),
.B(n_146),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_228),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_155),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_188),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_232),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_208),
.B(n_206),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_181),
.C(n_174),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_221),
.A2(n_201),
.B(n_202),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_233),
.A2(n_235),
.B(n_246),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_198),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_226),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_247),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_191),
.B1(n_201),
.B2(n_210),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_250),
.B1(n_227),
.B2(n_231),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_199),
.B1(n_192),
.B2(n_203),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_249),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_215),
.A2(n_199),
.B1(n_187),
.B2(n_192),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_215),
.A2(n_197),
.B1(n_186),
.B2(n_204),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_253),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_228),
.B1(n_212),
.B2(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_214),
.C(n_232),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_265),
.C(n_245),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_214),
.B1(n_227),
.B2(n_230),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_264),
.B1(n_250),
.B2(n_237),
.Y(n_272)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_222),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_260),
.B(n_261),
.Y(n_268)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_220),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_263),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_236),
.B(n_235),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_225),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_274),
.C(n_275),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_237),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_272),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_236),
.C(n_235),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_233),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_249),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_252),
.Y(n_279)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_251),
.Y(n_286)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_256),
.B1(n_262),
.B2(n_259),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_274),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_282),
.A2(n_283),
.B1(n_259),
.B2(n_256),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_248),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_287),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_267),
.C(n_276),
.Y(n_287)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_290),
.Y(n_293)
);

OAI221xp5_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_251),
.B1(n_289),
.B2(n_288),
.C(n_291),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_285),
.C(n_284),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_296),
.C(n_238),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_284),
.C(n_281),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_264),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_280),
.B1(n_277),
.B2(n_244),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_299),
.C(n_300),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_264),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_301),
.A2(n_264),
.B(n_218),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_303),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_301),
.A2(n_234),
.B(n_218),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_211),
.B(n_234),
.C(n_216),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_302),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_306),
.Y(n_309)
);


endmodule