module fake_jpeg_18321_n_39 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_39);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

AOI21xp33_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_9),
.B(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_20),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_16),
.B(n_18),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_4),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_13),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_5),
.C(n_10),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_11),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_28),
.Y(n_39)
);


endmodule