module real_jpeg_31832_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_23),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_2),
.B(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_4),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_5),
.B(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_6),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_7),
.B(n_67),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_69),
.Y(n_10)
);

OA21x2_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_48),
.B(n_68),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_26),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_14),
.B(n_26),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_21),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_15),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_15),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_39),
.B2(n_40),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_29),
.B(n_35),
.C(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_41),
.B(n_43),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_61),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_60),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_60),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_97),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_72),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_86),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

BUFx4f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_94),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);


endmodule