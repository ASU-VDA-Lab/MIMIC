module fake_aes_8521_n_32 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx3_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
AND3x2_ASAP7_75t_L g16 ( .A(n_2), .B(n_6), .C(n_1), .Y(n_16) );
O2A1O1Ixp5_ASAP7_75t_SL g17 ( .A1(n_11), .A2(n_0), .B(n_2), .C(n_3), .Y(n_17) );
AOI21x1_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_0), .B(n_3), .Y(n_18) );
OAI221xp5_ASAP7_75t_L g19 ( .A1(n_11), .A2(n_0), .B1(n_4), .B2(n_5), .C(n_6), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_12), .B(n_4), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_11), .B(n_10), .Y(n_21) );
NAND2xp5_ASAP7_75t_SL g22 ( .A(n_20), .B(n_11), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_21), .Y(n_23) );
BUFx3_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_22), .B(n_13), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_24), .Y(n_26) );
NAND3xp33_ASAP7_75t_L g27 ( .A(n_26), .B(n_17), .C(n_23), .Y(n_27) );
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_27), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_27), .Y(n_29) );
AOI22xp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_15), .B1(n_14), .B2(n_16), .Y(n_30) );
OAI21xp33_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_18), .B(n_16), .Y(n_31) );
AOI22xp33_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_8), .B1(n_9), .B2(n_30), .Y(n_32) );
endmodule