module fake_jpeg_17183_n_249 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_37),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_46),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_25),
.B1(n_26),
.B2(n_17),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_17),
.Y(n_46)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_19),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_26),
.B1(n_25),
.B2(n_18),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_32),
.B1(n_23),
.B2(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_32),
.B1(n_27),
.B2(n_21),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_57),
.B(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_77),
.B1(n_82),
.B2(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_30),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_27),
.B(n_18),
.C(n_21),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_30),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_17),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_20),
.B1(n_31),
.B2(n_45),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_35),
.B1(n_24),
.B2(n_23),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_45),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_19),
.B1(n_23),
.B2(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_80),
.Y(n_97)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_52),
.B(n_27),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_84),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_0),
.B(n_1),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_32),
.B1(n_54),
.B2(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_24),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_54),
.B(n_21),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_45),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_95),
.B1(n_103),
.B2(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_88),
.B(n_75),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_99),
.B1(n_105),
.B2(n_81),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_79),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_72),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_31),
.B1(n_22),
.B2(n_20),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_71),
.B1(n_64),
.B2(n_76),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_31),
.B1(n_22),
.B2(n_20),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_10),
.B1(n_15),
.B2(n_13),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_20),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_107),
.B(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_31),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

AOI22x1_ASAP7_75t_L g112 ( 
.A1(n_59),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_82),
.B(n_69),
.C(n_63),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_113),
.A2(n_127),
.B(n_95),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_116),
.B1(n_131),
.B2(n_138),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_59),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_125),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_86),
.Y(n_119)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_65),
.B(n_83),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_130),
.B(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_68),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_126),
.Y(n_154)
);

AOI31xp33_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_68),
.A3(n_80),
.B(n_71),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_87),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_67),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_0),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_109),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NOR2x1_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_0),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_1),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_134),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_97),
.B(n_107),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_89),
.A2(n_64),
.B(n_76),
.C(n_66),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_138)
);

NOR4xp25_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_98),
.C(n_93),
.D(n_95),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_146),
.C(n_163),
.Y(n_166)
);

AOI221xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_116),
.B1(n_130),
.B2(n_113),
.C(n_120),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_148),
.C(n_150),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_129),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_102),
.C(n_103),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_99),
.B1(n_104),
.B2(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_93),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_93),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_155),
.C(n_159),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_125),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_130),
.B(n_126),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_110),
.B1(n_104),
.B2(n_94),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_158),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_108),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_108),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_162),
.C(n_156),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_3),
.C(n_5),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_129),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_152),
.B(n_139),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_113),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_173),
.C(n_178),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_114),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_132),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_183),
.Y(n_194)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_179),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_180),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_120),
.A3(n_127),
.B1(n_115),
.B2(n_137),
.C1(n_138),
.C2(n_131),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_142),
.B1(n_139),
.B2(n_147),
.Y(n_187)
);

OAI322xp33_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_127),
.A3(n_137),
.B1(n_7),
.B2(n_8),
.C1(n_10),
.C2(n_3),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_162),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_185),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_140),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_170),
.B(n_174),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_166),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_152),
.B1(n_161),
.B2(n_149),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_200),
.B1(n_185),
.B2(n_182),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_148),
.B1(n_143),
.B2(n_153),
.Y(n_193)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_145),
.C(n_150),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_198),
.C(n_168),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_197),
.B(n_172),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_6),
.C(n_8),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_176),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_201),
.B(n_179),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_202),
.A2(n_204),
.B1(n_209),
.B2(n_213),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_212),
.C(n_196),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_210),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_173),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_207),
.A2(n_190),
.B1(n_193),
.B2(n_187),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_212),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_190),
.A2(n_175),
.B(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_211),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_168),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_178),
.B1(n_175),
.B2(n_171),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_203),
.B(n_197),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_221),
.C(n_216),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_202),
.C(n_210),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_213),
.C(n_207),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_195),
.B(n_194),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_191),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_186),
.B1(n_195),
.B2(n_200),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

AOI21x1_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_215),
.B(n_217),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_231),
.C(n_221),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_220),
.B(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_219),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_223),
.A2(n_191),
.B(n_199),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_230),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_222),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_235),
.C(n_236),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_SL g240 ( 
.A(n_237),
.B(n_231),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_238),
.A2(n_215),
.B1(n_225),
.B2(n_199),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_239),
.B(n_180),
.Y(n_243)
);

AOI21x1_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_11),
.B(n_12),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_184),
.C(n_181),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_245),
.C(n_242),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_12),
.C(n_13),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_247),
.Y(n_249)
);


endmodule