module fake_aes_7433_n_702 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_702);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_702;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_649;
wire n_276;
wire n_526;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_15), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_44), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_4), .Y(n_82) );
INVx1_ASAP7_75t_SL g83 ( .A(n_51), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_45), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_78), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_49), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_50), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_31), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_6), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_40), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_73), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_24), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_20), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_58), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_7), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_69), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_38), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_65), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_12), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_64), .Y(n_100) );
CKINVDCx14_ASAP7_75t_R g101 ( .A(n_75), .Y(n_101) );
BUFx2_ASAP7_75t_L g102 ( .A(n_42), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_33), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_41), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_14), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_0), .Y(n_106) );
INVxp33_ASAP7_75t_SL g107 ( .A(n_6), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_32), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_29), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_18), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_68), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_66), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_16), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_30), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_55), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_59), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_3), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_7), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_19), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_72), .Y(n_122) );
NOR2xp67_ASAP7_75t_L g123 ( .A(n_56), .B(n_47), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_11), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_23), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_62), .Y(n_126) );
CKINVDCx16_ASAP7_75t_R g127 ( .A(n_11), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_3), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_93), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_88), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_102), .B(n_1), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_88), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_102), .B(n_1), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_112), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_90), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_90), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_98), .B(n_2), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_114), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_112), .Y(n_139) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_91), .A2(n_35), .B(n_77), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_91), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_80), .B(n_2), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_116), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_116), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_92), .B(n_34), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_80), .B(n_4), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_92), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_89), .B(n_5), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_96), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_127), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_114), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_87), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_96), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_103), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_97), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_85), .Y(n_156) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_97), .A2(n_36), .B(n_76), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_85), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_89), .B(n_5), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_95), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_95), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_124), .B(n_8), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_101), .B(n_8), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_108), .B(n_9), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_104), .B(n_9), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_104), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_100), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_110), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_117), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_121), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_122), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_125), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_156), .B(n_81), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_138), .B(n_126), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_131), .B(n_128), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_131), .B(n_128), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_138), .B(n_126), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_158), .B(n_84), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_131), .B(n_124), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_134), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_132), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_168), .B(n_125), .Y(n_183) );
INVx6_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_134), .Y(n_186) );
BUFx4f_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVxp67_ASAP7_75t_L g188 ( .A(n_172), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_160), .B(n_82), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_168), .B(n_107), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_169), .B(n_107), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_132), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_145), .Y(n_193) );
INVx4_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_145), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_145), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_142), .Y(n_197) );
NAND3xp33_ASAP7_75t_L g198 ( .A(n_133), .B(n_137), .C(n_161), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_142), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_142), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_140), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_132), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_134), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_143), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_143), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_139), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_139), .Y(n_209) );
AND2x6_ASAP7_75t_L g210 ( .A(n_148), .B(n_99), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_169), .B(n_94), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_160), .B(n_111), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_137), .A2(n_106), .B1(n_120), .B2(n_119), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_139), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_144), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_148), .Y(n_216) );
INVx4_ASAP7_75t_SL g217 ( .A(n_145), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_148), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_144), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_148), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_170), .B(n_86), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_144), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_167), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_130), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_161), .B(n_118), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_130), .Y(n_226) );
OR2x6_ASAP7_75t_L g227 ( .A(n_133), .B(n_123), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_135), .B(n_115), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_135), .B(n_113), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_136), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_137), .B(n_105), .Y(n_231) );
OAI221xp5_ASAP7_75t_L g232 ( .A1(n_146), .A2(n_109), .B1(n_83), .B2(n_13), .C(n_14), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_136), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_167), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_141), .B(n_10), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_170), .B(n_10), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_141), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_147), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_235), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_210), .Y(n_240) );
INVxp67_ASAP7_75t_L g241 ( .A(n_174), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_235), .Y(n_242) );
NAND2x1p5_ASAP7_75t_L g243 ( .A(n_235), .B(n_164), .Y(n_243) );
AND2x2_ASAP7_75t_SL g244 ( .A(n_187), .B(n_164), .Y(n_244) );
NOR3xp33_ASAP7_75t_SL g245 ( .A(n_232), .B(n_129), .C(n_154), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_228), .B(n_164), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_193), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_181), .Y(n_248) );
INVx5_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_181), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_193), .Y(n_251) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_179), .B(n_163), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_231), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_194), .B(n_163), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_194), .B(n_153), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_188), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_194), .B(n_153), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_182), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_228), .B(n_149), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_182), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_231), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_177), .Y(n_262) );
NOR2xp67_ASAP7_75t_L g263 ( .A(n_213), .B(n_171), .Y(n_263) );
AND2x6_ASAP7_75t_L g264 ( .A(n_216), .B(n_147), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_227), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_195), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_192), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_227), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_228), .B(n_155), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_195), .B(n_155), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_192), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_229), .B(n_149), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_210), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_229), .B(n_166), .Y(n_274) );
INVx8_ASAP7_75t_L g275 ( .A(n_210), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_229), .B(n_166), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_210), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_179), .Y(n_278) );
INVx3_ASAP7_75t_L g279 ( .A(n_184), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_227), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_210), .Y(n_281) );
NOR2xp33_ASAP7_75t_R g282 ( .A(n_187), .B(n_151), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_198), .B(n_190), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_179), .Y(n_284) );
AO22x1_ASAP7_75t_L g285 ( .A1(n_216), .A2(n_145), .B1(n_152), .B2(n_159), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_175), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_203), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_195), .B(n_171), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_203), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_175), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_183), .B(n_167), .Y(n_291) );
NAND2xp33_ASAP7_75t_SL g292 ( .A(n_196), .B(n_150), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_184), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_176), .B(n_162), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_204), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_196), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_223), .Y(n_297) );
BUFx6f_ASAP7_75t_SL g298 ( .A(n_227), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_184), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_176), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_189), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_197), .A2(n_162), .B(n_159), .C(n_146), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_196), .B(n_157), .Y(n_303) );
BUFx2_ASAP7_75t_R g304 ( .A(n_191), .Y(n_304) );
NAND2xp33_ASAP7_75t_R g305 ( .A(n_189), .B(n_212), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_184), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_204), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_207), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_207), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_300), .B(n_212), .Y(n_310) );
INVxp67_ASAP7_75t_SL g311 ( .A(n_243), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_243), .B(n_225), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_283), .A2(n_220), .B1(n_218), .B2(n_225), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_252), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_278), .Y(n_315) );
INVx5_ASAP7_75t_L g316 ( .A(n_275), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_260), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_260), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_275), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_283), .A2(n_220), .B1(n_218), .B2(n_200), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_275), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_294), .B(n_211), .Y(n_322) );
OAI221xp5_ASAP7_75t_L g323 ( .A1(n_305), .A2(n_221), .B1(n_178), .B2(n_173), .C(n_236), .Y(n_323) );
INVx5_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_240), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_284), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_253), .B(n_237), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_256), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_252), .Y(n_329) );
BUFx8_ASAP7_75t_L g330 ( .A(n_298), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_261), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_241), .B(n_237), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_244), .A2(n_218), .B1(n_220), .B2(n_199), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_281), .B(n_187), .Y(n_334) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_303), .A2(n_233), .B(n_230), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_301), .B(n_233), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_305), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_240), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_292), .Y(n_339) );
NOR2x1_ASAP7_75t_SL g340 ( .A(n_249), .B(n_230), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_262), .B(n_238), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_246), .B(n_226), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_302), .B(n_226), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_286), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_266), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_249), .B(n_224), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_302), .A2(n_224), .B(n_234), .C(n_223), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_264), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_242), .A2(n_222), .B1(n_214), .B2(n_219), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_249), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_282), .Y(n_351) );
BUFx4f_ASAP7_75t_L g352 ( .A(n_264), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_267), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_239), .A2(n_222), .B1(n_214), .B2(n_219), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_264), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_282), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_267), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_266), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_290), .Y(n_359) );
BUFx3_ASAP7_75t_L g360 ( .A(n_249), .Y(n_360) );
BUFx10_ASAP7_75t_L g361 ( .A(n_264), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_271), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_304), .Y(n_363) );
INVx6_ASAP7_75t_L g364 ( .A(n_264), .Y(n_364) );
INVx5_ASAP7_75t_L g365 ( .A(n_364), .Y(n_365) );
INVx3_ASAP7_75t_SL g366 ( .A(n_364), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g367 ( .A1(n_347), .A2(n_255), .B(n_270), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_331), .Y(n_368) );
AO21x2_ASAP7_75t_L g369 ( .A1(n_335), .A2(n_303), .B(n_157), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_364), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_310), .A2(n_244), .B1(n_292), .B2(n_280), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_317), .Y(n_372) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_345), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_322), .B(n_263), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_317), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_318), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_318), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_337), .A2(n_298), .B1(n_268), .B2(n_265), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_312), .A2(n_239), .B1(n_254), .B2(n_299), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_359), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_352), .A2(n_269), .B1(n_274), .B2(n_272), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_364), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_345), .Y(n_383) );
INVx4_ASAP7_75t_L g384 ( .A(n_352), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_352), .A2(n_276), .B1(n_259), .B2(n_307), .Y(n_385) );
INVx3_ASAP7_75t_L g386 ( .A(n_361), .Y(n_386) );
AOI21xp33_ASAP7_75t_L g387 ( .A1(n_341), .A2(n_254), .B(n_277), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_343), .A2(n_270), .B(n_255), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_310), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_328), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_332), .A2(n_309), .B1(n_308), .B2(n_295), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_311), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_SL g393 ( .A1(n_347), .A2(n_291), .B(n_287), .C(n_250), .Y(n_393) );
AOI211xp5_ASAP7_75t_L g394 ( .A1(n_323), .A2(n_285), .B(n_165), .C(n_157), .Y(n_394) );
OAI22xp33_ASAP7_75t_L g395 ( .A1(n_328), .A2(n_273), .B1(n_271), .B2(n_258), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_312), .A2(n_245), .B1(n_299), .B2(n_306), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_353), .Y(n_397) );
INVx4_ASAP7_75t_L g398 ( .A(n_316), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_392), .B(n_336), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_389), .A2(n_339), .B1(n_344), .B2(n_314), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_391), .A2(n_339), .B1(n_336), .B2(n_327), .Y(n_401) );
NAND4xp25_ASAP7_75t_L g402 ( .A(n_374), .B(n_363), .C(n_327), .D(n_313), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_375), .B(n_353), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_392), .B(n_315), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_375), .B(n_329), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_368), .Y(n_406) );
OAI21x1_ASAP7_75t_L g407 ( .A1(n_367), .A2(n_348), .B(n_362), .Y(n_407) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_371), .A2(n_356), .B1(n_351), .B2(n_342), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_376), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_372), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_380), .A2(n_330), .B1(n_326), .B2(n_356), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g412 ( .A1(n_388), .A2(n_320), .B(n_333), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_395), .A2(n_330), .B1(n_145), .B2(n_306), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_393), .A2(n_362), .B(n_357), .Y(n_414) );
OAI21xp33_ASAP7_75t_L g415 ( .A1(n_394), .A2(n_357), .B(n_354), .Y(n_415) );
OAI21xp5_ASAP7_75t_L g416 ( .A1(n_376), .A2(n_349), .B(n_248), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_387), .A2(n_330), .B1(n_145), .B2(n_279), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_377), .Y(n_418) );
OAI21x1_ASAP7_75t_L g419 ( .A1(n_372), .A2(n_348), .B(n_346), .Y(n_419) );
OA21x2_ASAP7_75t_L g420 ( .A1(n_377), .A2(n_234), .B(n_289), .Y(n_420) );
INVx4_ASAP7_75t_SL g421 ( .A(n_366), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_396), .B(n_297), .Y(n_422) );
AOI222xp33_ASAP7_75t_L g423 ( .A1(n_390), .A2(n_348), .B1(n_355), .B2(n_334), .C1(n_186), .C2(n_205), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_397), .Y(n_424) );
INVx4_ASAP7_75t_L g425 ( .A(n_366), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_390), .A2(n_355), .B1(n_316), .B2(n_324), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_381), .A2(n_279), .B1(n_293), .B2(n_338), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_403), .B(n_397), .Y(n_428) );
AOI211xp5_ASAP7_75t_SL g429 ( .A1(n_401), .A2(n_385), .B(n_386), .C(n_180), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_409), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_409), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_402), .B(n_406), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_403), .B(n_369), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_399), .A2(n_378), .B1(n_366), .B2(n_379), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_399), .A2(n_384), .B1(n_398), .B2(n_370), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_405), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_405), .B(n_370), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_402), .B(n_208), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_420), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_400), .A2(n_384), .B1(n_398), .B2(n_365), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_425), .Y(n_441) );
NAND2xp33_ASAP7_75t_R g442 ( .A(n_420), .B(n_140), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_404), .Y(n_443) );
NAND4xp25_ASAP7_75t_SL g444 ( .A(n_411), .B(n_12), .C(n_13), .D(n_15), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_418), .B(n_369), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_418), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_408), .B(n_208), .Y(n_447) );
OR2x6_ASAP7_75t_L g448 ( .A(n_425), .B(n_384), .Y(n_448) );
INVxp67_ASAP7_75t_L g449 ( .A(n_410), .Y(n_449) );
OAI33xp33_ASAP7_75t_L g450 ( .A1(n_422), .A2(n_206), .A3(n_205), .B1(n_186), .B2(n_180), .B3(n_209), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_412), .A2(n_382), .B1(n_398), .B2(n_386), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_410), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_421), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_424), .B(n_383), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_425), .B(n_382), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_424), .Y(n_456) );
OAI21xp33_ASAP7_75t_L g457 ( .A1(n_413), .A2(n_206), .B(n_209), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_427), .A2(n_365), .B1(n_386), .B2(n_316), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_415), .A2(n_215), .B1(n_293), .B2(n_297), .C(n_185), .Y(n_459) );
OAI211xp5_ASAP7_75t_SL g460 ( .A1(n_423), .A2(n_215), .B(n_288), .C(n_257), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_420), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_420), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_416), .B(n_369), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_415), .A2(n_407), .B(n_414), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_436), .B(n_423), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_446), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_461), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_443), .B(n_416), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_461), .Y(n_469) );
NOR2x1p5_ASAP7_75t_L g470 ( .A(n_441), .B(n_421), .Y(n_470) );
INVx4_ASAP7_75t_L g471 ( .A(n_448), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_446), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_428), .B(n_407), .Y(n_473) );
AND2x2_ASAP7_75t_SL g474 ( .A(n_439), .B(n_421), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_428), .B(n_419), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_441), .B(n_421), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_462), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_438), .A2(n_417), .B(n_419), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_430), .B(n_426), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_462), .Y(n_480) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_454), .Y(n_481) );
INVxp33_ASAP7_75t_L g482 ( .A(n_432), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_439), .B(n_16), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_452), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_431), .B(n_17), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_445), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_444), .A2(n_365), .B1(n_140), .B2(n_358), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_429), .A2(n_346), .B(n_334), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_454), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_453), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_445), .Y(n_491) );
AND2x4_ASAP7_75t_SL g492 ( .A(n_448), .B(n_373), .Y(n_492) );
AOI322xp5_ASAP7_75t_L g493 ( .A1(n_453), .A2(n_17), .A3(n_18), .B1(n_185), .B2(n_202), .C1(n_201), .C2(n_365), .Y(n_493) );
NAND4xp25_ASAP7_75t_SL g494 ( .A(n_437), .B(n_361), .C(n_365), .D(n_316), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_433), .B(n_383), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_433), .B(n_383), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_452), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_456), .Y(n_498) );
INVx3_ASAP7_75t_L g499 ( .A(n_448), .Y(n_499) );
BUFx2_ASAP7_75t_SL g500 ( .A(n_440), .Y(n_500) );
INVx1_ASAP7_75t_SL g501 ( .A(n_437), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_463), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_449), .B(n_383), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_463), .B(n_383), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_464), .B(n_373), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_451), .B(n_185), .C(n_202), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_434), .B(n_373), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_448), .B(n_373), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_455), .B(n_373), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_447), .Y(n_510) );
BUFx2_ASAP7_75t_L g511 ( .A(n_435), .Y(n_511) );
AOI33xp33_ASAP7_75t_L g512 ( .A1(n_459), .A2(n_319), .A3(n_321), .B1(n_25), .B2(n_26), .B3(n_27), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_442), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_458), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_450), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_457), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_490), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_501), .B(n_202), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_502), .B(n_202), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_467), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_486), .B(n_202), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_467), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_469), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_472), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_502), .B(n_201), .Y(n_526) );
NAND2xp33_ASAP7_75t_SL g527 ( .A(n_470), .B(n_325), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_491), .B(n_21), .Y(n_528) );
NOR2x1_ASAP7_75t_L g529 ( .A(n_470), .B(n_460), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_483), .B(n_22), .Y(n_530) );
NAND2x1p5_ASAP7_75t_L g531 ( .A(n_476), .B(n_316), .Y(n_531) );
BUFx2_ASAP7_75t_SL g532 ( .A(n_471), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_468), .B(n_201), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_465), .B(n_201), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_502), .B(n_185), .Y(n_535) );
NOR2xp33_ASAP7_75t_SL g536 ( .A(n_471), .B(n_361), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_491), .B(n_185), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_491), .B(n_28), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_497), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_485), .B(n_338), .C(n_319), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_482), .B(n_37), .Y(n_541) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_478), .A2(n_288), .B(n_257), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_474), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_498), .B(n_340), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_473), .B(n_39), .Y(n_545) );
INVxp67_ASAP7_75t_L g546 ( .A(n_483), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_473), .B(n_43), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_484), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_489), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_474), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_489), .B(n_46), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_475), .B(n_48), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_469), .Y(n_553) );
NOR3xp33_ASAP7_75t_L g554 ( .A(n_512), .B(n_338), .C(n_321), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_489), .B(n_52), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_480), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_475), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_496), .B(n_53), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_489), .B(n_345), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_496), .B(n_54), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_511), .B(n_345), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_511), .B(n_358), .Y(n_563) );
INVx5_ASAP7_75t_L g564 ( .A(n_471), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_474), .B(n_324), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_477), .B(n_481), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_510), .B(n_358), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_477), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_481), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_471), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_504), .B(n_57), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_527), .Y(n_572) );
AOI221x1_ASAP7_75t_L g573 ( .A1(n_527), .A2(n_499), .B1(n_515), .B2(n_488), .C(n_500), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_558), .B(n_504), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_529), .A2(n_500), .B1(n_499), .B2(n_510), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_546), .B(n_481), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_545), .B(n_495), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_541), .A2(n_499), .B1(n_509), .B2(n_514), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_566), .B(n_481), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_543), .B(n_499), .Y(n_580) );
NAND4xp25_ASAP7_75t_L g581 ( .A(n_541), .B(n_493), .C(n_487), .D(n_479), .Y(n_581) );
OAI21xp33_ASAP7_75t_L g582 ( .A1(n_562), .A2(n_493), .B(n_507), .Y(n_582) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_520), .Y(n_583) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_543), .A2(n_506), .B1(n_515), .B2(n_514), .Y(n_584) );
AO21x1_ASAP7_75t_L g585 ( .A1(n_565), .A2(n_492), .B(n_508), .Y(n_585) );
OAI221xp5_ASAP7_75t_SL g586 ( .A1(n_550), .A2(n_513), .B1(n_509), .B2(n_515), .C(n_516), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_524), .B(n_481), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_540), .A2(n_495), .B1(n_513), .B2(n_508), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_525), .B(n_495), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_539), .B(n_495), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_570), .A2(n_508), .B1(n_494), .B2(n_516), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_556), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g593 ( .A1(n_570), .A2(n_492), .B(n_508), .C(n_506), .Y(n_593) );
INVxp67_ASAP7_75t_SL g594 ( .A(n_520), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_517), .A2(n_505), .B1(n_492), .B2(n_503), .C(n_358), .Y(n_595) );
AOI22xp33_ASAP7_75t_SL g596 ( .A1(n_532), .A2(n_505), .B1(n_503), .B2(n_324), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_557), .B(n_60), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_549), .B(n_61), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_548), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_522), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_522), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_564), .A2(n_324), .B1(n_325), .B2(n_350), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_523), .Y(n_603) );
AOI21xp33_ASAP7_75t_L g604 ( .A1(n_530), .A2(n_63), .B(n_67), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_559), .Y(n_605) );
OAI311xp33_ASAP7_75t_L g606 ( .A1(n_555), .A2(n_70), .A3(n_74), .B1(n_79), .C1(n_217), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_523), .B(n_325), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_565), .A2(n_324), .B(n_360), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_553), .Y(n_609) );
NOR4xp25_ASAP7_75t_L g610 ( .A(n_544), .B(n_217), .C(n_325), .D(n_360), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_553), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_534), .A2(n_350), .B1(n_266), .B2(n_296), .C(n_247), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_545), .B(n_217), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_568), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_547), .B(n_217), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_559), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_563), .B(n_247), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g618 ( .A1(n_531), .A2(n_247), .B1(n_251), .B2(n_266), .C(n_296), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_605), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_600), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_574), .B(n_547), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_582), .B(n_569), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_581), .B(n_552), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_581), .B(n_552), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_577), .B(n_552), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_592), .Y(n_626) );
AOI21xp33_ASAP7_75t_L g627 ( .A1(n_588), .A2(n_551), .B(n_571), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_606), .A2(n_531), .B(n_554), .C(n_571), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_599), .Y(n_629) );
INVxp67_ASAP7_75t_L g630 ( .A(n_576), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_601), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_603), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_589), .B(n_535), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_578), .B(n_564), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_590), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_616), .B(n_564), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_583), .Y(n_637) );
XNOR2xp5_ASAP7_75t_L g638 ( .A(n_591), .B(n_561), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_580), .B(n_564), .Y(n_639) );
OAI211xp5_ASAP7_75t_SL g640 ( .A1(n_575), .A2(n_560), .B(n_533), .C(n_518), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_579), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_609), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_594), .B(n_521), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_611), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_614), .Y(n_645) );
INVxp33_ASAP7_75t_SL g646 ( .A(n_572), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_585), .A2(n_561), .B1(n_564), .B2(n_528), .Y(n_647) );
NAND2x1_ASAP7_75t_L g648 ( .A(n_580), .B(n_528), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_572), .B(n_528), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_619), .B(n_595), .Y(n_650) );
AOI322xp5_ASAP7_75t_L g651 ( .A1(n_623), .A2(n_584), .A3(n_593), .B1(n_596), .B2(n_587), .C1(n_538), .C2(n_615), .Y(n_651) );
INVxp67_ASAP7_75t_SL g652 ( .A(n_637), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_644), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_623), .A2(n_624), .B1(n_638), .B2(n_646), .Y(n_654) );
NAND4xp75_ASAP7_75t_L g655 ( .A(n_624), .B(n_573), .C(n_608), .D(n_604), .Y(n_655) );
NOR4xp25_ASAP7_75t_L g656 ( .A(n_622), .B(n_586), .C(n_606), .D(n_598), .Y(n_656) );
OAI221xp5_ASAP7_75t_SL g657 ( .A1(n_628), .A2(n_610), .B1(n_613), .B2(n_612), .C(n_618), .Y(n_657) );
NAND2x1p5_ASAP7_75t_L g658 ( .A(n_648), .B(n_538), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_641), .B(n_617), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_646), .A2(n_536), .B1(n_597), .B2(n_542), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_649), .A2(n_610), .B(n_602), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_626), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_642), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_629), .Y(n_664) );
OAI211xp5_ASAP7_75t_SL g665 ( .A1(n_627), .A2(n_567), .B(n_607), .C(n_542), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_634), .B(n_542), .C(n_519), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_635), .Y(n_667) );
INVxp67_ASAP7_75t_SL g668 ( .A(n_620), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_634), .A2(n_526), .B1(n_537), .B2(n_247), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_645), .B(n_537), .Y(n_670) );
OAI221xp5_ASAP7_75t_SL g671 ( .A1(n_654), .A2(n_647), .B1(n_621), .B2(n_636), .C(n_625), .Y(n_671) );
AOI31xp33_ASAP7_75t_L g672 ( .A1(n_661), .A2(n_649), .A3(n_639), .B(n_630), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_652), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_663), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_663), .Y(n_675) );
NOR2x1p5_ASAP7_75t_L g676 ( .A(n_655), .B(n_633), .Y(n_676) );
OR3x1_ASAP7_75t_L g677 ( .A(n_665), .B(n_640), .C(n_643), .Y(n_677) );
INVx2_ASAP7_75t_SL g678 ( .A(n_653), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_665), .A2(n_631), .B1(n_632), .B2(n_251), .Y(n_679) );
NOR2xp33_ASAP7_75t_SL g680 ( .A(n_657), .B(n_251), .Y(n_680) );
INVx1_ASAP7_75t_SL g681 ( .A(n_650), .Y(n_681) );
XNOR2xp5_ASAP7_75t_L g682 ( .A(n_656), .B(n_296), .Y(n_682) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_668), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_660), .A2(n_667), .B1(n_659), .B2(n_666), .Y(n_684) );
O2A1O1Ixp5_ASAP7_75t_SL g685 ( .A1(n_662), .A2(n_664), .B(n_657), .C(n_670), .Y(n_685) );
AOI211x1_ASAP7_75t_L g686 ( .A1(n_651), .A2(n_661), .B(n_650), .C(n_666), .Y(n_686) );
OAI22xp5_ASAP7_75t_SL g687 ( .A1(n_658), .A2(n_654), .B1(n_646), .B2(n_624), .Y(n_687) );
XOR2x2_ASAP7_75t_L g688 ( .A(n_669), .B(n_654), .Y(n_688) );
OR2x2_ASAP7_75t_L g689 ( .A(n_681), .B(n_683), .Y(n_689) );
NOR2x2_ASAP7_75t_L g690 ( .A(n_686), .B(n_677), .Y(n_690) );
CKINVDCx5p33_ASAP7_75t_R g691 ( .A(n_688), .Y(n_691) );
INVx1_ASAP7_75t_SL g692 ( .A(n_673), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_687), .Y(n_693) );
OA22x2_ASAP7_75t_L g694 ( .A1(n_691), .A2(n_684), .B1(n_682), .B2(n_685), .Y(n_694) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_690), .B(n_680), .C(n_671), .D(n_679), .Y(n_695) );
AND3x4_ASAP7_75t_L g696 ( .A(n_693), .B(n_677), .C(n_676), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_694), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_696), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_698), .Y(n_699) );
NAND4xp75_ASAP7_75t_L g700 ( .A(n_697), .B(n_695), .C(n_674), .D(n_675), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_700), .A2(n_692), .B1(n_689), .B2(n_678), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_701), .A2(n_699), .B(n_672), .Y(n_702) );
endmodule