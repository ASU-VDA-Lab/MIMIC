module fake_jpeg_4983_n_208 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_35),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_21),
.Y(n_47)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_23),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_24),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_22),
.B1(n_14),
.B2(n_21),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_14),
.B(n_33),
.C(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_33),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_32),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_73),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_28),
.B1(n_52),
.B2(n_50),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_SL g111 ( 
.A(n_78),
.B(n_73),
.C(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_93),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_56),
.B(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_66),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_45),
.C(n_44),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_87),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_42),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_42),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_51),
.B1(n_48),
.B2(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_1),
.Y(n_108)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_102),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_109),
.Y(n_118)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_69),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_104),
.B(n_106),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_48),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_108),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_32),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_78),
.B1(n_75),
.B2(n_31),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_2),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_17),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_74),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_89),
.B1(n_88),
.B2(n_84),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_121),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_76),
.B1(n_82),
.B2(n_78),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_132),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_76),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_96),
.C(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_113),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_84),
.B1(n_86),
.B2(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_141),
.C(n_124),
.Y(n_155)
);

OR2x4_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_103),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_134),
.B(n_26),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_130),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_142),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_111),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_128),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_103),
.B(n_85),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_144),
.A2(n_119),
.B1(n_122),
.B2(n_118),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_153),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_140),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_19),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_157),
.C(n_163),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_128),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_158),
.B(n_146),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_123),
.C(n_131),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_19),
.Y(n_158)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_136),
.B1(n_147),
.B2(n_149),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_94),
.B1(n_19),
.B2(n_26),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_162),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_26),
.C(n_17),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_143),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_166),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_136),
.C(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_172),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_13),
.C(n_12),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_174),
.A2(n_162),
.B1(n_154),
.B2(n_150),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_161),
.B(n_159),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_177),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_184),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_171),
.A2(n_26),
.B1(n_17),
.B2(n_16),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_181),
.B1(n_4),
.B2(n_5),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_164),
.A2(n_2),
.B(n_3),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_2),
.B(n_3),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_187),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_182),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_6),
.Y(n_196)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_179),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_190),
.B(n_6),
.Y(n_197)
);

AOI21x1_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_174),
.B(n_170),
.Y(n_190)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_17),
.CI(n_16),
.CON(n_192),
.SN(n_192)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_7),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_181),
.B1(n_16),
.B2(n_7),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_5),
.B(n_6),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_197),
.B(n_198),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_188),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_202),
.B1(n_8),
.B2(n_9),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_197),
.C(n_8),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.C(n_9),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_207),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g207 ( 
.A(n_205),
.Y(n_207)
);


endmodule