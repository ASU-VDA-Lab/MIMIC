module real_jpeg_6788_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_1),
.A2(n_39),
.B1(n_61),
.B2(n_82),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_2),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_2),
.Y(n_131)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_2),
.Y(n_139)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_2),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_2),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_2),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_2),
.Y(n_261)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_2),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_3),
.A2(n_146),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_3),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_3),
.A2(n_194),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_3),
.A2(n_45),
.B1(n_194),
.B2(n_336),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_3),
.A2(n_194),
.B1(n_282),
.B2(n_368),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_5),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_5),
.A2(n_81),
.B1(n_177),
.B2(n_181),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_5),
.A2(n_81),
.B1(n_120),
.B2(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_6),
.A2(n_145),
.B1(n_146),
.B2(n_149),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_6),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_6),
.A2(n_145),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_6),
.A2(n_61),
.B1(n_145),
.B2(n_300),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_6),
.A2(n_145),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_8),
.Y(n_163)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_8),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_8),
.Y(n_274)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_8),
.Y(n_339)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_8),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_9),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_9),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_9),
.A2(n_140),
.B1(n_279),
.B2(n_282),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_9),
.A2(n_34),
.B1(n_140),
.B2(n_309),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_9),
.A2(n_140),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_10),
.Y(n_128)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_10),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_10),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_11),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_11),
.A2(n_55),
.B1(n_115),
.B2(n_119),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_11),
.A2(n_55),
.B1(n_266),
.B2(n_269),
.Y(n_265)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_13),
.A2(n_95),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_13),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_13),
.A2(n_112),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_13),
.A2(n_112),
.B1(n_148),
.B2(n_228),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_13),
.A2(n_112),
.B1(n_182),
.B2(n_373),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_14),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_14),
.A2(n_159),
.B1(n_170),
.B2(n_258),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_14),
.B(n_72),
.C(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_14),
.B(n_104),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_14),
.B(n_272),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_14),
.B(n_86),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_14),
.B(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_16),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_16),
.A2(n_33),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_232),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_231),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_204),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_20),
.B(n_204),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_152),
.C(n_165),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_21),
.B(n_152),
.CI(n_165),
.CON(n_287),
.SN(n_287)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_87),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_22),
.B(n_88),
.C(n_122),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_23),
.B(n_48),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_36),
.B2(n_38),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_24),
.A2(n_38),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_24),
.A2(n_264),
.B1(n_272),
.B2(n_275),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_24),
.A2(n_308),
.B(n_311),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_24),
.A2(n_258),
.B(n_311),
.Y(n_332)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_25),
.A2(n_176),
.B1(n_184),
.B2(n_185),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_25),
.B(n_312),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_25),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_25),
.A2(n_162),
.B1(n_265),
.B2(n_372),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_27),
.Y(n_373)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g183 ( 
.A(n_29),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_29),
.Y(n_271)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_30),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_32),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_36),
.Y(n_347)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_37),
.B(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_41),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_42),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_43),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_59),
.B1(n_80),
.B2(n_86),
.Y(n_48)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_49),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g376 ( 
.A(n_51),
.Y(n_376)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AO22x2_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_104)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_53),
.Y(n_172)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_54),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_54),
.Y(n_322)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_59),
.A2(n_80),
.B1(n_86),
.B2(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_59),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_59),
.A2(n_86),
.B1(n_155),
.B2(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_59),
.B(n_299),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_71),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_68),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_62),
.Y(n_300)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_68),
.Y(n_303)
);

INVx5_ASAP7_75t_SL g361 ( 
.A(n_68),
.Y(n_361)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_71),
.A2(n_319),
.B(n_323),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_71),
.A2(n_169),
.B(n_323),
.Y(n_418)
);

AOI22x1_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_82),
.Y(n_359)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_86),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_86),
.B(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_122),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_109),
.B1(n_113),
.B2(n_114),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g196 ( 
.A(n_89),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_89),
.A2(n_113),
.B1(n_278),
.B2(n_393),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_104),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_95),
.B1(n_100),
.B2(n_102),
.Y(n_90)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_91),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_94),
.Y(n_380)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_96),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.Y(n_133)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_99),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_99),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_103),
.Y(n_214)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_103),
.Y(n_249)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_103),
.Y(n_256)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_103),
.Y(n_365)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

AOI22x1_ASAP7_75t_L g195 ( 
.A1(n_104),
.A2(n_196),
.B1(n_197),
.B2(n_203),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_104),
.A2(n_196),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_113),
.B(n_198),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_113),
.A2(n_393),
.B(n_394),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_114),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g375 ( 
.A1(n_119),
.A2(n_367),
.A3(n_376),
.B1(n_377),
.B2(n_381),
.Y(n_375)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_121),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_138),
.B(n_143),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_123),
.A2(n_133),
.B1(n_138),
.B2(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_124),
.B(n_144),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_124),
.A2(n_412),
.B(n_415),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_133),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_128),
.Y(n_137)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_133),
.B(n_258),
.Y(n_396)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_134),
.A2(n_247),
.A3(n_250),
.B1(n_252),
.B2(n_257),
.Y(n_246)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_143),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_151),
.Y(n_143)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_147),
.Y(n_251)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_151),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_151),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_160),
.B2(n_164),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_154),
.B(n_160),
.Y(n_222)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g381 ( 
.A(n_159),
.B(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_160),
.A2(n_164),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_189),
.C(n_195),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_166),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_175),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_167),
.B(n_175),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_168),
.A2(n_297),
.B(n_298),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_168),
.A2(n_173),
.B1(n_319),
.B2(n_358),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_168),
.A2(n_298),
.B(n_358),
.Y(n_389)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx11_ASAP7_75t_L g320 ( 
.A(n_172),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_176),
.Y(n_275)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_177),
.Y(n_305)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_183),
.Y(n_337)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_189),
.A2(n_190),
.B1(n_195),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_191),
.A2(n_230),
.B(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_195),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_196),
.A2(n_277),
.B(n_286),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_196),
.A2(n_286),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_196),
.B(n_197),
.Y(n_394)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx6_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_220),
.B2(n_221),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_215),
.B(n_219),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_216),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_288),
.B(n_443),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_287),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_235),
.B(n_287),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.C(n_241),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_236),
.A2(n_237),
.B1(n_240),
.B2(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_240),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_241),
.B(n_433),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_276),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_242),
.A2(n_243),
.B1(n_276),
.B2(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_245),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_262),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_246),
.A2(n_262),
.B1(n_263),
.B2(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_246),
.Y(n_405)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_SL g412 ( 
.A1(n_257),
.A2(n_258),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_SL g364 ( 
.A1(n_258),
.A2(n_365),
.B(n_366),
.Y(n_364)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_271),
.Y(n_310)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_276),
.Y(n_428)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_285),
.Y(n_368)
);

BUFx24_ASAP7_75t_SL g445 ( 
.A(n_287),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_421),
.B(n_440),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_400),
.B(n_420),
.Y(n_290)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_384),
.B(n_399),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_352),
.B(n_383),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_326),
.B(n_351),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_306),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_295),
.B(n_306),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_301),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_296),
.A2(n_301),
.B1(n_302),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_316),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_307),
.B(n_317),
.C(n_325),
.Y(n_353)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_324),
.B2(n_325),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_343),
.B(n_350),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_333),
.B(n_342),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_341),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_341),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_338),
.B(n_340),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_335),
.Y(n_345)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_340),
.A2(n_371),
.B(n_374),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_348),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_348),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_353),
.B(n_354),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_369),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_362),
.B2(n_363),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_362),
.C(n_369),
.Y(n_385)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_375),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_375),
.Y(n_390)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx8_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_385),
.B(n_386),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_387),
.A2(n_388),
.B1(n_391),
.B2(n_398),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_389),
.B(n_390),
.C(n_398),
.Y(n_401)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_391),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_395),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_396),
.C(n_397),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_401),
.B(n_402),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_409),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_406),
.B1(n_407),
.B2(n_408),
.Y(n_403)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_404),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_406),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_407),
.C(n_409),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_411),
.B1(n_416),
.B2(n_419),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_417),
.C(n_418),
.Y(n_431)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx8_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_416),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_435),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_424),
.A2(n_441),
.B(n_442),
.Y(n_440)
);

NOR2x1_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_432),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_432),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_429),
.C(n_431),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_426),
.B(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_429),
.A2(n_430),
.B1(n_431),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_431),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_437),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);


endmodule