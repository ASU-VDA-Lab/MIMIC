module real_jpeg_27908_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_334, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_334;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_0),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_0),
.A2(n_31),
.B1(n_33),
.B2(n_119),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_0),
.A2(n_45),
.B1(n_46),
.B2(n_119),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_0),
.A2(n_61),
.B1(n_63),
.B2(n_119),
.Y(n_253)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_1),
.Y(n_104)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_1),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_1),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_2),
.A2(n_31),
.B1(n_33),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_2),
.A2(n_49),
.B1(n_61),
.B2(n_63),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_31),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_3),
.A2(n_52),
.B1(n_61),
.B2(n_63),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_52),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_5),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_5),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_5),
.A2(n_37),
.B1(n_61),
.B2(n_63),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_7),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_7),
.A2(n_31),
.B1(n_33),
.B2(n_180),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_180),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_7),
.A2(n_61),
.B1(n_63),
.B2(n_180),
.Y(n_266)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_9),
.B(n_30),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_9),
.B(n_33),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_9),
.A2(n_33),
.B(n_218),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_178),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_9),
.A2(n_58),
.B(n_61),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_9),
.B(n_86),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_9),
.A2(n_104),
.B1(n_125),
.B2(n_266),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_10),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_10),
.A2(n_35),
.B1(n_61),
.B2(n_63),
.Y(n_193)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_12),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_12),
.A2(n_31),
.B1(n_33),
.B2(n_146),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_146),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_12),
.A2(n_61),
.B1(n_63),
.B2(n_146),
.Y(n_258)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_14),
.A2(n_31),
.B1(n_33),
.B2(n_47),
.Y(n_54)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_14),
.Y(n_217)
);

INVx11_ASAP7_75t_SL g62 ( 
.A(n_15),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_93),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_91),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_19),
.B(n_78),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_68),
.C(n_72),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_20),
.A2(n_21),
.B1(n_68),
.B2(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_39),
.B1(n_40),
.B2(n_67),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_23),
.A2(n_118),
.B(n_120),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_23),
.A2(n_38),
.B1(n_118),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_23),
.A2(n_38),
.B1(n_145),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_24),
.B(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_24),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_24),
.A2(n_83),
.B(n_121),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_24),
.A2(n_30),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_25),
.B(n_33),
.Y(n_191)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g177 ( 
.A(n_27),
.B(n_178),
.CON(n_177),
.SN(n_177)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_29),
.A2(n_31),
.B1(n_177),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_30),
.B(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

AOI32xp33_ASAP7_75t_L g214 ( 
.A1(n_31),
.A2(n_45),
.A3(n_215),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_34),
.A2(n_38),
.B(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_36),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_38),
.B(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_55),
.B2(n_66),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_55),
.C(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_43),
.A2(n_74),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_44),
.A2(n_53),
.B1(n_76),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_44),
.A2(n_53),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_44),
.A2(n_53),
.B1(n_174),
.B2(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_44),
.A2(n_53),
.B1(n_202),
.B2(n_222),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_46),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g219 ( 
.A(n_46),
.B(n_216),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_46),
.A2(n_59),
.B(n_178),
.C(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_50),
.A2(n_86),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_55),
.A2(n_66),
.B1(n_73),
.B2(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_64),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_56),
.A2(n_60),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_56),
.A2(n_111),
.B(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_56),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_56),
.A2(n_64),
.B(n_129),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_56),
.A2(n_60),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_56),
.A2(n_152),
.B(n_226),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_56),
.A2(n_60),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_56),
.A2(n_60),
.B1(n_225),
.B2(n_243),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_60),
.A2(n_110),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_60),
.B(n_178),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_61),
.Y(n_63)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_63),
.B(n_271),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_65),
.B(n_131),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_68),
.C(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_68),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_68),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_72),
.B(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_73),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_77),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_74),
.A2(n_77),
.B(n_87),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI321xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_313),
.A3(n_325),
.B1(n_331),
.B2(n_332),
.C(n_334),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_163),
.B(n_312),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_147),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_96),
.B(n_147),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_122),
.C(n_133),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_97),
.A2(n_98),
.B1(n_122),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_112),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_99),
.B(n_114),
.C(n_116),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_100),
.B(n_109),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_107),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_101),
.A2(n_126),
.B(n_193),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_102),
.A2(n_108),
.B(n_138),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_102),
.A2(n_103),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_108),
.Y(n_107)
);

INVx11_ASAP7_75t_L g267 ( 
.A(n_103),
.Y(n_267)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_104),
.A2(n_125),
.B1(n_136),
.B2(n_193),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_126),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_107),
.A2(n_125),
.B(n_253),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_122),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_132),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_124),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_128),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_124),
.A2(n_157),
.B(n_160),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_127),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_136),
.B(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_125),
.A2(n_258),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_128),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_133),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_142),
.C(n_143),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_134),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_139),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_142),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_161),
.B2(n_162),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_156),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_150),
.B(n_156),
.C(n_162),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_153),
.B(n_155),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_153),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_155),
.B(n_315),
.C(n_321),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_155),
.A2(n_315),
.B1(n_316),
.B2(n_330),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_155),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_161),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_306),
.B(n_311),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_206),
.B(n_292),
.C(n_305),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_194),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_166),
.B(n_194),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_181),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_168),
.B(n_169),
.C(n_181),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_176),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_176),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_178),
.B(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_179),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_189),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_183),
.B(n_187),
.C(n_189),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_192),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.C(n_200),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_195),
.A2(n_196),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_200),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.C(n_205),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_205),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_291),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_284),
.B(n_290),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_236),
.B(n_283),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_227),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_210),
.B(n_227),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_220),
.C(n_223),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_211),
.A2(n_212),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_214),
.Y(n_234)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_228),
.B(n_234),
.C(n_235),
.Y(n_285)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_277),
.B(n_282),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_254),
.B(n_276),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_246),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_239),
.B(n_246),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_240),
.A2(n_241),
.B1(n_244),
.B2(n_261),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_244),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_252),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_251),
.C(n_252),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_253),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_262),
.B(n_275),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_260),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_256),
.B(n_260),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_268),
.B(n_274),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_264),
.B(n_265),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_285),
.B(n_286),
.Y(n_290)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_294),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_303),
.B2(n_304),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_300),
.C(n_304),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_323),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_321),
.A2(n_322),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);


endmodule