module fake_jpeg_413_n_133 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_46),
.Y(n_58)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_31),
.B(n_37),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_SL g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_12),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_10),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_20),
.A2(n_2),
.B(n_3),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_6),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx12_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_17),
.A2(n_6),
.B1(n_13),
.B2(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_15),
.A2(n_6),
.B1(n_22),
.B2(n_16),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_24),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_14),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_72),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_36),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_67),
.B1(n_72),
.B2(n_64),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_25),
.B(n_26),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_40),
.A3(n_52),
.B1(n_42),
.B2(n_34),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_42),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_86),
.B(n_71),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_35),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_57),
.B(n_59),
.Y(n_96)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_90),
.B1(n_57),
.B2(n_61),
.Y(n_100)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_74),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_55),
.B(n_60),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_99),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_85),
.B(n_86),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_78),
.C(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_110),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.C(n_104),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_79),
.B1(n_67),
.B2(n_63),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_96),
.B(n_99),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_114),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_104),
.B(n_95),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_97),
.C(n_98),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_102),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_116),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_111),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_116),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_117),
.C(n_101),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_106),
.Y(n_125)
);

AOI211xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_121),
.B(n_122),
.C(n_109),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_108),
.C(n_93),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_128),
.B(n_129),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_93),
.C(n_103),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_70),
.B(n_61),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_70),
.B1(n_77),
.B2(n_64),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_77),
.Y(n_133)
);


endmodule