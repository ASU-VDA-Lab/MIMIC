module fake_netlist_5_2571_n_39 (n_8, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_6, n_1, n_39);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_6;
input n_1;

output n_39;

wire n_29;
wire n_16;
wire n_12;
wire n_36;
wire n_25;
wire n_18;
wire n_27;
wire n_22;
wire n_10;
wire n_24;
wire n_28;
wire n_21;
wire n_34;
wire n_38;
wire n_35;
wire n_32;
wire n_11;
wire n_17;
wire n_19;
wire n_37;
wire n_26;
wire n_15;
wire n_30;
wire n_33;
wire n_14;
wire n_31;
wire n_23;
wire n_13;
wire n_20;

INVx2_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx5p33_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

OAI221xp5_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.C(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_14),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_18),
.B1(n_12),
.B2(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_19),
.Y(n_31)
);

OR2x4_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_33),
.Y(n_34)
);

OAI221xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_30),
.B1(n_28),
.B2(n_21),
.C(n_18),
.Y(n_35)
);

NOR2xp67_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_5),
.Y(n_36)
);

NOR3xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_23),
.C(n_15),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_10),
.B1(n_37),
.B2(n_32),
.Y(n_39)
);


endmodule