module fake_jpeg_28460_n_151 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_68),
.Y(n_73)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_0),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_53),
.Y(n_77)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_64),
.Y(n_87)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_57),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_49),
.B1(n_55),
.B2(n_60),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_86),
.B(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_87),
.B(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_53),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_55),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_97),
.C(n_25),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_51),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_59),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_62),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_5),
.C(n_6),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_3),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_85),
.B1(n_56),
.B2(n_61),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_108),
.B1(n_7),
.B2(n_8),
.Y(n_128)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_62),
.B1(n_58),
.B2(n_57),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_109),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_85),
.B1(n_56),
.B2(n_62),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_29),
.B1(n_37),
.B2(n_11),
.Y(n_127)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_112),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_4),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_114),
.B(n_117),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_45),
.B(n_24),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_21),
.C(n_40),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_119),
.C(n_28),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_42),
.B(n_20),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_18),
.C(n_39),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_120),
.B(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_118),
.B(n_17),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_128),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_16),
.C(n_38),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_111),
.C(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_124),
.B(n_126),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_6),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_7),
.B(n_8),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_113),
.B(n_110),
.C(n_31),
.D(n_32),
.Y(n_141)
);

AOI22x1_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_141),
.Y(n_144)
);

BUFx4f_ASAP7_75t_SL g140 ( 
.A(n_132),
.Y(n_140)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_133),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_130),
.C(n_138),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_144),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_136),
.B1(n_121),
.B2(n_137),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_125),
.B1(n_135),
.B2(n_142),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_125),
.C(n_142),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_131),
.Y(n_151)
);


endmodule