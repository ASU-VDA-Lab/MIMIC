module real_jpeg_15560_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_11;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_105;
wire n_40;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g79 ( 
.A(n_0),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_0),
.Y(n_119)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_1),
.Y(n_217)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_2),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_3),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_23),
.B1(n_96),
.B2(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_3),
.B(n_188),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_3),
.A2(n_202),
.A3(n_205),
.B1(n_206),
.B2(n_211),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_3),
.B(n_117),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_3),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_3),
.B(n_256),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_4),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_4),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22x1_ASAP7_75t_L g126 ( 
.A1(n_5),
.A2(n_60),
.B1(n_127),
.B2(n_130),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_5),
.A2(n_60),
.B1(n_227),
.B2(n_230),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_6),
.A2(n_109),
.B1(n_110),
.B2(n_115),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_6),
.B(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_6),
.A2(n_109),
.B1(n_173),
.B2(n_177),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_7),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_7),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_8),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_9),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_196),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_194),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_166),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_13),
.B(n_166),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_105),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_63),
.B1(n_103),
.B2(n_104),
.Y(n_14)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_15),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_43),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_29),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_19),
.B(n_44),
.Y(n_219)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_23),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_23),
.B(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_23),
.B(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_28),
.Y(n_121)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_29),
.Y(n_256)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_30),
.B(n_58),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_30),
.B(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_36),
.B1(n_38),
.B2(n_42),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_37),
.Y(n_210)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_37),
.Y(n_229)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_40),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_43),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_58),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_44),
.B(n_172),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_51),
.B2(n_55),
.Y(n_45)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_56),
.Y(n_204)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_87),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_64),
.A2(n_87),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_64),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_71),
.A3(n_74),
.B1(n_80),
.B2(n_84),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_68),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_72),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_84),
.B(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_87),
.Y(n_192)
);

OA21x2_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B(n_99),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_92),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_92),
.B(n_149),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_98),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_99),
.A2(n_222),
.B(n_225),
.Y(n_221)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_142),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_125),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_117),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_147),
.B(n_149),
.C(n_154),
.Y(n_146)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NOR2x1p5_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_117),
.B(n_126),
.Y(n_182)
);

AO22x2_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_135),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_133),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_133),
.Y(n_190)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_158),
.B2(n_159),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_145),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_146),
.B(n_225),
.Y(n_254)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_153),
.Y(n_232)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_181),
.C(n_191),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_167),
.A2(n_168),
.B1(n_181),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_181),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_190),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_191),
.B(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_266),
.B(n_272),
.Y(n_197)
);

AOI21x1_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_239),
.B(n_265),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_220),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_L g265 ( 
.A(n_200),
.B(n_220),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_218),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_201),
.B(n_218),
.Y(n_263)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_233),
.Y(n_220)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_221),
.Y(n_271)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_226),
.Y(n_252)
);

INVx4_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_236),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_236),
.B(n_237),
.C(n_271),
.Y(n_270)
);

OAI21x1_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_258),
.B(n_264),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_253),
.B(n_257),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_251),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_255),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_263),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_270),
.Y(n_272)
);


endmodule