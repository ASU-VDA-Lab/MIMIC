module fake_jpeg_17089_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_11),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_51),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_19),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_33),
.B1(n_17),
.B2(n_24),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_65),
.Y(n_85)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_33),
.B1(n_17),
.B2(n_24),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_33),
.B1(n_17),
.B2(n_24),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_33),
.B1(n_32),
.B2(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_43),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_36),
.C(n_56),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_81),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_36),
.C(n_39),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_103),
.B1(n_106),
.B2(n_25),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_86),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_97),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_47),
.B(n_23),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_87),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_90),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_92),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_45),
.B1(n_37),
.B2(n_38),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_100),
.B1(n_20),
.B2(n_25),
.Y(n_130)
);

OR2x4_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_26),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_28),
.B(n_34),
.Y(n_113)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_45),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_63),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_98),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_26),
.C(n_22),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_58),
.B1(n_50),
.B2(n_35),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_48),
.A2(n_58),
.B1(n_50),
.B2(n_47),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_105),
.Y(n_128)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_57),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_111),
.B1(n_116),
.B2(n_117),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_75),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_20),
.B(n_95),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_69),
.B(n_68),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_81),
.B(n_83),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_66),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_29),
.B1(n_21),
.B2(n_30),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_25),
.C(n_27),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_27),
.Y(n_163)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_29),
.B1(n_21),
.B2(n_30),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_95),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_16),
.B1(n_27),
.B2(n_25),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_29),
.B1(n_21),
.B2(n_20),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_100),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_88),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_138),
.B(n_140),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_80),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_141),
.B(n_142),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_162),
.B(n_115),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_130),
.B1(n_101),
.B2(n_100),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_149),
.B1(n_108),
.B2(n_123),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_74),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_156),
.B(n_165),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_158),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_79),
.B1(n_100),
.B2(n_101),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_157),
.B1(n_130),
.B2(n_112),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_93),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_93),
.B1(n_74),
.B2(n_96),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_67),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_26),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_159),
.B(n_152),
.Y(n_199)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

AOI222xp33_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_16),
.B1(n_27),
.B2(n_12),
.C1(n_15),
.C2(n_13),
.Y(n_161)
);

XNOR2x1_ASAP7_75t_SL g183 ( 
.A(n_161),
.B(n_117),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_0),
.B(n_1),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_137),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_16),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_0),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

BUFx8_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_168),
.B(n_0),
.Y(n_220)
);

NOR4xp25_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_119),
.C(n_113),
.D(n_115),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_170),
.A2(n_174),
.B(n_177),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_171),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_103),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_112),
.B(n_129),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_120),
.B(n_109),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_180),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_116),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_182),
.Y(n_226)
);

CKINVDCx12_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_183),
.A2(n_194),
.B(n_1),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_141),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_193),
.C(n_162),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_185),
.B(n_199),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_137),
.A2(n_126),
.B1(n_133),
.B2(n_111),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_188),
.A2(n_191),
.B1(n_197),
.B2(n_154),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_156),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_189),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_143),
.A2(n_133),
.B1(n_111),
.B2(n_107),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_107),
.C(n_127),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_114),
.B(n_131),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_143),
.A2(n_121),
.B1(n_102),
.B2(n_105),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_203),
.C(n_216),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_140),
.C(n_138),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_SL g204 ( 
.A(n_183),
.B(n_159),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_185),
.B1(n_178),
.B2(n_179),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_195),
.A2(n_153),
.B1(n_148),
.B2(n_149),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_205),
.A2(n_206),
.B1(n_211),
.B2(n_215),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_195),
.A2(n_148),
.B1(n_149),
.B2(n_114),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_165),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_180),
.A2(n_148),
.B1(n_131),
.B2(n_160),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_117),
.B1(n_127),
.B2(n_84),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_167),
.C(n_139),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_219),
.B1(n_225),
.B2(n_227),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_224),
.C(n_193),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_171),
.A2(n_166),
.B1(n_77),
.B2(n_2),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_178),
.Y(n_244)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_222),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_179),
.B(n_200),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_77),
.C(n_2),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_181),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_228),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_3),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

OAI31xp33_ASAP7_75t_SL g232 ( 
.A1(n_221),
.A2(n_194),
.A3(n_174),
.B(n_177),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_241),
.Y(n_262)
);

OAI21x1_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_170),
.B(n_199),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_237),
.B(n_253),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_212),
.A2(n_211),
.B1(n_219),
.B2(n_201),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_244),
.B(n_229),
.CI(n_220),
.CON(n_273),
.SN(n_273)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_248),
.C(n_249),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_250),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_173),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_188),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_225),
.A2(n_191),
.B1(n_175),
.B2(n_169),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_175),
.C(n_197),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_254),
.B(n_261),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_269),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_230),
.B(n_248),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_257),
.A2(n_238),
.B(n_250),
.Y(n_286)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_234),
.A2(n_216),
.B1(n_214),
.B2(n_205),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_272),
.B1(n_240),
.B2(n_232),
.Y(n_274)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_265),
.B(n_266),
.Y(n_284)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_203),
.C(n_207),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_270),
.C(n_271),
.Y(n_275)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_224),
.C(n_208),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_215),
.C(n_210),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_240),
.A2(n_206),
.B1(n_217),
.B2(n_213),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_247),
.Y(n_281)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_249),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_283),
.C(n_256),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_288),
.Y(n_291)
);

XNOR2x1_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_244),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_281),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_241),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_262),
.B(n_239),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_286),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_187),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_287),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_245),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_258),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_289),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_258),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_286),
.B(n_276),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_283),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_267),
.B(n_236),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_295),
.A2(n_300),
.B(n_285),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_270),
.C(n_268),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_299),
.C(n_278),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_263),
.B1(n_238),
.B2(n_262),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_273),
.C(n_198),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_239),
.B(n_198),
.Y(n_300)
);

OAI322xp33_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_273),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_303),
.B(n_4),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_282),
.Y(n_305)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_307),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_296),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_314),
.B(n_299),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_309),
.B(n_310),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_274),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_312),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_313),
.A2(n_304),
.A3(n_298),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_4),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_318),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_313),
.B1(n_7),
.B2(n_8),
.Y(n_323)
);

AOI31xp33_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_297),
.A3(n_304),
.B(n_302),
.Y(n_318)
);

A2O1A1O1Ixp25_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_302),
.B(n_308),
.C(n_306),
.D(n_309),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_323),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_294),
.C(n_5),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_325),
.A2(n_317),
.B(n_321),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_327),
.B(n_324),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_326),
.Y(n_329)
);

NOR3xp33_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_322),
.C(n_316),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_330),
.Y(n_331)
);


endmodule