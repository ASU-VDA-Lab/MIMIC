module fake_jpeg_5545_n_153 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_153);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_3),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_16),
.B1(n_14),
.B2(n_21),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_9),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_27),
.B(n_11),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_34),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_12),
.B(n_17),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_13),
.B(n_19),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_16),
.B1(n_14),
.B2(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_24),
.A2(n_16),
.B1(n_14),
.B2(n_19),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_50),
.B(n_37),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_31),
.B(n_32),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_32),
.B1(n_39),
.B2(n_35),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_64),
.B1(n_65),
.B2(n_41),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_55),
.B(n_59),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_40),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_22),
.B1(n_16),
.B2(n_14),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_24),
.B1(n_26),
.B2(n_22),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

NAND2x1_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_45),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_50),
.B1(n_49),
.B2(n_51),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_73),
.B1(n_76),
.B2(n_40),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_45),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_48),
.C(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_60),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_40),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_58),
.B1(n_77),
.B2(n_48),
.Y(n_98)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_67),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_75),
.C(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_74),
.Y(n_88)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_89),
.B(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_89),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_73),
.B1(n_70),
.B2(n_69),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_80),
.B1(n_87),
.B2(n_82),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_96),
.C(n_90),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_78),
.C(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_103),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_102),
.B(n_84),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_66),
.B(n_67),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_43),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_85),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_112),
.B(n_115),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_114),
.B1(n_18),
.B2(n_28),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_111),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_113),
.C(n_105),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_85),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_33),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_11),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_22),
.B1(n_42),
.B2(n_27),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_12),
.B(n_17),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_93),
.B(n_103),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_17),
.B(n_36),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_99),
.B1(n_42),
.B2(n_27),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_120),
.B1(n_121),
.B2(n_126),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_26),
.B1(n_13),
.B2(n_28),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_26),
.B1(n_36),
.B2(n_13),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_127),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_28),
.B1(n_18),
.B2(n_43),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_111),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_110),
.C(n_115),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_132),
.B(n_135),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_108),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_134),
.Y(n_142)
);

NOR2xp67_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_106),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_111),
.B1(n_109),
.B2(n_18),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_137),
.B(n_0),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_124),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_6),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_129),
.B1(n_136),
.B2(n_130),
.Y(n_143)
);

OAI321xp33_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_147),
.A3(n_146),
.B1(n_8),
.B2(n_3),
.C(n_4),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_6),
.B(n_10),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_145),
.C(n_1),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_23),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_148),
.A2(n_149),
.B(n_150),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_0),
.Y(n_149)
);

OAI221xp5_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_1),
.B1(n_4),
.B2(n_25),
.C(n_23),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);


endmodule