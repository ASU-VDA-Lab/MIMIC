module fake_jpeg_8782_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_0),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_34),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_16),
.B1(n_33),
.B2(n_32),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_48),
.A2(n_75),
.B1(n_25),
.B2(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_64),
.Y(n_89)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_61),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_16),
.B1(n_33),
.B2(n_30),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_36),
.A2(n_16),
.B1(n_33),
.B2(n_32),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_31),
.B(n_35),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_33),
.B1(n_24),
.B2(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_71),
.Y(n_79)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_22),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_35),
.B1(n_31),
.B2(n_30),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_40),
.A2(n_35),
.B1(n_31),
.B2(n_24),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_74),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_41),
.A2(n_18),
.B1(n_27),
.B2(n_22),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_47),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_37),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_82),
.A2(n_85),
.B(n_86),
.Y(n_124)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_83),
.B(n_87),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_36),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_90),
.A2(n_26),
.B(n_20),
.Y(n_137)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_47),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_27),
.B(n_18),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_19),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_38),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_110),
.Y(n_130)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_105),
.Y(n_123)
);

CKINVDCx12_ASAP7_75t_R g105 ( 
.A(n_69),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_49),
.B1(n_70),
.B2(n_67),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_38),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_108),
.Y(n_140)
);

CKINVDCx12_ASAP7_75t_R g108 ( 
.A(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_26),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_49),
.A2(n_29),
.B1(n_21),
.B2(n_37),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_25),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_56),
.B(n_26),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_60),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_59),
.B(n_26),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_77),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_120),
.A2(n_137),
.B(n_138),
.Y(n_181)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_122),
.Y(n_158)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_13),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_126),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_127),
.B(n_97),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_99),
.B1(n_95),
.B2(n_116),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_132),
.B(n_88),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_147),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_0),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_20),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_143),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g142 ( 
.A1(n_85),
.A2(n_61),
.B(n_67),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_142),
.A2(n_93),
.B1(n_84),
.B2(n_115),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_20),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_86),
.B(n_1),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_89),
.B(n_88),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_20),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_110),
.Y(n_170)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_155),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_141),
.A2(n_81),
.B1(n_96),
.B2(n_87),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_154),
.B1(n_135),
.B2(n_180),
.Y(n_187)
);

AO22x1_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_114),
.B1(n_101),
.B2(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_163),
.B1(n_175),
.B2(n_115),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_80),
.B1(n_114),
.B2(n_99),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_145),
.B1(n_93),
.B2(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_161),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_176),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_114),
.B1(n_79),
.B2(n_84),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_166),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_125),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_104),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_170),
.Y(n_196)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_79),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_173),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_93),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_174),
.B(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_102),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_138),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_124),
.B(n_15),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_84),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_119),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_124),
.C(n_119),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_188),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_127),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_186),
.B(n_187),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_146),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_190),
.B(n_198),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_154),
.A2(n_142),
.B1(n_120),
.B2(n_137),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_169),
.B1(n_176),
.B2(n_153),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_199),
.B1(n_203),
.B2(n_212),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_164),
.A2(n_154),
.B1(n_163),
.B2(n_157),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_171),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_210),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_145),
.B(n_126),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_207),
.A2(n_19),
.B(n_10),
.Y(n_239)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_149),
.B(n_129),
.C(n_109),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_152),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_164),
.A2(n_129),
.B1(n_113),
.B2(n_115),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_155),
.B(n_117),
.C(n_122),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_147),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_209),
.Y(n_248)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_218),
.B(n_221),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_178),
.B(n_160),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_184),
.B(n_208),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_194),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_206),
.A2(n_159),
.B1(n_166),
.B2(n_161),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_222),
.A2(n_231),
.B1(n_237),
.B2(n_189),
.Y(n_242)
);

AOI32xp33_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_169),
.A3(n_165),
.B1(n_150),
.B2(n_148),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_189),
.A3(n_202),
.B1(n_200),
.B2(n_192),
.C1(n_195),
.C2(n_182),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_227),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_185),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_193),
.B(n_151),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_228),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_150),
.B1(n_117),
.B2(n_103),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_240),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_136),
.B1(n_133),
.B2(n_152),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_1),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_7),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_182),
.B(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_204),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_243),
.B(n_234),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_244),
.B1(n_217),
.B2(n_214),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_196),
.B1(n_204),
.B2(n_210),
.Y(n_244)
);

HAxp5_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_238),
.CON(n_263),
.SN(n_263)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_188),
.B1(n_186),
.B2(n_91),
.Y(n_246)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_226),
.A2(n_209),
.B1(n_91),
.B2(n_19),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_247),
.A2(n_237),
.B1(n_222),
.B2(n_229),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_253),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_134),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_227),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_152),
.C(n_61),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_259),
.C(n_260),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_1),
.C(n_2),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_7),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_272),
.B1(n_261),
.B2(n_232),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_269),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_240),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_265),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_235),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_271),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_262),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_216),
.B(n_252),
.Y(n_284)
);

BUFx12_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_252),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_253),
.C(n_248),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_277),
.C(n_279),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_234),
.C(n_220),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_232),
.C(n_214),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_261),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_254),
.B1(n_245),
.B2(n_247),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_281),
.A2(n_287),
.B1(n_266),
.B2(n_280),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_289),
.B1(n_260),
.B2(n_259),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_284),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_276),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_6),
.C(n_3),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_239),
.B1(n_242),
.B2(n_250),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_272),
.A2(n_265),
.B1(n_270),
.B2(n_279),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_290),
.B(n_294),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_292),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_278),
.A2(n_244),
.B(n_225),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_266),
.A2(n_264),
.B1(n_277),
.B2(n_263),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_301),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_271),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_287),
.A2(n_268),
.B1(n_267),
.B2(n_275),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_255),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_267),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_283),
.A2(n_281),
.B(n_288),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_8),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_288),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_310),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_297),
.Y(n_310)
);

AOI21xp33_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_286),
.B(n_4),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_311),
.A2(n_301),
.B(n_4),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_15),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_302),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_319),
.A3(n_320),
.B1(n_312),
.B2(n_306),
.C1(n_308),
.C2(n_8),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_318),
.B(n_315),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_298),
.B1(n_295),
.B2(n_300),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_305),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g325 ( 
.A1(n_321),
.A2(n_322),
.A3(n_323),
.B1(n_5),
.B2(n_6),
.C1(n_8),
.C2(n_13),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_5),
.C(n_6),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_325),
.C(n_14),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_14),
.Y(n_328)
);


endmodule