module real_jpeg_5628_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_1),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_1),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_1),
.B(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_1),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_1),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_1),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_2),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_2),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_2),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_2),
.B(n_119),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_2),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_2),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_3),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_3),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_3),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_3),
.B(n_366),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_4),
.Y(n_129)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_4),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_5),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_5),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_5),
.B(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_5),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_5),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_5),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_5),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_5),
.B(n_357),
.Y(n_356)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_7),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_7),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_7),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_7),
.B(n_57),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_7),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_7),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g432 ( 
.A(n_7),
.B(n_433),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_8),
.Y(n_91)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_8),
.Y(n_135)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_9),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g444 ( 
.A(n_9),
.Y(n_444)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_11),
.B(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_11),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_11),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_11),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_11),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_11),
.B(n_310),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_11),
.B(n_444),
.Y(n_461)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_12),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_12),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_12),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_12),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_12),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_13),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_13),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_42),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_14),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_14),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_14),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_14),
.B(n_261),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_14),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_14),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_14),
.B(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_15),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_15),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_15),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_15),
.B(n_102),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_450),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_423),
.B(n_449),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_313),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_228),
.B(n_269),
.C(n_270),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_197),
.B(n_227),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_22),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_157),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_23),
.B(n_157),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_105),
.C(n_141),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_24),
.B(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_69),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_25),
.B(n_70),
.C(n_84),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_47),
.C(n_60),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_26),
.B(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_41),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_36),
.B2(n_40),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_28),
.A2(n_29),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_28),
.A2(n_29),
.B1(n_71),
.B2(n_72),
.Y(n_470)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_29),
.B(n_36),
.C(n_41),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_29),
.B(n_206),
.C(n_432),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OR2x2_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_49),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_30),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_30),
.B(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_34),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_34),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_34),
.Y(n_334)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_35),
.Y(n_195)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_35),
.Y(n_216)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_38),
.Y(n_167)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_39),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_39),
.Y(n_213)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_39),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_39),
.Y(n_311)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_45),
.B(n_108),
.Y(n_381)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_47),
.A2(n_60),
.B1(n_61),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_47),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.C(n_54),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_48),
.A2(n_54),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_48),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_48),
.A2(n_206),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_48),
.A2(n_206),
.B1(n_432),
.B2(n_434),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_48),
.B(n_127),
.C(n_279),
.Y(n_437)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_50),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_51),
.B(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_54),
.Y(n_207)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_58),
.Y(n_264)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_59),
.Y(n_294)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_62),
.A2(n_177),
.B1(n_178),
.B2(n_180),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_62),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_180),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_62),
.B(n_178),
.C(n_181),
.Y(n_267)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_84),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_72),
.B(n_78),
.C(n_82),
.Y(n_196)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_73),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_75),
.Y(n_220)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_79),
.B(n_127),
.Y(n_329)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_80),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_86),
.B(n_88),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_85),
.B(n_93),
.C(n_99),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_99),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_100),
.B(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_103),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_105),
.B(n_141),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_122),
.C(n_124),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_106),
.A2(n_122),
.B1(n_123),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_111),
.C(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_108),
.B(n_388),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_115),
.B1(n_116),
.B2(n_121),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_115),
.A2(n_116),
.B1(n_247),
.B2(n_251),
.Y(n_246)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_116),
.B(n_178),
.C(n_248),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_124),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.C(n_136),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_125),
.A2(n_126),
.B1(n_410),
.B2(n_411),
.Y(n_409)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_127),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_127),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_127),
.A2(n_237),
.B1(n_279),
.B2(n_282),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_127),
.B(n_240),
.C(n_245),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx8_ASAP7_75t_L g324 ( 
.A(n_129),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_130),
.A2(n_131),
.B1(n_136),
.B2(n_137),
.Y(n_411)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_135),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_135),
.Y(n_385)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_156),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_144),
.C(n_156),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_151),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_152),
.C(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_150),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_150),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_152),
.A2(n_292),
.B1(n_295),
.B2(n_296),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_152),
.Y(n_296)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_158),
.B(n_160),
.C(n_183),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_183),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_174),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_162),
.B(n_163),
.C(n_174),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_164),
.Y(n_235)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_169),
.B(n_172),
.C(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_181),
.B2(n_182),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_177),
.A2(n_178),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_177),
.A2(n_178),
.B1(n_321),
.B2(n_322),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_178),
.B(n_321),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_181),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_181),
.A2(n_182),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_182),
.B(n_443),
.C(n_446),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_184),
.B(n_186),
.C(n_187),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_196),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_189),
.B(n_191),
.C(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_225),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_198),
.B(n_225),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.C(n_222),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_199),
.A2(n_200),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_203),
.B(n_222),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.C(n_221),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_204),
.B(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_208),
.B(n_221),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.C(n_217),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_209),
.A2(n_210),
.B1(n_217),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_214),
.B(n_341),
.Y(n_340)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_216),
.Y(n_366)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_217),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_218),
.B(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_218),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_229),
.B(n_271),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_231),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_272),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_231),
.B(n_272),
.Y(n_422)
);

FAx1_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_252),
.CI(n_268),
.CON(n_231),
.SN(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_246),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_234),
.B(n_236),
.C(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_245),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_243),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_243),
.A2(n_245),
.B1(n_469),
.B2(n_470),
.Y(n_468)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_248),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_255),
.C(n_257),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_267),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_265),
.B2(n_266),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_260),
.B(n_265),
.C(n_267),
.Y(n_303)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_265),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_265),
.A2(n_266),
.B1(n_309),
.B2(n_312),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_266),
.B(n_305),
.C(n_312),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_273),
.B(n_275),
.C(n_298),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_298),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_283),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_276),
.B(n_284),
.C(n_285),
.Y(n_448)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_279),
.Y(n_282)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_291),
.B2(n_297),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_287),
.B(n_292),
.C(n_296),
.Y(n_438)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_291),
.Y(n_297)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_299),
.B(n_303),
.C(n_304),
.Y(n_426)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

AO22x1_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_309),
.Y(n_312)
);

INVx6_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

OAI31xp33_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_419),
.A3(n_420),
.B(n_422),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_413),
.B(n_418),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_400),
.B(n_412),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_360),
.B(n_399),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_343),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_318),
.B(n_343),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_330),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_319),
.B(n_331),
.C(n_340),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_325),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_320),
.B(n_326),
.C(n_329),
.Y(n_408)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_340),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.C(n_338),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_332),
.B(n_345),
.Y(n_344)
);

INVx11_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_335),
.A2(n_336),
.B1(n_338),
.B2(n_339),
.Y(n_345)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.C(n_359),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_344),
.B(n_396),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_346),
.A2(n_347),
.B1(n_359),
.B2(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_355),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_348),
.A2(n_349),
.B1(n_355),
.B2(n_356),
.Y(n_369)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_359),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_393),
.B(n_398),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_379),
.B(n_392),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_370),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_370),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_369),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_367),
.C(n_369),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_376),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_371),
.A2(n_372),
.B1(n_376),
.B2(n_377),
.Y(n_390)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_377),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_386),
.B(n_391),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx8_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_390),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_390),
.Y(n_391)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_395),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_402),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_403),
.A2(n_404),
.B1(n_406),
.B2(n_407),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_408),
.C(n_409),
.Y(n_417)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_417),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_417),
.Y(n_418)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_415),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_425),
.Y(n_449)
);

BUFx24_ASAP7_75t_SL g474 ( 
.A(n_425),
.Y(n_474)
);

FAx1_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_427),
.CI(n_439),
.CON(n_425),
.SN(n_425)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_427),
.C(n_439),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_435),
.B2(n_436),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_437),
.C(n_438),
.Y(n_456)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_432),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_448),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_441),
.B(n_442),
.C(n_448),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.Y(n_442)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_446),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_471),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_453),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_466),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_461),
.A2(n_462),
.B1(n_464),
.B2(n_465),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_461),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_462),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);


endmodule