module fake_jpeg_19620_n_312 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_8),
.B(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_49),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_43),
.B(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_18),
.B(n_2),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_50),
.Y(n_81)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_22),
.B(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_22),
.Y(n_77)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_56),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_36),
.B1(n_19),
.B2(n_28),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_77),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_36),
.B1(n_19),
.B2(n_29),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_60),
.A2(n_61),
.B1(n_89),
.B2(n_95),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_19),
.B1(n_30),
.B2(n_18),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_62),
.Y(n_96)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_33),
.B1(n_30),
.B2(n_24),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_66),
.A2(n_70),
.B1(n_94),
.B2(n_4),
.Y(n_116)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_33),
.B1(n_24),
.B2(n_34),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_74),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_38),
.B1(n_37),
.B2(n_31),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_78),
.A2(n_91),
.B1(n_2),
.B2(n_3),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_35),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_37),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_48),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_28),
.B1(n_35),
.B2(n_26),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_35),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_48),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_26),
.B1(n_23),
.B2(n_28),
.Y(n_91)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_20),
.B1(n_27),
.B2(n_39),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_42),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_97),
.Y(n_148)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_109),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_20),
.B(n_39),
.C(n_4),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_106),
.B(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_108),
.B(n_64),
.Y(n_142)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_112),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_80),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_48),
.B(n_23),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_12),
.C(n_13),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_117),
.B1(n_118),
.B2(n_126),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_116),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_57),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_57),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_57),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_124),
.Y(n_135)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_8),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_127),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_59),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_9),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_129),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_59),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_68),
.B(n_11),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_11),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_91),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_79),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_87),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_136),
.A2(n_163),
.B(n_108),
.Y(n_184)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_155),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_71),
.C(n_75),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_126),
.C(n_128),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_71),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_121),
.A2(n_72),
.B1(n_86),
.B2(n_63),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_96),
.B1(n_129),
.B2(n_123),
.Y(n_165)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_86),
.B1(n_13),
.B2(n_14),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_63),
.B1(n_58),
.B2(n_65),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_130),
.B1(n_114),
.B2(n_99),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_96),
.B(n_65),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_160),
.Y(n_169)
);

OR2x2_ASAP7_75t_SL g157 ( 
.A(n_106),
.B(n_14),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_14),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_158),
.B(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_102),
.B(n_15),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_175),
.B1(n_154),
.B2(n_151),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_112),
.B1(n_130),
.B2(n_100),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_167),
.A2(n_179),
.B(n_182),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_150),
.B(n_160),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_171),
.Y(n_202)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_103),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_178),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_139),
.B(n_111),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_141),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_152),
.Y(n_182)
);

BUFx24_ASAP7_75t_SL g183 ( 
.A(n_146),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_183),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_187),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_131),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_190),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_142),
.C(n_143),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_159),
.C(n_148),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_136),
.B(n_107),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_191),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_99),
.Y(n_194)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_145),
.A2(n_100),
.B1(n_105),
.B2(n_98),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_195),
.A2(n_140),
.B1(n_134),
.B2(n_164),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_109),
.Y(n_196)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_147),
.B(n_158),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_198),
.A2(n_199),
.B(n_211),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_157),
.B(n_143),
.C(n_163),
.D(n_147),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_135),
.B(n_156),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_219),
.B(n_178),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_223),
.C(n_169),
.Y(n_235)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_148),
.B(n_159),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_165),
.B1(n_168),
.B2(n_175),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_168),
.A2(n_134),
.B1(n_162),
.B2(n_105),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_180),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_216),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_162),
.B(n_138),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_138),
.C(n_187),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_198),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_174),
.Y(n_225)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_179),
.Y(n_228)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_215),
.B(n_173),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_234),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_223),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_241),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_207),
.C(n_218),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_210),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_237),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_173),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_205),
.B(n_169),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_172),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_185),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_245),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_238),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_244),
.A2(n_211),
.B1(n_213),
.B2(n_197),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_243),
.B1(n_200),
.B2(n_229),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_256),
.C(n_246),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_235),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_212),
.B1(n_204),
.B2(n_220),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_219),
.B1(n_200),
.B2(n_203),
.Y(n_268)
);

INVxp33_ASAP7_75t_SL g260 ( 
.A(n_226),
.Y(n_260)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_224),
.C(n_238),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_230),
.C(n_229),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_245),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_276),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_170),
.Y(n_266)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_262),
.B(n_226),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_269),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_273),
.C(n_246),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_274),
.B(n_247),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_248),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_272),
.A2(n_255),
.B(n_258),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_243),
.C(n_242),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_248),
.A2(n_257),
.B(n_199),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_188),
.C(n_230),
.Y(n_275)
);

OAI21x1_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_201),
.B(n_251),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_250),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_283),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_286),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_273),
.C(n_261),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_271),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_269),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_288),
.B(n_264),
.Y(n_297)
);

AOI21xp33_ASAP7_75t_SL g292 ( 
.A1(n_287),
.A2(n_274),
.B(n_268),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_263),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_263),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_294),
.A2(n_295),
.B(n_267),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_298),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_283),
.C(n_286),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_277),
.C(n_279),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_300),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_279),
.C(n_281),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_301),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_294),
.B(n_271),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_166),
.B(n_222),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_304),
.A2(n_240),
.A3(n_249),
.B1(n_186),
.B2(n_166),
.C1(n_176),
.C2(n_192),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_307),
.C(n_308),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_302),
.A2(n_240),
.B1(n_182),
.B2(n_176),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_309),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_310),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_311),
.A2(n_305),
.B(n_191),
.Y(n_312)
);


endmodule