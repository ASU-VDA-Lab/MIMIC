module fake_netlist_1_8424_n_50 (n_11, n_1, n_2, n_13, n_16, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_50);
input n_11;
input n_1;
input n_2;
input n_13;
input n_16;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_50;
wire n_45;
wire n_38;
wire n_20;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_48;
wire n_46;
wire n_25;
wire n_30;
wire n_26;
wire n_33;
wire n_49;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
OAI22xp5_ASAP7_75t_SL g17 ( .A1(n_12), .A2(n_8), .B1(n_6), .B2(n_2), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_9), .B(n_4), .Y(n_18) );
BUFx12f_ASAP7_75t_L g19 ( .A(n_4), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_3), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_11), .Y(n_22) );
AOI22xp5_ASAP7_75t_L g23 ( .A1(n_7), .A2(n_10), .B1(n_13), .B2(n_11), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_10), .B(n_0), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_8), .Y(n_25) );
OAI22xp5_ASAP7_75t_L g26 ( .A1(n_22), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_1), .B1(n_3), .B2(n_5), .Y(n_27) );
BUFx6f_ASAP7_75t_L g28 ( .A(n_21), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_21), .B(n_5), .Y(n_29) );
INVx2_ASAP7_75t_SL g30 ( .A(n_28), .Y(n_30) );
CKINVDCx6p67_ASAP7_75t_R g31 ( .A(n_29), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_24), .Y(n_33) );
INVx2_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
AND2x2_ASAP7_75t_L g35 ( .A(n_33), .B(n_31), .Y(n_35) );
NAND2xp5_ASAP7_75t_L g36 ( .A(n_35), .B(n_31), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_34), .B(n_27), .Y(n_38) );
AOI221xp5_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_26), .B1(n_24), .B2(n_18), .C(n_17), .Y(n_39) );
AOI322xp5_ASAP7_75t_L g40 ( .A1(n_36), .A2(n_23), .A3(n_20), .B1(n_22), .B2(n_25), .C1(n_24), .C2(n_18), .Y(n_40) );
AOI22xp5_ASAP7_75t_L g41 ( .A1(n_37), .A2(n_19), .B1(n_23), .B2(n_24), .Y(n_41) );
OAI221xp5_ASAP7_75t_L g42 ( .A1(n_39), .A2(n_28), .B1(n_30), .B2(n_9), .C(n_6), .Y(n_42) );
INVx2_ASAP7_75t_SL g43 ( .A(n_40), .Y(n_43) );
INVxp67_ASAP7_75t_L g44 ( .A(n_41), .Y(n_44) );
BUFx2_ASAP7_75t_L g45 ( .A(n_44), .Y(n_45) );
AOI222xp33_ASAP7_75t_L g46 ( .A1(n_43), .A2(n_28), .B1(n_7), .B2(n_30), .C1(n_15), .C2(n_16), .Y(n_46) );
INVx1_ASAP7_75t_L g47 ( .A(n_42), .Y(n_47) );
INVx2_ASAP7_75t_L g48 ( .A(n_42), .Y(n_48) );
HB1xp67_ASAP7_75t_L g49 ( .A(n_45), .Y(n_49) );
AOI22xp5_ASAP7_75t_SL g50 ( .A1(n_49), .A2(n_48), .B1(n_47), .B2(n_46), .Y(n_50) );
endmodule