module real_jpeg_933_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_244;
wire n_128;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_1),
.A2(n_39),
.B1(n_60),
.B2(n_61),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_3),
.A2(n_55),
.B1(n_57),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_68),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_68),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_68),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_27),
.B1(n_29),
.B2(n_49),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_5),
.B(n_69),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_5),
.B(n_27),
.C(n_75),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_5),
.B(n_74),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_5),
.B(n_32),
.C(n_35),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_111),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_5),
.B(n_45),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_5),
.B(n_40),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_5),
.A2(n_60),
.B1(n_61),
.B2(n_111),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_7),
.A2(n_60),
.B1(n_61),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_7),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_7),
.A2(n_55),
.B1(n_57),
.B2(n_79),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_79),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_79),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_12),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_54),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_54),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_26),
.B1(n_60),
.B2(n_61),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_14),
.A2(n_26),
.B1(n_35),
.B2(n_36),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_15),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_140),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_116),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_21),
.B(n_116),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_84),
.C(n_93),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_22),
.B(n_84),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_50),
.B1(n_82),
.B2(n_83),
.Y(n_22)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_24),
.B(n_41),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_38),
.B2(n_40),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_25),
.Y(n_176)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_27),
.A2(n_29),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_27),
.B(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_30),
.A2(n_38),
.B1(n_40),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_30),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_30),
.A2(n_155),
.B(n_157),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_30),
.B(n_159),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_34),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_34),
.A2(n_176),
.B(n_177),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_34),
.A2(n_177),
.B(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_34),
.A2(n_132),
.B1(n_156),
.B2(n_197),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_35),
.B(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_40),
.B(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_42),
.A2(n_45),
.B(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_42),
.A2(n_111),
.B(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_43),
.A2(n_44),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_43),
.A2(n_44),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_43),
.A2(n_44),
.B1(n_114),
.B2(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_43),
.B(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_43),
.A2(n_189),
.B(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_43),
.A2(n_44),
.B1(n_189),
.B2(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_44),
.A2(n_153),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_44),
.B(n_167),
.Y(n_191)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_45),
.A2(n_166),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_70),
.B2(n_71),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_52),
.B(n_70),
.C(n_82),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_58),
.B1(n_67),
.B2(n_69),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_66)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_55),
.A2(n_61),
.A3(n_63),
.B1(n_109),
.B2(n_112),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_111),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_55),
.A2(n_110),
.B(n_111),
.C(n_126),
.Y(n_172)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_66),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_59),
.B(n_100),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_61),
.B1(n_75),
.B2(n_76),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g112 ( 
.A(n_60),
.B(n_64),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_60),
.B(n_163),
.Y(n_162)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B(n_77),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_72),
.A2(n_73),
.B1(n_104),
.B2(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_73),
.A2(n_77),
.B(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_73),
.A2(n_103),
.B1(n_104),
.B2(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_74),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_78),
.Y(n_105)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_92),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_93),
.A2(n_94),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.C(n_106),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_244)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B(n_105),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_104),
.A2(n_105),
.B(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_106),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_113),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_113),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_139),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_130),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_129),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_127),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_128),
.B(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_131),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_132),
.A2(n_158),
.B(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_135),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_240),
.B(n_254),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_183),
.B(n_239),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_168),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_144),
.B(n_168),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_154),
.C(n_160),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_145),
.B(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_149),
.C(n_152),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_154),
.B(n_160),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_161),
.A2(n_162),
.B1(n_164),
.B2(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_179),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_169),
.B(n_180),
.C(n_182),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_178),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_170),
.B(n_174),
.C(n_175),
.Y(n_247)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_234),
.B(n_238),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_224),
.B(n_233),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_206),
.B(n_223),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_200),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_200),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_192),
.B1(n_198),
.B2(n_199),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_195),
.C(n_198),
.Y(n_225)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_217),
.B(n_222),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_212),
.B(n_216),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_215),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_214),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_220),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_226),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_230),
.C(n_231),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_237),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_249),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_248),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_248),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_246),
.C(n_247),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_253),
.Y(n_256)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);


endmodule