module fake_jpeg_4697_n_174 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_28),
.B(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_23),
.B1(n_24),
.B2(n_14),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_34),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_53),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_46),
.B1(n_15),
.B2(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_48),
.B(n_27),
.Y(n_65)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_19),
.B1(n_24),
.B2(n_15),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_50),
.Y(n_62)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_18),
.B1(n_19),
.B2(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_53),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_65),
.B1(n_68),
.B2(n_21),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_35),
.B1(n_37),
.B2(n_34),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_66),
.B1(n_16),
.B2(n_44),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_34),
.B1(n_37),
.B2(n_27),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_52),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_35),
.B1(n_22),
.B2(n_26),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_26),
.B(n_22),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_68),
.B(n_21),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_70),
.B(n_71),
.Y(n_100)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_43),
.B1(n_29),
.B2(n_50),
.Y(n_72)
);

AOI21x1_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_43),
.B(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_81),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_16),
.B(n_32),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_49),
.C(n_45),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_58),
.C(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_56),
.B1(n_63),
.B2(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_82),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_32),
.Y(n_80)
);

A2O1A1O1Ixp25_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_32),
.B(n_49),
.C(n_43),
.D(n_52),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_49),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_88),
.C(n_75),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_65),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_66),
.B1(n_62),
.B2(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_93),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_94),
.B(n_95),
.Y(n_115)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_32),
.B(n_49),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_79),
.B(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_60),
.Y(n_106)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_56),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_74),
.B(n_82),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_108),
.B(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_71),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_112),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_76),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_78),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_89),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_74),
.B(n_73),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_69),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_85),
.C(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_85),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_125),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_97),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_103),
.CI(n_100),
.CON(n_134),
.SN(n_134)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_4),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_99),
.B1(n_93),
.B2(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_114),
.B1(n_92),
.B2(n_101),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_136),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_99),
.B(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_137),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_95),
.B1(n_2),
.B2(n_3),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_12),
.Y(n_136)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_1),
.B(n_2),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_118),
.B(n_124),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_140),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_117),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_131),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_150),
.B(n_118),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_123),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_138),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_155),
.C(n_143),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_145),
.A2(n_133),
.B1(n_121),
.B2(n_132),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_127),
.B(n_134),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_144),
.B1(n_142),
.B2(n_137),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_156),
.B1(n_157),
.B2(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_160),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_155),
.B(n_137),
.C(n_126),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_143),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_135),
.Y(n_166)
);

OAI21x1_ASAP7_75t_SL g169 ( 
.A1(n_164),
.A2(n_157),
.B(n_116),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_167),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_170),
.B(n_8),
.Y(n_172)
);

NOR4xp25_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_163),
.C(n_12),
.D(n_7),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_166),
.A3(n_5),
.B1(n_8),
.B2(n_10),
.C1(n_11),
.C2(n_4),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_SL g173 ( 
.A(n_171),
.B(n_172),
.C(n_10),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_10),
.Y(n_174)
);


endmodule