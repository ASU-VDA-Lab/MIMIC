module fake_jpeg_12878_n_565 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_565);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_565;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_10),
.B(n_14),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_54),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_60),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_59),
.B(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_17),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_62),
.A2(n_103),
.B(n_108),
.Y(n_127)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_65),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_32),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_67),
.B(n_76),
.Y(n_133)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_71),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_72),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_37),
.B(n_1),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_2),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_78),
.B(n_81),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_87),
.Y(n_134)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_32),
.B(n_3),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_40),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_91),
.Y(n_124)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_92),
.Y(n_174)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_93),
.Y(n_169)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_19),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_98),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_37),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_36),
.B(n_3),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_23),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_49),
.Y(n_151)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_23),
.B(n_4),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_63),
.A2(n_109),
.B1(n_64),
.B2(n_70),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_126),
.A2(n_29),
.B1(n_24),
.B2(n_104),
.Y(n_205)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_132),
.Y(n_208)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_140),
.B(n_151),
.Y(n_200)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_62),
.B(n_29),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_143),
.A2(n_41),
.B(n_51),
.Y(n_196)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_149),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_78),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_155),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_62),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_57),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_163),
.Y(n_214)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_60),
.B(n_36),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_165),
.B(n_171),
.Y(n_203)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_65),
.B(n_41),
.Y(n_171)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_55),
.Y(n_173)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_54),
.Y(n_175)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_65),
.Y(n_224)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_179),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_180),
.B(n_183),
.Y(n_258)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_181),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_127),
.A2(n_69),
.B1(n_101),
.B2(n_100),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_182),
.A2(n_198),
.B1(n_205),
.B2(n_228),
.Y(n_294)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_45),
.C(n_44),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_131),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_184),
.B(n_204),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_112),
.A2(n_86),
.B1(n_75),
.B2(n_73),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_188),
.A2(n_240),
.B1(n_160),
.B2(n_159),
.Y(n_254)
);

CKINVDCx9p33_ASAP7_75t_R g189 ( 
.A(n_172),
.Y(n_189)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_189),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_43),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_190),
.B(n_206),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_123),
.A2(n_96),
.B1(n_88),
.B2(n_24),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_191),
.Y(n_296)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_56),
.B1(n_66),
.B2(n_71),
.Y(n_192)
);

AO22x2_ASAP7_75t_L g293 ( 
.A1(n_192),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_293)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_193),
.Y(n_284)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

INVx11_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_196),
.B(n_228),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_126),
.A2(n_77),
.B1(n_72),
.B2(n_26),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_121),
.B(n_129),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_201),
.B(n_135),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_202),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_134),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_130),
.B(n_45),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_141),
.B(n_44),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_213),
.Y(n_245)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_111),
.Y(n_209)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_113),
.Y(n_210)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_210),
.Y(n_292)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_117),
.B(n_118),
.Y(n_213)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_115),
.Y(n_216)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_217),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g218 ( 
.A1(n_153),
.A2(n_93),
.B1(n_91),
.B2(n_53),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_218),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_267)
);

CKINVDCx12_ASAP7_75t_R g219 ( 
.A(n_146),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_221),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_153),
.A2(n_26),
.B1(n_34),
.B2(n_49),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_119),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_110),
.A2(n_26),
.B1(n_52),
.B2(n_51),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_110),
.A2(n_49),
.B1(n_52),
.B2(n_43),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_224),
.B(n_235),
.Y(n_275)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_142),
.Y(n_226)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_137),
.B(n_35),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_227),
.B(n_230),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_49),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_152),
.A2(n_35),
.B1(n_92),
.B2(n_48),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_229),
.A2(n_169),
.B1(n_124),
.B2(n_174),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_132),
.B(n_4),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_142),
.Y(n_231)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_231),
.Y(n_276)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_128),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_232),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_128),
.B(n_4),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_233),
.B(n_189),
.Y(n_290)
);

CKINVDCx12_ASAP7_75t_R g235 ( 
.A(n_124),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_114),
.B(n_122),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_201),
.Y(n_269)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_147),
.Y(n_237)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_144),
.Y(n_238)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_238),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_152),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_116),
.Y(n_241)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_125),
.B1(n_166),
.B2(n_120),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_247),
.A2(n_192),
.B1(n_179),
.B2(n_228),
.Y(n_301)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_178),
.Y(n_251)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_190),
.B(n_138),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_253),
.B(n_269),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_254),
.A2(n_272),
.B1(n_238),
.B2(n_226),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_220),
.A2(n_136),
.B1(n_169),
.B2(n_174),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_255),
.Y(n_343)
);

BUFx24_ASAP7_75t_SL g257 ( 
.A(n_203),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_257),
.B(n_282),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_262),
.Y(n_316)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_263),
.Y(n_300)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_212),
.A2(n_150),
.B(n_6),
.C(n_8),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_278),
.Y(n_302)
);

OAI22x1_ASAP7_75t_L g270 ( 
.A1(n_191),
.A2(n_168),
.B1(n_164),
.B2(n_162),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_270),
.A2(n_194),
.B1(n_215),
.B2(n_217),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_200),
.A2(n_160),
.B1(n_159),
.B2(n_162),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_218),
.A2(n_192),
.B1(n_213),
.B2(n_207),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_274),
.A2(n_294),
.B1(n_192),
.B2(n_229),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_206),
.B(n_168),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_280),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_164),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_9),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_234),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_12),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_225),
.B(n_144),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_288),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_208),
.B(n_135),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_297),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_11),
.Y(n_333)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_211),
.Y(n_295)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_295),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_209),
.B(n_8),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_274),
.B(n_283),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_299),
.A2(n_312),
.B(n_339),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_301),
.A2(n_307),
.B1(n_314),
.B2(n_318),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_248),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_303),
.B(n_338),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_306),
.A2(n_319),
.B1(n_331),
.B2(n_341),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_193),
.B1(n_231),
.B2(n_210),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_327),
.Y(n_356)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_283),
.A2(n_185),
.B(n_199),
.Y(n_312)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_277),
.Y(n_317)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_247),
.A2(n_185),
.B1(n_232),
.B2(n_199),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_245),
.A2(n_194),
.B1(n_197),
.B2(n_187),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_248),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_321),
.Y(n_351)
);

MAJx2_ASAP7_75t_L g322 ( 
.A(n_269),
.B(n_197),
.C(n_187),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g384 ( 
.A(n_322),
.B(n_276),
.C(n_289),
.Y(n_384)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_277),
.Y(n_323)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_286),
.B(n_208),
.C(n_195),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_278),
.C(n_270),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_265),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_325),
.B(n_332),
.Y(n_385)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_326),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_245),
.A2(n_216),
.B1(n_202),
.B2(n_181),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_340),
.Y(n_360)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_267),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_249),
.Y(n_332)
);

AO21x1_ASAP7_75t_L g371 ( 
.A1(n_333),
.A2(n_291),
.B(n_276),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_334),
.Y(n_379)
);

INVx8_ASAP7_75t_L g335 ( 
.A(n_260),
.Y(n_335)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_335),
.Y(n_353)
);

INVx4_ASAP7_75t_SL g336 ( 
.A(n_260),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_336),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_242),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_264),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_283),
.A2(n_12),
.B(n_13),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_244),
.B(n_12),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_267),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_341)
);

FAx1_ASAP7_75t_SL g342 ( 
.A(n_244),
.B(n_15),
.CI(n_16),
.CON(n_342),
.SN(n_342)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_344),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_258),
.B(n_15),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_275),
.B(n_15),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_289),
.Y(n_367)
);

XNOR2x1_ASAP7_75t_L g407 ( 
.A(n_346),
.B(n_384),
.Y(n_407)
);

OAI32xp33_ASAP7_75t_L g349 ( 
.A1(n_302),
.A2(n_268),
.A3(n_293),
.B1(n_295),
.B2(n_279),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_363),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_271),
.C(n_252),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_350),
.B(n_352),
.C(n_357),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_250),
.C(n_285),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_264),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_306),
.A2(n_293),
.B1(n_279),
.B2(n_242),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_359),
.A2(n_362),
.B1(n_348),
.B2(n_371),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_330),
.A2(n_302),
.B1(n_331),
.B2(n_341),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_293),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_321),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_367),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_320),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_328),
.B(n_250),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_369),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_285),
.Y(n_369)
);

O2A1O1Ixp33_ASAP7_75t_L g370 ( 
.A1(n_299),
.A2(n_246),
.B(n_261),
.C(n_256),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_370),
.B(n_336),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_371),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_273),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_378),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g375 ( 
.A1(n_333),
.A2(n_246),
.B(n_261),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_375),
.A2(n_343),
.B(n_309),
.Y(n_388)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_334),
.Y(n_377)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_377),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_305),
.B(n_273),
.Y(n_378)
);

NOR2x1_ASAP7_75t_R g380 ( 
.A(n_342),
.B(n_312),
.Y(n_380)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_384),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_327),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_386),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_342),
.B(n_303),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_383),
.B(n_339),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_319),
.Y(n_386)
);

INVx13_ASAP7_75t_L g387 ( 
.A(n_351),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_387),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_388),
.A2(n_353),
.B(n_374),
.Y(n_442)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_381),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

INVx13_ASAP7_75t_L g390 ( 
.A(n_381),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_390),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_347),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_391),
.B(n_392),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_385),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_359),
.A2(n_307),
.B1(n_343),
.B2(n_309),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_393),
.A2(n_403),
.B1(n_421),
.B2(n_375),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_395),
.B(n_414),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_378),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_396),
.B(n_419),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_397),
.B(n_422),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_383),
.A2(n_333),
.B(n_311),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_398),
.A2(n_401),
.B(n_369),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_358),
.A2(n_338),
.B(n_332),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_348),
.A2(n_308),
.B1(n_313),
.B2(n_300),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_356),
.A2(n_335),
.B1(n_316),
.B2(n_310),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_406),
.A2(n_417),
.B1(n_353),
.B2(n_379),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_350),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_411),
.C(n_412),
.Y(n_430)
);

MAJx2_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_313),
.C(n_304),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_352),
.B(n_320),
.C(n_300),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_413),
.A2(n_416),
.B(n_394),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_298),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_357),
.B(n_298),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_420),
.C(n_355),
.Y(n_440)
);

AND2x6_ASAP7_75t_L g416 ( 
.A(n_370),
.B(n_336),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_386),
.A2(n_316),
.B1(n_326),
.B2(n_323),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_363),
.B(n_317),
.Y(n_418)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_418),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_376),
.B(n_256),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_376),
.B(n_315),
.C(n_284),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_402),
.A2(n_362),
.B1(n_372),
.B2(n_346),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_423),
.A2(n_393),
.B1(n_403),
.B2(n_392),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_424),
.A2(n_439),
.B1(n_425),
.B2(n_432),
.Y(n_477)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_400),
.Y(n_426)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_426),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_427),
.A2(n_402),
.B(n_401),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_358),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_428),
.B(n_437),
.Y(n_460)
);

NOR3xp33_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_454),
.C(n_398),
.Y(n_466)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_404),
.Y(n_431)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_431),
.Y(n_465)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_405),
.Y(n_432)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_433),
.B(n_379),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_397),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_407),
.B(n_360),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_395),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_421),
.A2(n_375),
.B1(n_356),
.B2(n_349),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_444),
.C(n_447),
.Y(n_457)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_441),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_442),
.A2(n_413),
.B(n_388),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_399),
.B(n_360),
.C(n_368),
.Y(n_444)
);

AO22x1_ASAP7_75t_SL g445 ( 
.A1(n_394),
.A2(n_380),
.B1(n_355),
.B2(n_354),
.Y(n_445)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_445),
.Y(n_469)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_417),
.Y(n_446)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_446),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_407),
.B(n_354),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_418),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_448),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_391),
.B(n_315),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_452),
.B(n_453),
.Y(n_461)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_410),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_410),
.Y(n_454)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_449),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_456),
.B(n_466),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_412),
.C(n_415),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_459),
.C(n_468),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_428),
.C(n_447),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_462),
.A2(n_427),
.B(n_445),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_463),
.A2(n_471),
.B(n_387),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_411),
.C(n_422),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_449),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_481),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_442),
.A2(n_413),
.B(n_416),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_474),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_420),
.C(n_396),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_480),
.C(n_458),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_475),
.A2(n_477),
.B1(n_450),
.B2(n_423),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_443),
.Y(n_478)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_478),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_444),
.B(n_374),
.C(n_390),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_443),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_SL g483 ( 
.A(n_459),
.B(n_434),
.C(n_436),
.Y(n_483)
);

AOI21xp33_ASAP7_75t_L g504 ( 
.A1(n_483),
.A2(n_468),
.B(n_475),
.Y(n_504)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_478),
.Y(n_486)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_486),
.Y(n_509)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_465),
.Y(n_487)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_487),
.Y(n_512)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_464),
.Y(n_488)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_488),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_493),
.C(n_497),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_491),
.A2(n_495),
.B1(n_501),
.B2(n_456),
.Y(n_505)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_461),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_SL g518 ( 
.A1(n_492),
.A2(n_476),
.B1(n_474),
.B2(n_463),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_438),
.C(n_435),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_479),
.A2(n_441),
.B1(n_429),
.B2(n_424),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_496),
.B(n_500),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_457),
.B(n_435),
.C(n_451),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_445),
.C(n_439),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_502),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_499),
.A2(n_471),
.B(n_476),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_473),
.B(n_390),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_479),
.A2(n_408),
.B1(n_377),
.B2(n_389),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_460),
.B(n_389),
.C(n_408),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_460),
.B(n_361),
.C(n_387),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_462),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_504),
.B(n_497),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_505),
.A2(n_516),
.B1(n_509),
.B2(n_502),
.Y(n_523)
);

CKINVDCx14_ASAP7_75t_R g507 ( 
.A(n_482),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_514),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_485),
.A2(n_469),
.B1(n_455),
.B2(n_467),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_508),
.A2(n_516),
.B1(n_518),
.B2(n_292),
.Y(n_536)
);

INVx13_ASAP7_75t_L g513 ( 
.A(n_501),
.Y(n_513)
);

INVx11_ASAP7_75t_L g528 ( 
.A(n_513),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_494),
.B(n_467),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_495),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_498),
.A2(n_469),
.B1(n_475),
.B2(n_455),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_517),
.B(n_519),
.Y(n_531)
);

INVx13_ASAP7_75t_L g519 ( 
.A(n_496),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_520),
.B(n_521),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_522),
.B(n_527),
.Y(n_539)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_523),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_519),
.A2(n_491),
.B(n_503),
.Y(n_524)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_524),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_517),
.A2(n_493),
.B(n_490),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_526),
.B(n_510),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_507),
.B(n_500),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_506),
.B(n_489),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_529),
.B(n_530),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_514),
.B(n_490),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_505),
.A2(n_484),
.B1(n_472),
.B2(n_334),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_532),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_511),
.B(n_484),
.C(n_361),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_534),
.B(n_535),
.C(n_512),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_511),
.B(n_292),
.C(n_16),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_536),
.A2(n_509),
.B1(n_512),
.B2(n_515),
.Y(n_540)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_537),
.Y(n_548)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_540),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_532),
.C(n_506),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_541),
.B(n_542),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_525),
.A2(n_515),
.B1(n_513),
.B2(n_519),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_523),
.B(n_510),
.C(n_521),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_544),
.B(n_524),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_547),
.B(n_533),
.Y(n_551)
);

AOI31xp67_ASAP7_75t_L g549 ( 
.A1(n_539),
.A2(n_528),
.A3(n_533),
.B(n_508),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_549),
.A2(n_538),
.B1(n_528),
.B2(n_544),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_550),
.B(n_551),
.Y(n_554)
);

NOR2x1_ASAP7_75t_L g555 ( 
.A(n_548),
.B(n_525),
.Y(n_555)
);

NOR2x1_ASAP7_75t_L g559 ( 
.A(n_555),
.B(n_553),
.Y(n_559)
);

NOR2xp67_ASAP7_75t_L g556 ( 
.A(n_552),
.B(n_546),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_556),
.A2(n_557),
.B(n_554),
.Y(n_558)
);

AOI322xp5_ASAP7_75t_L g560 ( 
.A1(n_558),
.A2(n_559),
.A3(n_543),
.B1(n_549),
.B2(n_520),
.C1(n_513),
.C2(n_541),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_537),
.C(n_531),
.Y(n_561)
);

OA21x2_ASAP7_75t_SL g562 ( 
.A1(n_561),
.A2(n_545),
.B(n_547),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_SL g563 ( 
.A(n_562),
.B(n_531),
.C(n_526),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_563),
.B(n_535),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_564),
.B(n_17),
.C(n_554),
.Y(n_565)
);


endmodule