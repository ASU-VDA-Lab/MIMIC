module real_jpeg_32398_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_10;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_0),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_0),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_1),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_1),
.A2(n_17),
.B1(n_86),
.B2(n_88),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_1),
.A2(n_17),
.B1(n_138),
.B2(n_142),
.Y(n_137)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_2),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_3),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_4),
.B(n_62),
.Y(n_61)
);

AO22x1_ASAP7_75t_SL g79 ( 
.A1(n_4),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_4),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_4),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_4),
.A2(n_83),
.B1(n_150),
.B2(n_153),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_4),
.A2(n_173),
.A3(n_176),
.B1(n_178),
.B2(n_183),
.Y(n_172)
);

OAI22x1_ASAP7_75t_SL g190 ( 
.A1(n_4),
.A2(n_83),
.B1(n_191),
.B2(n_194),
.Y(n_190)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_7),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_8),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_8),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_8),
.A2(n_55),
.B1(n_212),
.B2(n_215),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_167),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_166),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp67_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_100),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_13),
.B(n_100),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_60),
.C(n_72),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_14),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_48),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_25),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_16),
.B(n_49),
.Y(n_133)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_19),
.A2(n_64),
.B1(n_66),
.B2(n_71),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_20),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_25),
.B(n_50),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_25),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_R g221 ( 
.A(n_37),
.B(n_83),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_40),
.Y(n_186)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_43),
.Y(n_231)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_47),
.Y(n_182)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_47),
.Y(n_217)
);

NAND2x1_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_51),
.B(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_54),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_59),
.Y(n_193)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_62),
.B(n_137),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AO21x2_ASAP7_75t_L g157 ( 
.A1(n_63),
.A2(n_112),
.B(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_73),
.B(n_200),
.Y(n_199)
);

AND2x4_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_84),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_79),
.B(n_92),
.Y(n_228)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_104),
.A3(n_107),
.B1(n_111),
.B2(n_119),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_83),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_83),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_84),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_85),
.B(n_206),
.Y(n_205)
);

BUFx4f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_92),
.B(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21x1_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_125),
.B(n_129),
.Y(n_124)
);

NAND2x1_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_130),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_123),
.B2(n_124),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_165),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_146),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_157),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_202),
.B(n_236),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_199),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_170),
.B(n_199),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_187),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_171),
.A2(n_172),
.B1(n_187),
.B2(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx2_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_219),
.B(n_235),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_218),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_218),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_227),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_SL g233 ( 
.A(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_225),
.B(n_234),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_222),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);


endmodule