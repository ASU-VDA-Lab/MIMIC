module fake_jpeg_3385_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx11_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_9),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_22),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_20),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_29),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_35),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_17),
.B1(n_16),
.B2(n_18),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_25),
.B1(n_10),
.B2(n_11),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_28),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_18),
.B1(n_25),
.B2(n_9),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_27),
.B(n_26),
.Y(n_37)
);

A2O1A1O1Ixp25_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_10),
.B(n_11),
.C(n_13),
.D(n_6),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_45),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_47),
.B(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_49),
.B(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_51),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_46),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_54)
);


endmodule