module real_aes_7373_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_87), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g447 ( .A(n_0), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_1), .Y(n_748) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_2), .A2(n_141), .B(n_144), .C(n_219), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_3), .A2(n_169), .B(n_170), .Y(n_168) );
INVx1_ASAP7_75t_L g498 ( .A(n_4), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_5), .B(n_180), .Y(n_179) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_6), .A2(n_169), .B(n_476), .Y(n_475) );
AND2x6_ASAP7_75t_L g141 ( .A(n_7), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g244 ( .A(n_8), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_9), .B(n_42), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_10), .A2(n_268), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_11), .B(n_153), .Y(n_221) );
INVx1_ASAP7_75t_L g480 ( .A(n_12), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_13), .B(n_174), .Y(n_531) );
INVx1_ASAP7_75t_L g133 ( .A(n_14), .Y(n_133) );
INVx1_ASAP7_75t_L g543 ( .A(n_15), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_16), .A2(n_188), .B(n_229), .C(n_231), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_17), .B(n_180), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_18), .B(n_469), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_19), .A2(n_102), .B1(n_111), .B2(n_751), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_20), .B(n_169), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_21), .B(n_276), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_22), .A2(n_174), .B(n_205), .C(n_208), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_23), .B(n_180), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_24), .B(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_25), .A2(n_207), .B(n_231), .C(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_26), .B(n_153), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g135 ( .A(n_27), .Y(n_135) );
INVx1_ASAP7_75t_L g186 ( .A(n_28), .Y(n_186) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_29), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_30), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_31), .B(n_153), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_32), .Y(n_449) );
INVx1_ASAP7_75t_L g273 ( .A(n_33), .Y(n_273) );
INVx1_ASAP7_75t_L g488 ( .A(n_34), .Y(n_488) );
INVx2_ASAP7_75t_L g139 ( .A(n_35), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_36), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_37), .A2(n_174), .B(n_175), .C(n_177), .Y(n_173) );
INVxp67_ASAP7_75t_L g274 ( .A(n_38), .Y(n_274) );
CKINVDCx14_ASAP7_75t_R g171 ( .A(n_39), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_40), .A2(n_144), .B(n_185), .C(n_192), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_41), .A2(n_141), .B(n_144), .C(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g487 ( .A(n_43), .Y(n_487) );
OAI22xp5_ASAP7_75t_SL g440 ( .A1(n_44), .A2(n_50), .B1(n_441), .B2(n_442), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_44), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_45), .A2(n_63), .B1(n_741), .B2(n_742), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_45), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_46), .A2(n_155), .B(n_242), .C(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_47), .B(n_153), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_48), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_49), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_50), .Y(n_441) );
INVx1_ASAP7_75t_L g203 ( .A(n_51), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_52), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_53), .B(n_169), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_54), .A2(n_144), .B1(n_208), .B2(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_55), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_56), .Y(n_495) );
CKINVDCx14_ASAP7_75t_R g240 ( .A(n_57), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_58), .A2(n_177), .B(n_242), .C(n_479), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_59), .Y(n_523) );
INVx1_ASAP7_75t_L g477 ( .A(n_60), .Y(n_477) );
INVx1_ASAP7_75t_L g142 ( .A(n_61), .Y(n_142) );
INVx1_ASAP7_75t_L g132 ( .A(n_62), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_63), .Y(n_741) );
INVx1_ASAP7_75t_SL g176 ( .A(n_64), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_65), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_66), .B(n_180), .Y(n_210) );
INVx1_ASAP7_75t_L g148 ( .A(n_67), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_SL g468 ( .A1(n_68), .A2(n_177), .B(n_469), .C(n_470), .Y(n_468) );
INVxp67_ASAP7_75t_L g471 ( .A(n_69), .Y(n_471) );
INVx1_ASAP7_75t_L g110 ( .A(n_70), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_71), .A2(n_169), .B(n_239), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_72), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_73), .A2(n_169), .B(n_226), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_74), .Y(n_491) );
INVx1_ASAP7_75t_L g517 ( .A(n_75), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_76), .A2(n_268), .B(n_269), .Y(n_267) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_77), .Y(n_183) );
INVx1_ASAP7_75t_L g227 ( .A(n_78), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_79), .A2(n_141), .B(n_144), .C(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_80), .A2(n_169), .B(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g230 ( .A(n_81), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_82), .B(n_187), .Y(n_511) );
INVx2_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
INVx1_ASAP7_75t_L g220 ( .A(n_84), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_85), .B(n_469), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_86), .A2(n_141), .B(n_144), .C(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g444 ( .A(n_87), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g455 ( .A(n_87), .Y(n_455) );
OR2x2_ASAP7_75t_L g738 ( .A(n_87), .B(n_446), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_88), .A2(n_144), .B(n_147), .C(n_157), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_89), .B(n_162), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_90), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_91), .A2(n_141), .B(n_144), .C(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_92), .Y(n_535) );
INVx1_ASAP7_75t_L g467 ( .A(n_93), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_94), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_95), .B(n_187), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_96), .B(n_128), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_97), .B(n_128), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g206 ( .A(n_99), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_100), .A2(n_169), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx12_ASAP7_75t_R g753 ( .A(n_104), .Y(n_753) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g446 ( .A(n_105), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_117), .B(n_450), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g750 ( .A(n_115), .Y(n_750) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_443), .B(n_448), .Y(n_117) );
XNOR2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_440), .Y(n_118) );
INVx3_ASAP7_75t_L g739 ( .A(n_119), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_119), .A2(n_453), .B1(n_737), .B2(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_SL g119 ( .A(n_120), .B(n_395), .Y(n_119) );
NOR4xp25_ASAP7_75t_L g120 ( .A(n_121), .B(n_332), .C(n_366), .D(n_382), .Y(n_120) );
NAND4xp25_ASAP7_75t_SL g121 ( .A(n_122), .B(n_258), .C(n_296), .D(n_312), .Y(n_121) );
AOI222xp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_195), .B1(n_233), .B2(n_246), .C1(n_251), .C2(n_257), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI31xp33_ASAP7_75t_L g428 ( .A1(n_124), .A2(n_429), .A3(n_430), .B(n_432), .Y(n_428) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_163), .Y(n_124) );
AND2x2_ASAP7_75t_L g403 ( .A(n_125), .B(n_165), .Y(n_403) );
BUFx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_SL g250 ( .A(n_126), .Y(n_250) );
AND2x2_ASAP7_75t_L g257 ( .A(n_126), .B(n_181), .Y(n_257) );
AND2x2_ASAP7_75t_L g317 ( .A(n_126), .B(n_166), .Y(n_317) );
AO21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_134), .B(n_159), .Y(n_126) );
INVx3_ASAP7_75t_L g180 ( .A(n_127), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_127), .B(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_127), .B(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_SL g513 ( .A(n_127), .B(n_514), .Y(n_513) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_128), .A2(n_465), .B(n_472), .Y(n_464) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g266 ( .A(n_129), .Y(n_266) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g162 ( .A(n_130), .B(n_131), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_143), .Y(n_134) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_136), .A2(n_162), .B(n_183), .C(n_184), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_136), .A2(n_217), .B(n_218), .Y(n_216) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_136), .A2(n_158), .B1(n_485), .B2(n_489), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_136), .A2(n_495), .B(n_496), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_136), .A2(n_517), .B(n_518), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
AND2x4_ASAP7_75t_L g169 ( .A(n_137), .B(n_141), .Y(n_169) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g191 ( .A(n_138), .Y(n_191) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
INVx1_ASAP7_75t_L g209 ( .A(n_139), .Y(n_209) );
INVx1_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_140), .Y(n_153) );
INVx3_ASAP7_75t_L g188 ( .A(n_140), .Y(n_188) );
INVx1_ASAP7_75t_L g469 ( .A(n_140), .Y(n_469) );
INVx4_ASAP7_75t_SL g158 ( .A(n_141), .Y(n_158) );
BUFx3_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
INVx5_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx3_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_145), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_152), .C(n_154), .Y(n_147) );
O2A1O1Ixp5_ASAP7_75t_L g219 ( .A1(n_149), .A2(n_154), .B(n_220), .C(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g486 ( .A1(n_150), .A2(n_151), .B1(n_487), .B2(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx4_ASAP7_75t_L g207 ( .A(n_151), .Y(n_207) );
INVx4_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
INVx2_ASAP7_75t_L g242 ( .A(n_153), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_154), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_154), .A2(n_520), .B(n_521), .Y(n_519) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g231 ( .A(n_156), .Y(n_231) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g170 ( .A1(n_158), .A2(n_171), .B(n_172), .C(n_173), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_SL g202 ( .A1(n_158), .A2(n_172), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_SL g226 ( .A1(n_158), .A2(n_172), .B(n_227), .C(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_SL g239 ( .A1(n_158), .A2(n_172), .B(n_240), .C(n_241), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g269 ( .A1(n_158), .A2(n_172), .B(n_270), .C(n_271), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_158), .A2(n_172), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_158), .A2(n_172), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_158), .A2(n_172), .B(n_540), .C(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx1_ASAP7_75t_L g276 ( .A(n_161), .Y(n_276) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_161), .A2(n_527), .B(n_534), .Y(n_526) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_162), .A2(n_238), .B(n_245), .Y(n_237) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_162), .A2(n_538), .B(n_544), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_163), .B(n_347), .Y(n_346) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_164), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_164), .B(n_261), .Y(n_307) );
AND2x2_ASAP7_75t_L g400 ( .A(n_164), .B(n_340), .Y(n_400) );
OAI321xp33_ASAP7_75t_L g434 ( .A1(n_164), .A2(n_250), .A3(n_407), .B1(n_435), .B2(n_437), .C(n_438), .Y(n_434) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_164), .B(n_236), .C(n_347), .D(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_181), .Y(n_164) );
AND2x2_ASAP7_75t_L g302 ( .A(n_165), .B(n_248), .Y(n_302) );
AND2x2_ASAP7_75t_L g321 ( .A(n_165), .B(n_250), .Y(n_321) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g249 ( .A(n_166), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g277 ( .A(n_166), .B(n_181), .Y(n_277) );
AND2x2_ASAP7_75t_L g363 ( .A(n_166), .B(n_248), .Y(n_363) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_179), .Y(n_166) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_167), .A2(n_201), .B(n_210), .Y(n_200) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_167), .A2(n_225), .B(n_232), .Y(n_224) );
BUFx2_ASAP7_75t_L g268 ( .A(n_169), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_174), .B(n_176), .Y(n_175) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_178), .Y(n_532) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_180), .A2(n_475), .B(n_481), .Y(n_474) );
INVx3_ASAP7_75t_SL g248 ( .A(n_181), .Y(n_248) );
AND2x2_ASAP7_75t_L g295 ( .A(n_181), .B(n_282), .Y(n_295) );
OR2x2_ASAP7_75t_L g328 ( .A(n_181), .B(n_250), .Y(n_328) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_181), .Y(n_335) );
AND2x2_ASAP7_75t_L g364 ( .A(n_181), .B(n_249), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_181), .B(n_337), .Y(n_379) );
AND2x2_ASAP7_75t_L g411 ( .A(n_181), .B(n_403), .Y(n_411) );
AND2x2_ASAP7_75t_L g420 ( .A(n_181), .B(n_262), .Y(n_420) );
OR2x6_ASAP7_75t_L g181 ( .A(n_182), .B(n_193), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_189), .C(n_190), .Y(n_185) );
OAI22xp33_ASAP7_75t_L g272 ( .A1(n_187), .A2(n_207), .B1(n_273), .B2(n_274), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_187), .A2(n_498), .B(n_499), .C(n_500), .Y(n_497) );
INVx5_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_188), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_188), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_188), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_191), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_211), .Y(n_196) );
INVx1_ASAP7_75t_SL g388 ( .A(n_197), .Y(n_388) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g253 ( .A(n_198), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g235 ( .A(n_199), .B(n_213), .Y(n_235) );
AND2x2_ASAP7_75t_L g324 ( .A(n_199), .B(n_237), .Y(n_324) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g294 ( .A(n_200), .B(n_224), .Y(n_294) );
OR2x2_ASAP7_75t_L g305 ( .A(n_200), .B(n_237), .Y(n_305) );
AND2x2_ASAP7_75t_L g331 ( .A(n_200), .B(n_237), .Y(n_331) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_200), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_207), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_207), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g500 ( .A(n_208), .Y(n_500) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_211), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_211), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g304 ( .A(n_212), .B(n_305), .Y(n_304) );
AOI322xp5_ASAP7_75t_L g390 ( .A1(n_212), .A2(n_294), .A3(n_300), .B1(n_331), .B2(n_381), .C1(n_391), .C2(n_393), .Y(n_390) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_224), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_213), .B(n_236), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_213), .B(n_237), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_213), .B(n_254), .Y(n_311) );
AND2x2_ASAP7_75t_L g365 ( .A(n_213), .B(n_331), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_213), .Y(n_369) );
AND2x2_ASAP7_75t_L g381 ( .A(n_213), .B(n_224), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_213), .B(n_253), .Y(n_413) );
INVx4_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g278 ( .A(n_214), .B(n_224), .Y(n_278) );
BUFx3_ASAP7_75t_L g292 ( .A(n_214), .Y(n_292) );
AND3x2_ASAP7_75t_L g374 ( .A(n_214), .B(n_354), .C(n_375), .Y(n_374) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_222), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_215), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_215), .B(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_215), .B(n_535), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g234 ( .A(n_224), .B(n_235), .C(n_236), .Y(n_234) );
INVx1_ASAP7_75t_SL g254 ( .A(n_224), .Y(n_254) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_224), .Y(n_359) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g353 ( .A(n_235), .B(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g360 ( .A(n_235), .Y(n_360) );
AND2x2_ASAP7_75t_L g398 ( .A(n_236), .B(n_376), .Y(n_398) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
BUFx3_ASAP7_75t_L g279 ( .A(n_237), .Y(n_279) );
AND2x2_ASAP7_75t_L g354 ( .A(n_237), .B(n_254), .Y(n_354) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
OR2x2_ASAP7_75t_L g298 ( .A(n_248), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g417 ( .A(n_248), .B(n_317), .Y(n_417) );
AND2x2_ASAP7_75t_L g431 ( .A(n_248), .B(n_250), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_249), .B(n_262), .Y(n_372) );
AND2x2_ASAP7_75t_L g419 ( .A(n_249), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g282 ( .A(n_250), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g299 ( .A(n_250), .B(n_262), .Y(n_299) );
INVx1_ASAP7_75t_L g309 ( .A(n_250), .Y(n_309) );
AND2x2_ASAP7_75t_L g340 ( .A(n_250), .B(n_262), .Y(n_340) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_252), .A2(n_383), .B1(n_387), .B2(n_389), .C(n_390), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_253), .B(n_255), .Y(n_252) );
AND2x2_ASAP7_75t_L g286 ( .A(n_253), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_256), .B(n_293), .Y(n_436) );
AOI322xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_278), .A3(n_279), .B1(n_280), .B2(n_286), .C1(n_288), .C2(n_295), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_277), .Y(n_260) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_261), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_261), .B(n_327), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g350 ( .A1(n_261), .A2(n_277), .B(n_351), .C(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_261), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_261), .B(n_321), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_261), .B(n_403), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_261), .B(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_262), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_262), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g392 ( .A(n_262), .B(n_279), .Y(n_392) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_267), .B(n_275), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_264), .A2(n_284), .B(n_285), .Y(n_283) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_264), .A2(n_516), .B(n_522), .Y(n_515) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AOI21xp5_ASAP7_75t_SL g507 ( .A1(n_265), .A2(n_508), .B(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_266), .A2(n_484), .B(n_490), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_266), .B(n_491), .Y(n_490) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_266), .A2(n_494), .B(n_501), .Y(n_493) );
INVx1_ASAP7_75t_L g284 ( .A(n_267), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_275), .Y(n_285) );
INVx1_ASAP7_75t_L g367 ( .A(n_277), .Y(n_367) );
OAI31xp33_ASAP7_75t_L g377 ( .A1(n_277), .A2(n_302), .A3(n_378), .B(n_380), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_277), .B(n_283), .Y(n_429) );
INVx1_ASAP7_75t_SL g290 ( .A(n_278), .Y(n_290) );
AND2x2_ASAP7_75t_L g323 ( .A(n_278), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g404 ( .A(n_278), .B(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g289 ( .A(n_279), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g314 ( .A(n_279), .Y(n_314) );
AND2x2_ASAP7_75t_L g341 ( .A(n_279), .B(n_294), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_279), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g433 ( .A(n_279), .B(n_381), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_281), .B(n_351), .Y(n_424) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g320 ( .A(n_283), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g338 ( .A(n_283), .Y(n_338) );
NAND2xp33_ASAP7_75t_SL g288 ( .A(n_289), .B(n_291), .Y(n_288) );
OAI211xp5_ASAP7_75t_SL g332 ( .A1(n_290), .A2(n_333), .B(n_339), .C(n_355), .Y(n_332) );
OR2x2_ASAP7_75t_L g407 ( .A(n_290), .B(n_388), .Y(n_407) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_292), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_292), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g313 ( .A(n_294), .B(n_314), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_300), .B(n_303), .C(n_306), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_SL g347 ( .A(n_299), .Y(n_347) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_302), .B(n_340), .Y(n_345) );
INVx1_ASAP7_75t_L g351 ( .A(n_302), .Y(n_351) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g310 ( .A(n_305), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g343 ( .A(n_305), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g405 ( .A(n_305), .Y(n_405) );
AOI21xp33_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_308), .B(n_310), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_308), .A2(n_319), .B(n_322), .Y(n_318) );
AOI211xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_315), .B(n_318), .C(n_325), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_313), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_316), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_SL g329 ( .A(n_317), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_319), .A2(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_324), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g349 ( .A(n_324), .Y(n_349) );
AOI21xp33_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_329), .B(n_330), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g380 ( .A(n_331), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_337), .B(n_363), .Y(n_389) );
AND2x2_ASAP7_75t_L g402 ( .A(n_337), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g416 ( .A(n_337), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g426 ( .A(n_337), .B(n_364), .Y(n_426) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI211xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B(n_342), .C(n_350), .Y(n_339) );
INVx1_ASAP7_75t_L g386 ( .A(n_340), .Y(n_386) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .B1(n_346), .B2(n_348), .Y(n_342) );
OR2x2_ASAP7_75t_L g348 ( .A(n_344), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_344), .B(n_405), .Y(n_427) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g421 ( .A(n_354), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_361), .B1(n_364), .B2(n_365), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g439 ( .A(n_359), .Y(n_439) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g385 ( .A(n_363), .Y(n_385) );
OAI211xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_368), .B(n_370), .C(n_377), .Y(n_366) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_385), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NOR5xp2_ASAP7_75t_L g395 ( .A(n_396), .B(n_414), .C(n_422), .D(n_428), .E(n_434), .Y(n_395) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_397), .A2(n_399), .B(n_401), .C(n_408), .Y(n_396) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B(n_406), .Y(n_401) );
OAI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B(n_412), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_411), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AOI21xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_418), .B(n_421), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g437 ( .A(n_417), .Y(n_437) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2xp33_ASAP7_75t_SL g448 ( .A(n_444), .B(n_449), .Y(n_448) );
NOR2x2_ASAP7_75t_L g747 ( .A(n_445), .B(n_455), .Y(n_747) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g454 ( .A(n_446), .B(n_455), .Y(n_454) );
OAI21xp5_ASAP7_75t_SL g450 ( .A1(n_448), .A2(n_451), .B(n_749), .Y(n_450) );
OAI222xp33_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_740), .B1(n_743), .B2(n_745), .C1(n_746), .C2(n_748), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_456), .B1(n_737), .B2(n_739), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g744 ( .A(n_456), .Y(n_744) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND4x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_655), .C(n_702), .D(n_722), .Y(n_457) );
NOR3xp33_ASAP7_75t_SL g458 ( .A(n_459), .B(n_585), .C(n_610), .Y(n_458) );
OAI211xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_503), .B(n_545), .C(n_575), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_482), .Y(n_461) );
INVx3_ASAP7_75t_SL g627 ( .A(n_462), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_462), .B(n_558), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_462), .B(n_492), .Y(n_708) );
AND2x2_ASAP7_75t_L g731 ( .A(n_462), .B(n_597), .Y(n_731) );
AND2x4_ASAP7_75t_L g462 ( .A(n_463), .B(n_473), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g549 ( .A(n_464), .B(n_474), .Y(n_549) );
INVx3_ASAP7_75t_L g562 ( .A(n_464), .Y(n_562) );
AND2x2_ASAP7_75t_L g567 ( .A(n_464), .B(n_473), .Y(n_567) );
OR2x2_ASAP7_75t_L g618 ( .A(n_464), .B(n_559), .Y(n_618) );
BUFx2_ASAP7_75t_L g638 ( .A(n_464), .Y(n_638) );
AND2x2_ASAP7_75t_L g648 ( .A(n_464), .B(n_559), .Y(n_648) );
AND2x2_ASAP7_75t_L g654 ( .A(n_464), .B(n_483), .Y(n_654) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_474), .B(n_559), .Y(n_573) );
INVx2_ASAP7_75t_L g583 ( .A(n_474), .Y(n_583) );
AND2x2_ASAP7_75t_L g596 ( .A(n_474), .B(n_562), .Y(n_596) );
OR2x2_ASAP7_75t_L g607 ( .A(n_474), .B(n_559), .Y(n_607) );
AND2x2_ASAP7_75t_SL g653 ( .A(n_474), .B(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g665 ( .A(n_474), .Y(n_665) );
AND2x2_ASAP7_75t_L g711 ( .A(n_474), .B(n_483), .Y(n_711) );
INVx3_ASAP7_75t_SL g584 ( .A(n_482), .Y(n_584) );
OR2x2_ASAP7_75t_L g637 ( .A(n_482), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_492), .Y(n_482) );
INVx3_ASAP7_75t_L g559 ( .A(n_483), .Y(n_559) );
AND2x2_ASAP7_75t_L g626 ( .A(n_483), .B(n_493), .Y(n_626) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_483), .Y(n_694) );
AOI33xp33_ASAP7_75t_L g698 ( .A1(n_483), .A2(n_627), .A3(n_634), .B1(n_643), .B2(n_699), .B3(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g547 ( .A(n_492), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_492), .B(n_562), .Y(n_561) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_492), .B(n_622), .C(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_L g647 ( .A(n_492), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_492), .B(n_654), .Y(n_657) );
AND2x2_ASAP7_75t_L g710 ( .A(n_492), .B(n_711), .Y(n_710) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g566 ( .A(n_493), .Y(n_566) );
OR2x2_ASAP7_75t_L g660 ( .A(n_493), .B(n_559), .Y(n_660) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_524), .Y(n_503) );
AOI32xp33_ASAP7_75t_L g611 ( .A1(n_504), .A2(n_612), .A3(n_614), .B1(n_616), .B2(n_619), .Y(n_611) );
NOR2xp67_ASAP7_75t_L g684 ( .A(n_504), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g714 ( .A(n_504), .Y(n_714) );
INVx4_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g646 ( .A(n_505), .B(n_630), .Y(n_646) );
AND2x2_ASAP7_75t_L g666 ( .A(n_505), .B(n_592), .Y(n_666) );
AND2x2_ASAP7_75t_L g734 ( .A(n_505), .B(n_652), .Y(n_734) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
INVx3_ASAP7_75t_L g555 ( .A(n_506), .Y(n_555) );
AND2x2_ASAP7_75t_L g569 ( .A(n_506), .B(n_553), .Y(n_569) );
OR2x2_ASAP7_75t_L g574 ( .A(n_506), .B(n_552), .Y(n_574) );
INVx1_ASAP7_75t_L g581 ( .A(n_506), .Y(n_581) );
AND2x2_ASAP7_75t_L g589 ( .A(n_506), .B(n_563), .Y(n_589) );
AND2x2_ASAP7_75t_L g591 ( .A(n_506), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_506), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g644 ( .A(n_506), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_506), .B(n_729), .Y(n_728) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_513), .Y(n_506) );
INVx2_ASAP7_75t_L g553 ( .A(n_515), .Y(n_553) );
AND2x2_ASAP7_75t_L g599 ( .A(n_515), .B(n_525), .Y(n_599) );
AND2x2_ASAP7_75t_L g609 ( .A(n_515), .B(n_537), .Y(n_609) );
INVx2_ASAP7_75t_L g729 ( .A(n_524), .Y(n_729) );
OR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_536), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_525), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g570 ( .A(n_525), .Y(n_570) );
AND2x2_ASAP7_75t_L g614 ( .A(n_525), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g630 ( .A(n_525), .B(n_593), .Y(n_630) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g578 ( .A(n_526), .Y(n_578) );
AND2x2_ASAP7_75t_L g592 ( .A(n_526), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g643 ( .A(n_526), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_526), .B(n_553), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_532), .Y(n_529) );
AND2x2_ASAP7_75t_L g554 ( .A(n_536), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g615 ( .A(n_536), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_536), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g652 ( .A(n_536), .Y(n_652) );
INVx1_ASAP7_75t_L g685 ( .A(n_536), .Y(n_685) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g563 ( .A(n_537), .B(n_553), .Y(n_563) );
INVx1_ASAP7_75t_L g593 ( .A(n_537), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_550), .B1(n_556), .B2(n_563), .C(n_564), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_547), .B(n_567), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_547), .B(n_630), .Y(n_707) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_549), .B(n_597), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_549), .B(n_558), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_549), .B(n_572), .Y(n_701) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g623 ( .A(n_553), .Y(n_623) );
AND2x2_ASAP7_75t_L g598 ( .A(n_554), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g676 ( .A(n_554), .Y(n_676) );
AND2x2_ASAP7_75t_L g608 ( .A(n_555), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_555), .B(n_578), .Y(n_624) );
AND2x2_ASAP7_75t_L g688 ( .A(n_555), .B(n_614), .Y(n_688) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g597 ( .A(n_559), .B(n_566), .Y(n_597) );
AND2x2_ASAP7_75t_L g693 ( .A(n_560), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_562), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_563), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_563), .B(n_570), .Y(n_658) );
AND2x2_ASAP7_75t_L g678 ( .A(n_563), .B(n_578), .Y(n_678) );
AND2x2_ASAP7_75t_L g699 ( .A(n_563), .B(n_643), .Y(n_699) );
OAI32xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .A3(n_570), .B1(n_571), .B2(n_574), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_SL g572 ( .A(n_566), .Y(n_572) );
NAND2x1_ASAP7_75t_L g613 ( .A(n_566), .B(n_596), .Y(n_613) );
OR2x2_ASAP7_75t_L g617 ( .A(n_566), .B(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_566), .B(n_665), .Y(n_718) );
INVx1_ASAP7_75t_L g586 ( .A(n_567), .Y(n_586) );
OAI221xp5_ASAP7_75t_SL g704 ( .A1(n_568), .A2(n_659), .B1(n_705), .B2(n_708), .C(n_709), .Y(n_704) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g576 ( .A(n_569), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g619 ( .A(n_569), .B(n_592), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_569), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g697 ( .A(n_569), .B(n_630), .Y(n_697) );
INVxp67_ASAP7_75t_L g633 ( .A(n_570), .Y(n_633) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AND2x2_ASAP7_75t_L g703 ( .A(n_572), .B(n_690), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_572), .B(n_653), .Y(n_726) );
INVx1_ASAP7_75t_L g601 ( .A(n_574), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_574), .B(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g719 ( .A(n_574), .B(n_720), .Y(n_719) );
OAI21xp5_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_579), .B(n_582), .Y(n_575) );
AND2x2_ASAP7_75t_L g588 ( .A(n_577), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g672 ( .A(n_581), .B(n_592), .Y(n_672) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AND2x2_ASAP7_75t_L g690 ( .A(n_583), .B(n_648), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_583), .B(n_647), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_584), .B(n_596), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_590), .C(n_600), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_586), .A2(n_621), .B1(n_625), .B2(n_628), .C(n_631), .Y(n_620) );
AOI31xp33_ASAP7_75t_L g715 ( .A1(n_586), .A2(n_716), .A3(n_717), .B(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_594), .B1(n_596), .B2(n_598), .Y(n_590) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g716 ( .A(n_596), .Y(n_716) );
INVx1_ASAP7_75t_L g679 ( .A(n_597), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g722 ( .A1(n_599), .A2(n_723), .B(n_725), .C(n_727), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_604), .B2(n_608), .Y(n_600) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_605), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI221xp5_ASAP7_75t_SL g695 ( .A1(n_607), .A2(n_641), .B1(n_660), .B2(n_696), .C(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g691 ( .A(n_608), .Y(n_691) );
INVx1_ASAP7_75t_L g645 ( .A(n_609), .Y(n_645) );
NAND3xp33_ASAP7_75t_SL g610 ( .A(n_611), .B(n_620), .C(n_635), .Y(n_610) );
OAI21xp33_ASAP7_75t_L g661 ( .A1(n_612), .A2(n_662), .B(n_666), .Y(n_661) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_614), .B(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g721 ( .A(n_615), .Y(n_721) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g659 ( .A(n_622), .B(n_642), .Y(n_659) );
INVx1_ASAP7_75t_L g634 ( .A(n_623), .Y(n_634) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g632 ( .A(n_626), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_626), .B(n_664), .Y(n_663) );
NOR4xp25_ASAP7_75t_L g631 ( .A(n_627), .B(n_632), .C(n_633), .D(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI222xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_640), .B1(n_646), .B2(n_647), .C1(n_649), .C2(n_653), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g733 ( .A(n_637), .Y(n_733) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_645), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_649), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI21xp5_ASAP7_75t_SL g709 ( .A1(n_654), .A2(n_710), .B(n_712), .Y(n_709) );
NOR4xp25_ASAP7_75t_L g655 ( .A(n_656), .B(n_667), .C(n_680), .D(n_695), .Y(n_655) );
OAI221xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_658), .B1(n_659), .B2(n_660), .C(n_661), .Y(n_656) );
INVx1_ASAP7_75t_L g736 ( .A(n_657), .Y(n_736) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_664), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
OAI222xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B1(n_673), .B2(n_674), .C1(n_677), .C2(n_679), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g702 ( .A1(n_672), .A2(n_703), .B(n_704), .C(n_715), .Y(n_702) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
OAI222xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_686), .B1(n_687), .B2(n_689), .C1(n_691), .C2(n_692), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_697), .A2(n_700), .B1(n_733), .B2(n_734), .Y(n_732) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI211xp5_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_730), .B(n_732), .C(n_735), .Y(n_727) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g745 ( .A(n_740), .Y(n_745) );
INVx3_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
endmodule