module fake_jpeg_8615_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_19),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_53),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_24),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_29),
.C(n_22),
.Y(n_68)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_48),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_28),
.B1(n_21),
.B2(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_59),
.B1(n_31),
.B2(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_60),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_31),
.B1(n_27),
.B2(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_30),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_4),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_75),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_29),
.B(n_30),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_6),
.C(n_14),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_68),
.B(n_71),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_34),
.B(n_33),
.C(n_22),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_52),
.B1(n_61),
.B2(n_56),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_76),
.B1(n_77),
.B2(n_80),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_22),
.B1(n_34),
.B2(n_33),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_81),
.B1(n_50),
.B2(n_47),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_34),
.B1(n_8),
.B2(n_9),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_91),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_90),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_93),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_56),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_50),
.B(n_48),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_70),
.B(n_78),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_67),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_106),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_52),
.B1(n_45),
.B2(n_44),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_45),
.B1(n_44),
.B2(n_55),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_55),
.B1(n_49),
.B2(n_62),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_103),
.A2(n_78),
.B1(n_67),
.B2(n_81),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_6),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_0),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_68),
.Y(n_114)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_115),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_66),
.C(n_77),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_128),
.B1(n_103),
.B2(n_14),
.Y(n_149)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_119),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_80),
.C(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_114),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_87),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_105),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_0),
.B(n_1),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_0),
.B(n_1),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_127),
.B1(n_85),
.B2(n_105),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_78),
.B1(n_70),
.B2(n_11),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_49),
.B1(n_78),
.B2(n_9),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_95),
.A3(n_96),
.B1(n_114),
.B2(n_115),
.C1(n_104),
.C2(n_97),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_138),
.C(n_146),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_132),
.B1(n_149),
.B2(n_141),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_99),
.B1(n_86),
.B2(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_133),
.B(n_134),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_119),
.B(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_139),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_104),
.A3(n_97),
.B1(n_102),
.B2(n_4),
.C1(n_14),
.C2(n_101),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_102),
.Y(n_140)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_97),
.B1(n_98),
.B2(n_92),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_148),
.B1(n_128),
.B2(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_101),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_105),
.C(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_123),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_127),
.B(n_122),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_139),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_124),
.B(n_123),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_110),
.B1(n_116),
.B2(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_164),
.B(n_134),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_114),
.A3(n_112),
.B1(n_125),
.B2(n_111),
.C1(n_113),
.C2(n_3),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_166),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_112),
.B(n_2),
.C(n_3),
.D(n_1),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_177),
.B(n_181),
.Y(n_188)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_137),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_167),
.B(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_148),
.C(n_137),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_182),
.C(n_150),
.Y(n_190)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_142),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_160),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_190),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_158),
.B(n_163),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_171),
.B(n_180),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_178),
.A2(n_149),
.B1(n_131),
.B2(n_154),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_143),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_172),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_193),
.C(n_174),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_153),
.Y(n_193)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_174),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_200),
.C(n_190),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_188),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_203),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_187),
.A2(n_168),
.B(n_175),
.C(n_154),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_202),
.C(n_183),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_201),
.B(n_194),
.Y(n_210)
);

OA21x2_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_146),
.B(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_112),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_184),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_202),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_199),
.Y(n_216)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_192),
.B(n_193),
.Y(n_209)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_194),
.B(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_210),
.B(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_214),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_199),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_216),
.B(n_199),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_207),
.C(n_205),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_218),
.B(n_215),
.C(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_222),
.A2(n_223),
.B(n_2),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_2),
.C(n_3),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_225),
.Y(n_227)
);


endmodule