module real_jpeg_15314_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_539),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_0),
.B(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_1),
.Y(n_85)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_1),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_2),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_2),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_2),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_2),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_3),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_3),
.A2(n_37),
.B1(n_290),
.B2(n_292),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_3),
.A2(n_37),
.B1(n_192),
.B2(n_392),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_3),
.A2(n_37),
.B1(n_431),
.B2(n_434),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_143),
.B1(n_146),
.B2(n_150),
.Y(n_142)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_4),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_4),
.A2(n_150),
.B1(n_228),
.B2(n_232),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_4),
.A2(n_150),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g524 ( 
.A1(n_4),
.A2(n_150),
.B1(n_359),
.B2(n_525),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_5),
.A2(n_157),
.B1(n_160),
.B2(n_163),
.Y(n_156)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_5),
.A2(n_163),
.B1(n_258),
.B2(n_261),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_5),
.A2(n_105),
.B1(n_163),
.B2(n_344),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_6),
.Y(n_141)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_6),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_6),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g438 ( 
.A(n_6),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_7),
.A2(n_191),
.B1(n_192),
.B2(n_196),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_7),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_7),
.A2(n_191),
.B1(n_216),
.B2(n_221),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_7),
.A2(n_191),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_7),
.A2(n_191),
.B1(n_359),
.B2(n_361),
.Y(n_358)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_8),
.Y(n_540)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_9),
.Y(n_176)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_9),
.Y(n_195)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_9),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_9),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_9),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_9),
.Y(n_410)
);

BUFx5_ASAP7_75t_L g465 ( 
.A(n_9),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_10),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_10),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_10),
.A2(n_104),
.B1(n_268),
.B2(n_271),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_10),
.A2(n_104),
.B1(n_397),
.B2(n_398),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g458 ( 
.A1(n_10),
.A2(n_104),
.B1(n_459),
.B2(n_461),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_11),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_11),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_11),
.A2(n_111),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_11),
.A2(n_111),
.B1(n_247),
.B2(n_250),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_11),
.A2(n_111),
.B1(n_201),
.B2(n_327),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_13),
.A2(n_116),
.A3(n_118),
.B1(n_119),
.B2(n_125),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_13),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_13),
.A2(n_124),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_13),
.B(n_42),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_13),
.B(n_71),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_13),
.B(n_189),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_13),
.B(n_448),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g467 ( 
.A1(n_13),
.A2(n_120),
.B1(n_124),
.B2(n_206),
.Y(n_467)
);

OAI32xp33_ASAP7_75t_L g469 ( 
.A1(n_13),
.A2(n_470),
.A3(n_473),
.B1(n_476),
.B2(n_477),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_16),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_16),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_16),
.Y(n_220)
);

BUFx4f_ASAP7_75t_L g446 ( 
.A(n_16),
.Y(n_446)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g270 ( 
.A(n_17),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_514),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_508),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_366),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_303),
.C(n_333),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_281),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_237),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_26),
.B(n_237),
.C(n_510),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_164),
.C(n_210),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_27),
.B(n_302),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_114),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_68),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_29),
.B(n_68),
.C(n_114),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_40),
.B1(n_42),
.B2(n_60),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_31),
.A2(n_41),
.B1(n_200),
.B2(n_203),
.Y(n_199)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g360 ( 
.A(n_34),
.Y(n_360)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_36),
.Y(n_129)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_40),
.B(n_358),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_41),
.A2(n_61),
.B1(n_203),
.B2(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_41),
.A2(n_267),
.B(n_325),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_41),
.A2(n_356),
.B(n_357),
.Y(n_355)
);

OR2x6_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_42),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_42),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_42),
.B(n_358),
.Y(n_357)
);

AO22x2_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_45),
.Y(n_209)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_46),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_48),
.Y(n_279)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_48),
.Y(n_472)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_55),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_56),
.Y(n_271)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_61)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_62),
.Y(n_202)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_64),
.A2(n_67),
.B1(n_100),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_64),
.A2(n_67),
.B1(n_407),
.B2(n_409),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_64),
.A2(n_67),
.B1(n_417),
.B2(n_421),
.Y(n_416)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_65),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_98),
.B(n_107),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_69),
.A2(n_71),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

AOI21x1_ASAP7_75t_SL g529 ( 
.A1(n_69),
.A2(n_343),
.B(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_70),
.A2(n_99),
.B1(n_108),
.B2(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_70),
.A2(n_109),
.B(n_273),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_70),
.A2(n_108),
.B1(n_205),
.B2(n_289),
.Y(n_288)
);

OAI22x1_ASAP7_75t_L g317 ( 
.A1(n_70),
.A2(n_108),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_70),
.A2(n_108),
.B1(n_289),
.B2(n_467),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_82),
.Y(n_70)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_71),
.B(n_274),
.Y(n_273)
);

AO22x2_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B1(n_78),
.B2(n_80),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g168 ( 
.A1(n_75),
.A2(n_169),
.B1(n_172),
.B2(n_174),
.Y(n_168)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_77),
.Y(n_198)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_77),
.Y(n_231)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_89),
.B2(n_94),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_97),
.Y(n_480)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_106),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_113),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_131),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_115),
.B(n_131),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_123),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_124),
.B(n_192),
.Y(n_381)
);

OAI21xp33_ASAP7_75t_SL g386 ( 
.A1(n_124),
.A2(n_381),
.B(n_387),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_124),
.A2(n_133),
.B1(n_430),
.B2(n_437),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_124),
.B(n_373),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_129),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_142),
.B1(n_151),
.B2(n_156),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_132),
.A2(n_156),
.B(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_132),
.A2(n_415),
.B1(n_423),
.B2(n_424),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_132),
.A2(n_212),
.B(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_133),
.B(n_215),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_133),
.A2(n_246),
.B(n_310),
.Y(n_309)
);

AOI21x1_ASAP7_75t_L g395 ( 
.A1(n_133),
.A2(n_396),
.B(n_403),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_133),
.A2(n_416),
.B1(n_430),
.B2(n_435),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_134),
.Y(n_434)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_136),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_138),
.Y(n_310)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_140),
.Y(n_245)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_141),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_142),
.A2(n_254),
.B(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_149),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_149),
.Y(n_422)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_149),
.Y(n_433)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_164),
.B(n_210),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_199),
.C(n_204),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_165),
.B(n_204),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_182),
.B(n_188),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_166),
.A2(n_177),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g312 ( 
.A1(n_166),
.A2(n_188),
.B(n_257),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_166),
.A2(n_177),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_167),
.B(n_190),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_167),
.A2(n_189),
.B1(n_386),
.B2(n_391),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_167),
.A2(n_189),
.B1(n_391),
.B2(n_406),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_167),
.A2(n_350),
.B(n_499),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_167),
.A2(n_183),
.B(n_189),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_177),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_175),
.Y(n_393)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_176),
.Y(n_376)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_177),
.B(n_184),
.Y(n_350)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_179),
.Y(n_253)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_180),
.Y(n_397)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_181),
.Y(n_383)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_187),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_227),
.Y(n_226)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_199),
.B(n_284),
.Y(n_283)
);

OAI21x1_ASAP7_75t_SL g523 ( 
.A1(n_203),
.A2(n_524),
.B(n_526),
.Y(n_523)
);

INVx3_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_209),
.Y(n_323)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_209),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_225),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_211),
.B(n_225),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_219),
.Y(n_402)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_236),
.Y(n_225)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_231),
.Y(n_475)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_236),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_238),
.B(n_262),
.C(n_280),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_262),
.B1(n_263),
.B2(n_280),
.Y(n_239)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_255),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_241),
.B(n_255),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_254),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_242),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_246),
.Y(n_487)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_253),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_R g330 ( 
.A(n_264),
.B(n_266),
.C(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_272),
.Y(n_265)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_270),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_272),
.Y(n_331)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_273),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_301),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_282),
.B(n_301),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.C(n_287),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_283),
.B(n_504),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_287),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_294),
.C(n_296),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_288),
.B(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_296),
.Y(n_495)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_300),
.Y(n_424)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g508 ( 
.A1(n_304),
.A2(n_509),
.B(n_511),
.C(n_512),
.D(n_513),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_305),
.B(n_306),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_329),
.B1(n_330),
.B2(n_332),
.Y(n_306)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_314),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_314),
.C(n_329),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_309),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_309),
.A2(n_313),
.B1(n_355),
.B2(n_364),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_309),
.B(n_312),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI21xp33_ASAP7_75t_L g535 ( 
.A1(n_313),
.A2(n_364),
.B(n_536),
.Y(n_535)
);

XNOR2x1_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_324),
.C(n_337),
.Y(n_336)
);

XNOR2x1_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_324),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_317),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_326),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_333),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_334),
.B(n_335),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_336),
.B(n_339),
.C(n_353),
.Y(n_517)
);

XNOR2x1_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_353),
.Y(n_338)
);

OA21x2_ASAP7_75t_SL g339 ( 
.A1(n_340),
.A2(n_349),
.B(n_352),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_349),
.Y(n_352)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_352),
.A2(n_521),
.B1(n_532),
.B2(n_533),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_352),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_365),
.Y(n_353)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_355),
.Y(n_364)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_365),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_502),
.B(n_507),
.Y(n_366)
);

AOI21x1_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_489),
.B(n_501),
.Y(n_367)
);

OAI21x1_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_452),
.B(n_488),
.Y(n_368)
);

AOI21x1_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_412),
.B(n_451),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_394),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_371),
.B(n_394),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_384),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_372),
.A2(n_384),
.B1(n_385),
.B2(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_372),
.Y(n_426)
);

OAI32xp33_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_377),
.A3(n_379),
.B1(n_381),
.B2(n_382),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_378),
.B(n_383),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_404),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_395),
.B(n_405),
.C(n_411),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_411),
.Y(n_404)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_406),
.Y(n_457)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_409),
.Y(n_460)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_413),
.A2(n_427),
.B(n_450),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_425),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_425),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

AOI21x1_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_440),
.B(n_449),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_439),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_439),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx6_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

BUFx12f_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_447),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_453),
.B(n_454),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_468),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_466),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_456),
.B(n_466),
.C(n_468),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_458),
.Y(n_499)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_486),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_486),
.Y(n_497)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_481),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_SL g501 ( 
.A(n_490),
.B(n_491),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_493),
.B1(n_496),
.B2(n_500),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_497),
.C(n_498),
.Y(n_506)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_496),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NOR2xp67_ASAP7_75t_SL g502 ( 
.A(n_503),
.B(n_506),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_506),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_538),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

NOR2xp67_ASAP7_75t_SL g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_517),
.B(n_518),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_519),
.A2(n_520),
.B1(n_534),
.B2(n_535),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_521),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_523),
.B1(n_527),
.B2(n_531),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_527),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.Y(n_527)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);


endmodule