module real_jpeg_25794_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_32),
.B1(n_37),
.B2(n_41),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_3),
.A2(n_32),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_32),
.B1(n_52),
.B2(n_56),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_5),
.A2(n_52),
.B1(n_56),
.B2(n_60),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_5),
.A2(n_37),
.B1(n_41),
.B2(n_60),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_60),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_8),
.A2(n_25),
.B1(n_37),
.B2(n_41),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_10),
.A2(n_37),
.B1(n_41),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_10),
.A2(n_44),
.B1(n_52),
.B2(n_56),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_44),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_10),
.A2(n_55),
.B(n_103),
.C(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_10),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_10),
.B(n_51),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_10),
.A2(n_56),
.B(n_72),
.C(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_10),
.B(n_24),
.C(n_40),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_10),
.B(n_127),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_10),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_10),
.B(n_42),
.Y(n_200)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_11),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_11),
.B(n_183),
.Y(n_188)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_11),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_130),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_128),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_106),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_15),
.B(n_106),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_91),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_79),
.B2(n_80),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_47),
.B2(n_48),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_21),
.B(n_33),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_28),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_22),
.A2(n_30),
.B(n_90),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_23),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_24),
.B(n_194),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_26),
.B(n_31),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_26),
.B(n_89),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_26),
.A2(n_89),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_26),
.B(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_29),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_29),
.B(n_181),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_45),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_34),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_43),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_35),
.B(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_35),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_35),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_36)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_37),
.A2(n_41),
.B1(n_72),
.B2(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_37),
.B(n_171),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_41),
.A2(n_44),
.B(n_74),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_42),
.B(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_44),
.A2(n_54),
.B(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_45),
.B(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_68),
.B1(n_69),
.B2(n_78),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_61),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_65),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_56),
.B1(n_72),
.B2(n_74),
.Y(n_71)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_55),
.B1(n_59),
.B2(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_62),
.Y(n_95)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_117),
.Y(n_116)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_75),
.B(n_76),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_70),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_70),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_75),
.B(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_77),
.B(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_82),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_82),
.B(n_121),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_84),
.B(n_168),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_86),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_90),
.B(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_101),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_105),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_112),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_107),
.A2(n_108),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_228),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_111),
.Y(n_228)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_122),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_115),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_126),
.B(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_229),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_223),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_162),
.B(n_222),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_152),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_134),
.B(n_152),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_142),
.C(n_147),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_135),
.B(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_138),
.C(n_140),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_139),
.B(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_142),
.B(n_147),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_143),
.A2(n_145),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_143),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_145),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_155),
.B(n_156),
.C(n_157),
.Y(n_224)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_217),
.B(n_221),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_205),
.B(n_216),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_185),
.B(n_204),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_166),
.B(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_169),
.B1(n_170),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_179),
.B2(n_184),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_178),
.C(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_179),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_191),
.B(n_203),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_189),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_188),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_199),
.B(n_202),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_200),
.B(n_201),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_206),
.B(n_207),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);


endmodule