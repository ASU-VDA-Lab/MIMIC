module fake_jpeg_18059_n_62 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_7),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_8),
.C(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_12),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_12),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_10),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_20),
.B1(n_19),
.B2(n_9),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_20),
.B1(n_9),
.B2(n_14),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_1),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_1),
.B(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_5),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_21),
.C(n_22),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_4),
.Y(n_37)
);

XOR2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_44),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_43),
.B(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_13),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_42),
.C(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_52),
.B(n_27),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_51),
.B(n_13),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_50),
.C(n_21),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_18),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_57),
.B(n_5),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_59),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_15),
.C(n_18),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_15),
.Y(n_62)
);


endmodule