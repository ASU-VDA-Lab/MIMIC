module fake_jpeg_22039_n_77 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_46),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_3),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_33),
.B1(n_6),
.B2(n_9),
.Y(n_55)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_50),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_53),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_34),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_15),
.B(n_16),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_5),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_10),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_63),
.C(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_65),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_67),
.B1(n_64),
.B2(n_69),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_31),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_21),
.B(n_23),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_30),
.Y(n_77)
);


endmodule