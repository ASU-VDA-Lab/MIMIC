module fake_jpeg_10077_n_258 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx8_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_17),
.B1(n_25),
.B2(n_29),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_22),
.B1(n_29),
.B2(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_55),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_43),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_18),
.B1(n_32),
.B2(n_30),
.Y(n_59)
);

AO22x1_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_22),
.B1(n_28),
.B2(n_27),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_37),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_74),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_43),
.B1(n_40),
.B2(n_17),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_72),
.B1(n_85),
.B2(n_40),
.Y(n_95)
);

XNOR2x1_ASAP7_75t_SL g115 ( 
.A(n_68),
.B(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_40),
.B1(n_17),
.B2(n_50),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_23),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_84),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_18),
.B1(n_24),
.B2(n_26),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_0),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_31),
.B(n_23),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_34),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_28),
.Y(n_107)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_56),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_91),
.A2(n_113),
.B(n_81),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_95),
.A2(n_111),
.B1(n_64),
.B2(n_24),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_64),
.B(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_104),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_36),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_105),
.C(n_116),
.Y(n_128)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_106),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_37),
.B(n_39),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_103),
.B1(n_115),
.B2(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_20),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_61),
.C(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_81),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_20),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_109),
.B(n_110),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_31),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_1),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_36),
.C(n_57),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_119),
.Y(n_157)
);

AO21x2_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_68),
.B(n_65),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_141),
.B(n_84),
.C(n_80),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_67),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_135),
.C(n_142),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_69),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_127),
.B(n_134),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_130),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

NAND2x1p5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_85),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_112),
.B(n_34),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_93),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_133),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_70),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_92),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_91),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_143),
.B(n_113),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_92),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_78),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_112),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_73),
.B1(n_37),
.B2(n_39),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_36),
.C(n_78),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_145),
.B(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_153),
.B(n_160),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_96),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_168),
.Y(n_177)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_100),
.B1(n_95),
.B2(n_113),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_161),
.A2(n_137),
.B1(n_121),
.B2(n_123),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_114),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_103),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_129),
.C(n_34),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_37),
.B1(n_39),
.B2(n_88),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_166),
.B(n_169),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_118),
.B(n_26),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_138),
.B(n_143),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_131),
.B1(n_126),
.B2(n_127),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_172),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_187),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_128),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_166),
.B(n_156),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_184),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_181),
.B1(n_191),
.B2(n_159),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_137),
.B1(n_133),
.B2(n_30),
.Y(n_181)
);

OA21x2_ASAP7_75t_SL g183 ( 
.A1(n_165),
.A2(n_34),
.B(n_12),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_183),
.B(n_168),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_167),
.C(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_146),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_192),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_160),
.A2(n_32),
.B1(n_86),
.B2(n_16),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_16),
.C(n_15),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_205),
.B(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_196),
.B(n_199),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_151),
.B1(n_164),
.B2(n_144),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_181),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_159),
.B1(n_161),
.B2(n_155),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_171),
.B1(n_174),
.B2(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_170),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_204),
.C(n_209),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_167),
.C(n_163),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_150),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_176),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_147),
.C(n_145),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_216),
.C(n_217),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_213),
.B(n_215),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_174),
.C(n_175),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_179),
.C(n_186),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_221),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_173),
.B(n_179),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_197),
.B1(n_193),
.B2(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_157),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_228),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_212),
.B(n_209),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_227),
.Y(n_242)
);

AO21x1_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_198),
.B(n_200),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_196),
.C(n_194),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_214),
.C(n_217),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_13),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_233),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_86),
.B1(n_2),
.B2(n_3),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_216),
.A3(n_211),
.B1(n_13),
.B2(n_12),
.C1(n_7),
.C2(n_10),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_238),
.C(n_241),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_31),
.C(n_3),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_225),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_239),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_31),
.C(n_5),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_233),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_247),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_237),
.A2(n_224),
.B1(n_5),
.B2(n_6),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_245),
.B1(n_248),
.B2(n_242),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_1),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_244),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_249),
.A2(n_252),
.B(n_10),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_6),
.C(n_10),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_6),
.B(n_7),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_247),
.B(n_244),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_253),
.A2(n_255),
.B(n_11),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_254),
.A2(n_11),
.B(n_245),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.Y(n_258)
);


endmodule