module fake_jpeg_2041_n_611 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_611);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_611;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_59),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_60),
.B(n_61),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_67),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_26),
.B(n_18),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_69),
.B(n_27),
.C(n_49),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_70),
.Y(n_187)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx11_ASAP7_75t_L g218 ( 
.A(n_71),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_72),
.Y(n_168)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g175 ( 
.A(n_73),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_13),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_99),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_75),
.B(n_77),
.Y(n_184)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_79),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_80),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_19),
.B(n_16),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_109),
.Y(n_137)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_82),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_83),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

CKINVDCx6p67_ASAP7_75t_R g165 ( 
.A(n_86),
.Y(n_165)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_88),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_91),
.Y(n_204)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_92),
.Y(n_149)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_93),
.Y(n_212)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_94),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_95),
.Y(n_215)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_97),
.Y(n_203)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_21),
.B(n_13),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_13),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_101),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_16),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_102),
.Y(n_216)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_103),
.Y(n_205)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_104),
.Y(n_211)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_26),
.B(n_10),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_113),
.Y(n_219)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_32),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_34),
.B(n_10),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_0),
.Y(n_148)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_37),
.Y(n_119)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_34),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_121),
.B(n_27),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_39),
.B(n_0),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_124),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_24),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_37),
.Y(n_125)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_32),
.Y(n_127)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_56),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_140),
.B(n_143),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_56),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_148),
.B(n_159),
.Y(n_257)
);

BUFx12_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_150),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_101),
.A2(n_123),
.B1(n_74),
.B2(n_42),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g300 ( 
.A1(n_151),
.A2(n_210),
.B1(n_216),
.B2(n_215),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_42),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_155),
.B(n_157),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_92),
.B(n_41),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_39),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_107),
.B(n_41),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_160),
.B(n_177),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_84),
.A2(n_25),
.B1(n_54),
.B2(n_51),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_164),
.A2(n_49),
.B1(n_44),
.B2(n_31),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_25),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_166),
.B(n_176),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_110),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_170),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_111),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_73),
.B(n_55),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_95),
.B(n_24),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_178),
.B(n_0),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_188),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_102),
.B(n_28),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_96),
.B(n_55),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_192),
.B(n_194),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_62),
.B(n_54),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_58),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_202),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_108),
.B(n_23),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_68),
.B(n_33),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g295 ( 
.A(n_206),
.B(n_220),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_122),
.B(n_51),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_214),
.Y(n_230)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_79),
.Y(n_209)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_70),
.A2(n_50),
.B1(n_28),
.B2(n_30),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_125),
.B(n_33),
.Y(n_214)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_93),
.Y(n_217)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_72),
.B(n_50),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_119),
.B(n_30),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_44),
.Y(n_237)
);

CKINVDCx9p33_ASAP7_75t_R g222 ( 
.A(n_165),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_222),
.Y(n_313)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_223),
.Y(n_316)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_141),
.Y(n_224)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_224),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_151),
.A2(n_85),
.B1(n_91),
.B2(n_88),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_227),
.A2(n_233),
.B1(n_265),
.B2(n_168),
.Y(n_303)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_139),
.Y(n_229)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_229),
.Y(n_312)
);

BUFx12_ASAP7_75t_L g234 ( 
.A(n_150),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g327 ( 
.A(n_234),
.Y(n_327)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_235),
.Y(n_319)
);

CKINVDCx9p33_ASAP7_75t_R g236 ( 
.A(n_165),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_236),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_237),
.B(n_242),
.Y(n_334)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_144),
.Y(n_238)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_238),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_132),
.A2(n_31),
.B1(n_23),
.B2(n_32),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_239),
.A2(n_271),
.B1(n_275),
.B2(n_281),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_240),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_241),
.B(n_244),
.Y(n_340)
);

CKINVDCx12_ASAP7_75t_R g242 ( 
.A(n_179),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_144),
.Y(n_243)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_243),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_133),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_138),
.A2(n_112),
.B(n_32),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_245),
.A2(n_210),
.B(n_175),
.Y(n_307)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_174),
.Y(n_248)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_248),
.Y(n_301)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_249),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_184),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_250),
.B(n_253),
.Y(n_344)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_129),
.Y(n_251)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_147),
.Y(n_252)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_252),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_176),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_134),
.B(n_112),
.C(n_2),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_254),
.B(n_263),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_147),
.Y(n_255)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_255),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_156),
.Y(n_258)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_258),
.Y(n_322)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_145),
.Y(n_259)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_259),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_156),
.Y(n_260)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_260),
.Y(n_338)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_218),
.Y(n_261)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_261),
.Y(n_345)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_161),
.Y(n_262)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_262),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_130),
.B(n_1),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_263),
.B(n_273),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_132),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_190),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_266),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_138),
.B(n_5),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_268),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_155),
.B(n_6),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_177),
.A2(n_188),
.B1(n_208),
.B2(n_164),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_269),
.A2(n_172),
.B1(n_191),
.B2(n_204),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_183),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_195),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_274),
.Y(n_308)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_161),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_193),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_152),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_161),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_276),
.B(n_278),
.Y(n_311)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_207),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_285),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_140),
.B(n_7),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_187),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_282),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_162),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_201),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_196),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_283),
.B(n_284),
.Y(n_346)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_131),
.Y(n_284)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_215),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_130),
.B(n_9),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_287),
.A2(n_298),
.B(n_153),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_192),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_288),
.B(n_289),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_168),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_143),
.B(n_157),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_291),
.B(n_293),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_165),
.A2(n_199),
.B1(n_149),
.B2(n_167),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g330 ( 
.A1(n_292),
.A2(n_154),
.B1(n_182),
.B2(n_219),
.Y(n_330)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_133),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_202),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_294),
.B(n_296),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_137),
.B(n_135),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_203),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_299),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_142),
.B(n_136),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_205),
.B(n_211),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_300),
.A2(n_266),
.B1(n_248),
.B2(n_249),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_303),
.A2(n_305),
.B1(n_333),
.B2(n_335),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_146),
.B1(n_212),
.B2(n_171),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_307),
.B(n_315),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_309),
.B(n_244),
.Y(n_359)
);

AO22x2_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_189),
.B1(n_181),
.B2(n_173),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_300),
.A2(n_216),
.B1(n_146),
.B2(n_171),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_324),
.A2(n_326),
.B1(n_339),
.B2(n_238),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_295),
.A2(n_212),
.B1(n_172),
.B2(n_197),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_328),
.B(n_353),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_247),
.B(n_198),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_329),
.B(n_332),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_330),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_231),
.B(n_198),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_230),
.A2(n_204),
.B1(n_191),
.B2(n_197),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_228),
.A2(n_185),
.B1(n_270),
.B2(n_280),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_185),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_343),
.C(n_351),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_257),
.B(n_185),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_241),
.A2(n_290),
.B1(n_287),
.B2(n_226),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_348),
.A2(n_354),
.B1(n_275),
.B2(n_255),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_298),
.B(n_232),
.Y(n_351)
);

AO22x2_ASAP7_75t_L g353 ( 
.A1(n_224),
.A2(n_235),
.B1(n_259),
.B2(n_243),
.Y(n_353)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_358),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_359),
.B(n_368),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_356),
.B(n_348),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_360),
.B(n_361),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_318),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_349),
.B(n_225),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_362),
.B(n_366),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_246),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_364),
.B(n_365),
.C(n_367),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_264),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_328),
.B(n_351),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_240),
.C(n_286),
.Y(n_367)
);

AND2x6_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_286),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_304),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_369),
.B(n_371),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_301),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_370),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_306),
.B(n_293),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_319),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_372),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_355),
.B(n_297),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_373),
.B(n_375),
.Y(n_438)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_314),
.Y(n_374)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_374),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_334),
.B(n_279),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_307),
.A2(n_292),
.B(n_261),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_376),
.A2(n_315),
.B(n_320),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_311),
.B(n_262),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_380),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_341),
.B(n_340),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_393),
.Y(n_415)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_379),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_316),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_SL g433 ( 
.A1(n_381),
.A2(n_322),
.B1(n_337),
.B2(n_317),
.Y(n_433)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_347),
.Y(n_384)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_384),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_302),
.B(n_273),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_385),
.B(n_386),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_316),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_321),
.B(n_276),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_388),
.Y(n_414)
);

AND2x2_ASAP7_75t_SL g390 ( 
.A(n_340),
.B(n_289),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_390),
.B(n_391),
.Y(n_428)
);

AO22x1_ASAP7_75t_L g391 ( 
.A1(n_326),
.A2(n_285),
.B1(n_271),
.B2(n_281),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_336),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_392),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_346),
.B(n_252),
.Y(n_393)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_347),
.Y(n_395)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_395),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_396),
.A2(n_315),
.B1(n_305),
.B2(n_301),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_341),
.B(n_234),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_397),
.B(n_330),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_303),
.B(n_258),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_399),
.Y(n_419)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_325),
.B(n_260),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_402),
.Y(n_427)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_352),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_363),
.B(n_354),
.C(n_312),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_409),
.B(n_426),
.C(n_429),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_394),
.A2(n_324),
.B1(n_350),
.B2(n_335),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_411),
.A2(n_413),
.B1(n_425),
.B2(n_382),
.Y(n_446)
);

AO22x1_ASAP7_75t_L g412 ( 
.A1(n_389),
.A2(n_400),
.B1(n_396),
.B2(n_374),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_412),
.B(n_431),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_387),
.Y(n_421)
);

INVx13_ASAP7_75t_L g468 ( 
.A(n_421),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_389),
.A2(n_315),
.B1(n_333),
.B2(n_353),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_422),
.A2(n_391),
.B1(n_376),
.B2(n_383),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_382),
.A2(n_320),
.B1(n_353),
.B2(n_352),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_363),
.B(n_312),
.C(n_310),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_366),
.B(n_353),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_365),
.B(n_345),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_432),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_362),
.B(n_338),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_433),
.A2(n_379),
.B1(n_402),
.B2(n_399),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_400),
.A2(n_330),
.B(n_327),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_439),
.A2(n_359),
.B(n_378),
.Y(n_467)
);

BUFx10_ASAP7_75t_L g442 ( 
.A(n_421),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_442),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_358),
.Y(n_443)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_443),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_400),
.Y(n_444)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_444),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_414),
.B(n_371),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_445),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_446),
.A2(n_467),
.B(n_439),
.Y(n_483)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_427),
.Y(n_447)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_447),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_416),
.B(n_401),
.Y(n_448)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_448),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_435),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_449),
.B(n_406),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_416),
.A2(n_381),
.B1(n_389),
.B2(n_398),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_450),
.B(n_457),
.Y(n_480)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_451),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_438),
.B(n_360),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g492 ( 
.A(n_453),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_408),
.B(n_364),
.Y(n_454)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_454),
.Y(n_500)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_417),
.Y(n_455)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_455),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_456),
.A2(n_472),
.B1(n_428),
.B2(n_422),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_424),
.A2(n_367),
.B1(n_368),
.B2(n_391),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_420),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_466),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_436),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_461),
.Y(n_481)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_419),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_460),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_408),
.B(n_390),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_405),
.B(n_397),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_464),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_437),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_463),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_403),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_404),
.A2(n_390),
.B1(n_372),
.B2(n_395),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_471),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_403),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_470),
.B(n_473),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_404),
.A2(n_419),
.B1(n_420),
.B2(n_429),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_412),
.A2(n_384),
.B1(n_370),
.B2(n_313),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_423),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_443),
.B(n_460),
.Y(n_474)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_474),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_483),
.A2(n_494),
.B(n_498),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_447),
.B(n_415),
.Y(n_484)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_484),
.Y(n_514)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_487),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_426),
.C(n_407),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_488),
.B(n_489),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_407),
.C(n_430),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_452),
.B(n_409),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_491),
.B(n_462),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_454),
.B(n_434),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_493),
.B(n_444),
.C(n_467),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_441),
.A2(n_432),
.B(n_428),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_452),
.B(n_415),
.C(n_410),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_496),
.B(n_461),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_441),
.A2(n_428),
.B(n_412),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_SL g526 ( 
.A1(n_501),
.A2(n_442),
.B1(n_463),
.B2(n_459),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_466),
.B(n_423),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_504),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_505),
.B(n_507),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_497),
.B(n_457),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_478),
.B(n_470),
.Y(n_508)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_508),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_478),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_509),
.B(n_520),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_510),
.A2(n_511),
.B1(n_530),
.B2(n_490),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_501),
.A2(n_456),
.B1(n_450),
.B2(n_440),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_503),
.B(n_448),
.Y(n_513)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_513),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_491),
.B(n_440),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_515),
.B(n_517),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_475),
.Y(n_516)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_516),
.Y(n_536)
);

AOI21x1_ASAP7_75t_L g517 ( 
.A1(n_494),
.A2(n_469),
.B(n_473),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_518),
.B(n_519),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_500),
.B(n_472),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_481),
.Y(n_520)
);

XOR2x1_ASAP7_75t_L g522 ( 
.A(n_477),
.B(n_468),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_522),
.B(n_498),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_500),
.B(n_488),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_523),
.B(n_484),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_480),
.A2(n_451),
.B1(n_455),
.B2(n_468),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_524),
.A2(n_497),
.B1(n_485),
.B2(n_477),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_463),
.Y(n_525)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_525),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_526),
.A2(n_528),
.B1(n_507),
.B2(n_511),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_479),
.Y(n_529)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_529),
.Y(n_548)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_481),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_489),
.C(n_504),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_533),
.B(n_546),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_535),
.A2(n_543),
.B1(n_547),
.B2(n_525),
.Y(n_552)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_537),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_539),
.B(n_508),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_541),
.A2(n_539),
.B1(n_545),
.B2(n_531),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_506),
.A2(n_480),
.B1(n_490),
.B2(n_485),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_523),
.B(n_515),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_544),
.B(n_533),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_518),
.B(n_528),
.C(n_517),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_506),
.A2(n_486),
.B1(n_476),
.B2(n_495),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_SL g557 ( 
.A(n_549),
.B(n_519),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_507),
.B(n_483),
.C(n_486),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_550),
.B(n_529),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_551),
.B(n_556),
.Y(n_571)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_552),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_557),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_549),
.B(n_522),
.Y(n_556)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_542),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_558),
.B(n_560),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_538),
.B(n_524),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_559),
.B(n_564),
.Y(n_576)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_535),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_561),
.B(n_563),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_562),
.A2(n_547),
.B1(n_534),
.B2(n_514),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_546),
.B(n_530),
.C(n_482),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_536),
.B(n_527),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_538),
.B(n_482),
.C(n_512),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_565),
.B(n_540),
.C(n_532),
.Y(n_567)
);

INVx13_ASAP7_75t_L g566 ( 
.A(n_548),
.Y(n_566)
);

INVxp33_ASAP7_75t_L g579 ( 
.A(n_566),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_567),
.B(n_572),
.Y(n_588)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_566),
.Y(n_569)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_569),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_551),
.B(n_550),
.C(n_544),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_563),
.B(n_532),
.C(n_543),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_574),
.B(n_556),
.Y(n_584)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_575),
.Y(n_587)
);

FAx1_ASAP7_75t_SL g577 ( 
.A(n_565),
.B(n_474),
.CI(n_476),
.CON(n_577),
.SN(n_577)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_577),
.A2(n_555),
.B1(n_568),
.B2(n_553),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_554),
.B(n_492),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_578),
.B(n_499),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_571),
.B(n_562),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_581),
.B(n_584),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_583),
.B(n_586),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_573),
.A2(n_495),
.B1(n_513),
.B2(n_502),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_585),
.B(n_589),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_571),
.B(n_559),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_576),
.A2(n_557),
.B1(n_502),
.B2(n_499),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_590),
.B(n_580),
.Y(n_591)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_591),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_588),
.B(n_572),
.Y(n_593)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_593),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_583),
.A2(n_567),
.B(n_574),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_594),
.A2(n_581),
.B1(n_587),
.B2(n_589),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_586),
.B(n_570),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_595),
.B(n_579),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_599),
.B(n_601),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_592),
.A2(n_579),
.B1(n_582),
.B2(n_569),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_602),
.B(n_597),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_599),
.Y(n_604)
);

AOI322xp5_ASAP7_75t_L g606 ( 
.A1(n_604),
.A2(n_605),
.A3(n_597),
.B1(n_600),
.B2(n_596),
.C1(n_598),
.C2(n_577),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_606),
.Y(n_607)
);

A2O1A1O1Ixp25_ASAP7_75t_L g608 ( 
.A1(n_607),
.A2(n_603),
.B(n_577),
.C(n_575),
.D(n_442),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_608),
.B(n_442),
.C(n_418),
.Y(n_609)
);

OAI311xp33_ASAP7_75t_L g610 ( 
.A1(n_609),
.A2(n_418),
.A3(n_437),
.B1(n_327),
.C1(n_234),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_610),
.B(n_327),
.Y(n_611)
);


endmodule