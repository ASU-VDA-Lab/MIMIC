module real_jpeg_18648_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_2),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_2),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_3),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_3),
.A2(n_92),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_3),
.A2(n_92),
.B1(n_156),
.B2(n_160),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g193 ( 
.A1(n_3),
.A2(n_92),
.B1(n_194),
.B2(n_198),
.Y(n_193)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_4),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_5),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_5),
.Y(n_166)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_5),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_5),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_6),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_7),
.A2(n_322),
.B1(n_326),
.B2(n_327),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_7),
.Y(n_326)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_8),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_9),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_9),
.A2(n_52),
.B1(n_98),
.B2(n_102),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_9),
.A2(n_46),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_9),
.B(n_177),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_9),
.A2(n_68),
.A3(n_226),
.B1(n_227),
.B2(n_230),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_9),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_9),
.B(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_10),
.Y(n_159)
);

BUFx4f_ASAP7_75t_L g325 ( 
.A(n_10),
.Y(n_325)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_11),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_11),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_311),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_217),
.B(n_308),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_182),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_16),
.B(n_182),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.C(n_174),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_17),
.B(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_95),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_54),
.B2(n_55),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_20),
.B(n_54),
.C(n_95),
.Y(n_216)
);

AOI21x1_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_30),
.B(n_44),
.Y(n_20)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_21),
.Y(n_281)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2x1_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_33),
.Y(n_32)
);

AO22x2_ASAP7_75t_L g192 ( 
.A1(n_22),
.A2(n_32),
.B1(n_45),
.B2(n_193),
.Y(n_192)
);

AO22x1_ASAP7_75t_L g243 ( 
.A1(n_22),
.A2(n_32),
.B1(n_45),
.B2(n_193),
.Y(n_243)
);

AO22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_29),
.Y(n_22)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_24),
.Y(n_154)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_25),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_26),
.Y(n_209)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_28),
.Y(n_263)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_35),
.Y(n_199)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_42),
.Y(n_226)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_42),
.Y(n_232)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B(n_51),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_51),
.A2(n_154),
.A3(n_250),
.B1(n_254),
.B2(n_258),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_52),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_54),
.A2(n_55),
.B1(n_192),
.B2(n_214),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_54),
.B(n_192),
.C(n_224),
.Y(n_301)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_66),
.B1(n_78),
.B2(n_87),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_56),
.A2(n_66),
.B1(n_78),
.B2(n_87),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_56),
.A2(n_66),
.B(n_78),
.Y(n_334)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_62),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_62),
.Y(n_280)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_64),
.A2(n_118),
.B1(n_120),
.B2(n_122),
.Y(n_117)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

NAND2x1p5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_78),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_78),
.Y(n_245)
);

OA22x2_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_83),
.Y(n_253)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_90),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_96),
.B(n_334),
.Y(n_333)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_105),
.B1(n_117),
.B2(n_123),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g186 ( 
.A1(n_97),
.A2(n_105),
.B1(n_117),
.B2(n_123),
.Y(n_186)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21x1_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_112),
.B(n_117),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_127),
.B(n_174),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_148),
.B2(n_149),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_129),
.B(n_148),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_148),
.A2(n_149),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_149),
.B(n_242),
.C(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_149),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_149),
.B(n_279),
.Y(n_282)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_155),
.B1(n_163),
.B2(n_167),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_150),
.A2(n_202),
.B1(n_321),
.B2(n_328),
.Y(n_320)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_168),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_151),
.B(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_179),
.B(n_181),
.Y(n_178)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_159),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_159),
.Y(n_327)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_167),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.C(n_178),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_175),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_175),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_175),
.A2(n_185),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_175),
.B(n_186),
.C(n_188),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_176),
.A2(n_178),
.B1(n_284),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_176),
.Y(n_299)
);

NOR2x1_ASAP7_75t_L g269 ( 
.A(n_178),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_178),
.Y(n_284)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_202),
.B(n_210),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_183),
.B(n_191),
.C(n_215),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_186),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_215),
.B2(n_216),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_200),
.B1(n_201),
.B2(n_214),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_192),
.B(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_192),
.A2(n_214),
.B1(n_249),
.B2(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_192),
.B(n_201),
.Y(n_335)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_213),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_303),
.B(n_307),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_290),
.B(n_302),
.Y(n_220)
);

OAI21x1_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_246),
.B(n_289),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_241),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_223),
.B(n_241),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_240),
.Y(n_223)
);

XOR2x2_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_233),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_225),
.B(n_233),
.Y(n_293)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_236),
.Y(n_277)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_242),
.A2(n_243),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_242),
.B(n_293),
.C(n_295),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_242),
.A2(n_243),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_244),
.Y(n_266)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_267),
.B(n_288),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_264),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_SL g288 ( 
.A(n_248),
.B(n_264),
.Y(n_288)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_283),
.B(n_287),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_278),
.B(n_282),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_276),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_284),
.B(n_285),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_301),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_301),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_295),
.B1(n_296),
.B2(n_300),
.Y(n_291)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_336),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_315),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_332),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2x1_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);


endmodule