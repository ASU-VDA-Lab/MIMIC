module real_jpeg_13287_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_249;
wire n_286;
wire n_166;
wire n_78;
wire n_176;
wire n_215;
wire n_221;
wire n_292;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_262;
wire n_148;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_213;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx10_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_3),
.A2(n_41),
.B1(n_47),
.B2(n_51),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_3),
.A2(n_41),
.B1(n_66),
.B2(n_67),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_5),
.A2(n_66),
.B1(n_67),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_5),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_47),
.B1(n_51),
.B2(n_88),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_88),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_54),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_7),
.A2(n_47),
.B1(n_51),
.B2(n_54),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_7),
.A2(n_54),
.B1(n_66),
.B2(n_67),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_8),
.A2(n_27),
.B(n_33),
.C(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_8),
.B(n_42),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_8),
.B(n_28),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_8),
.A2(n_28),
.B(n_139),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_8),
.B(n_62),
.C(n_67),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_8),
.A2(n_38),
.B1(n_47),
.B2(n_51),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_8),
.A2(n_82),
.B1(n_83),
.B2(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_8),
.B(n_110),
.Y(n_190)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_56),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_10),
.A2(n_47),
.B1(n_51),
.B2(n_56),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_10),
.A2(n_56),
.B1(n_66),
.B2(n_67),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_56),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_11),
.A2(n_66),
.B1(n_67),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_11),
.A2(n_47),
.B1(n_51),
.B2(n_86),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_86),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_86),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_13),
.A2(n_47),
.B1(n_51),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_13),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_13),
.A2(n_66),
.B1(n_67),
.B2(n_74),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_74),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_74),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_14),
.A2(n_47),
.B1(n_51),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_71),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_14),
.A2(n_66),
.B1(n_67),
.B2(n_71),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_71),
.Y(n_249)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_276),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_254),
.B(n_275),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_227),
.B(n_253),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_122),
.B(n_203),
.C(n_226),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_101),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_21),
.B(n_101),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_77),
.C(n_92),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_22),
.B(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_43),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_23),
.B(n_57),
.C(n_76),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_24),
.B(n_272),
.Y(n_291)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_25),
.A2(n_26),
.B1(n_40),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_25),
.A2(n_26),
.B1(n_105),
.B2(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_25),
.A2(n_220),
.B(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_25),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_26),
.A2(n_290),
.B(n_291),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_28),
.A2(n_29),
.B1(n_49),
.B2(n_50),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_28),
.A2(n_31),
.B(n_38),
.Y(n_91)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_SL g140 ( 
.A(n_29),
.B(n_49),
.C(n_51),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_38),
.B(n_83),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_38),
.B(n_65),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_42),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_42),
.B(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_57),
.B1(n_58),
.B2(n_76),
.Y(n_43)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_53),
.B2(n_55),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_45),
.A2(n_46),
.B1(n_53),
.B2(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_45),
.A2(n_55),
.B(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_45),
.A2(n_46),
.B1(n_100),
.B2(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_45),
.A2(n_109),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_45),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_45),
.A2(n_222),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.Y(n_45)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_46),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g51 ( 
.A(n_47),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_47),
.A2(n_50),
.B(n_138),
.C(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_47),
.B(n_163),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_69),
.B(n_72),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_59),
.A2(n_132),
.B(n_134),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_59),
.A2(n_65),
.B(n_69),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_73),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_60),
.A2(n_75),
.B1(n_133),
.B2(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_60),
.A2(n_75),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_60),
.A2(n_75),
.B1(n_156),
.B2(n_166),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_60),
.A2(n_75),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_60),
.A2(n_213),
.B(n_237),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_66),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_70),
.B(n_75),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_72),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_77),
.A2(n_78),
.B1(n_92),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_89),
.B2(n_90),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_89),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_81),
.A2(n_120),
.B(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_81),
.A2(n_84),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_82),
.A2(n_83),
.B1(n_169),
.B2(n_177),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_82),
.A2(n_171),
.B(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_82),
.A2(n_83),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_96),
.Y(n_120)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_85),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_84),
.B(n_143),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_99),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_95),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_112),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_102),
.B(n_113),
.C(n_121),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_111),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_104),
.B(n_106),
.C(n_111),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_110),
.B(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_110),
.A2(n_246),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_121),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_114),
.B(n_117),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_115),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_116),
.B(n_134),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_201),
.B(n_202),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_144),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_125),
.B(n_128),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.C(n_135),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_135),
.B1(n_136),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_141),
.B1(n_142),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_143),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_157),
.B(n_200),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_149),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_155),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_152),
.A2(n_153),
.B1(n_155),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_194),
.B(n_199),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_183),
.B(n_193),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_172),
.B(n_182),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_167),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_164),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_178),
.B(n_181),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_180),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_185),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_189),
.C(n_192),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_198),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_225),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_225),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_207),
.C(n_215),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_215),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_214),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_218),
.C(n_224),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_224),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_223),
.B(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_229),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_252),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_238),
.B1(n_250),
.B2(n_251),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_251),
.C(n_252),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_232),
.A2(n_233),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_235),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g280 ( 
.A1(n_233),
.A2(n_266),
.B(n_268),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_243),
.C(n_247),
.Y(n_257)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_244),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_274),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_274),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_273),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_259),
.C(n_265),
.Y(n_278)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_265),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_263),
.B(n_264),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_263),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_280),
.CI(n_281),
.CON(n_279),
.SN(n_279)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_293),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_279),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_279),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_289),
.B2(n_292),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_287),
.B2(n_288),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_289),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);


endmodule