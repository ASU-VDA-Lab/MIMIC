module real_jpeg_27326_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_341, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_341;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_0),
.A2(n_27),
.B1(n_31),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_0),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_113),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_0),
.A2(n_53),
.B1(n_54),
.B2(n_113),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_0),
.A2(n_58),
.B1(n_60),
.B2(n_113),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_1),
.Y(n_99)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_1),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_2),
.B(n_26),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_2),
.B(n_31),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_2),
.A2(n_31),
.B(n_161),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_2),
.A2(n_53),
.B1(n_54),
.B2(n_118),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_2),
.A2(n_55),
.B(n_58),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_2),
.B(n_77),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_2),
.A2(n_97),
.B1(n_135),
.B2(n_212),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_3),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_27),
.B1(n_31),
.B2(n_120),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_120),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_3),
.A2(n_58),
.B1(n_60),
.B2(n_120),
.Y(n_212)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_5),
.A2(n_27),
.B1(n_31),
.B2(n_37),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_5),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_5),
.A2(n_37),
.B1(n_58),
.B2(n_60),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_8),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_8),
.A2(n_46),
.B1(n_58),
.B2(n_60),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_8),
.A2(n_27),
.B1(n_31),
.B2(n_46),
.Y(n_269)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_10),
.A2(n_27),
.B1(n_31),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_10),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_115),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_10),
.A2(n_58),
.B1(n_60),
.B2(n_115),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_115),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_11),
.A2(n_48),
.B1(n_58),
.B2(n_60),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_11),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_11),
.A2(n_27),
.B1(n_31),
.B2(n_48),
.Y(n_290)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_13),
.A2(n_27),
.B1(n_31),
.B2(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_14),
.A2(n_25),
.B1(n_53),
.B2(n_54),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_14),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_14),
.A2(n_25),
.B1(n_58),
.B2(n_60),
.Y(n_158)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_15),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_339),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_82),
.B(n_337),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_20),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_21),
.A2(n_44),
.B(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_22),
.A2(n_33),
.B(n_81),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_22),
.A2(n_26),
.B(n_33),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_26),
.B(n_29),
.C(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_29),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g117 ( 
.A(n_23),
.B(n_118),
.CON(n_117),
.SN(n_117)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_26),
.A2(n_33),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_27),
.A2(n_34),
.B1(n_117),
.B2(n_132),
.Y(n_131)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_27),
.A2(n_53),
.A3(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_159)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_29),
.B(n_31),
.Y(n_132)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_32),
.A2(n_45),
.B(n_49),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_33),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_36),
.B(n_49),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_39),
.B(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_74),
.C(n_79),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_40),
.A2(n_41),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_50),
.C(n_63),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_42),
.A2(n_43),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_44),
.A2(n_49),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_44),
.A2(n_49),
.B1(n_126),
.B2(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_50),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_50),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_50),
.A2(n_63),
.B1(n_305),
.B2(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_57),
.B(n_61),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_61),
.B(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_51),
.A2(n_57),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_51),
.A2(n_169),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_51),
.A2(n_57),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_51),
.A2(n_57),
.B1(n_168),
.B2(n_187),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_51),
.A2(n_57),
.B1(n_92),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_51),
.A2(n_108),
.B(n_245),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_54),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g162 ( 
.A(n_54),
.B(n_66),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_54),
.A2(n_56),
.B(n_118),
.C(n_189),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_57),
.B(n_118),
.Y(n_210)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_60),
.B(n_217),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_62),
.B(n_109),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_63),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_64),
.A2(n_76),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_65),
.A2(n_71),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_65),
.A2(n_71),
.B1(n_112),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_65),
.A2(n_71),
.B1(n_144),
.B2(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_65),
.B(n_70),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_65),
.A2(n_71),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_66),
.Y(n_160)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_69),
.A2(n_77),
.B(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_74),
.A2(n_75),
.B1(n_79),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_76),
.A2(n_78),
.B(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_76),
.A2(n_255),
.B(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_79),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_330),
.B(n_336),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_300),
.A3(n_322),
.B1(n_328),
.B2(n_329),
.C(n_341),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_281),
.B(n_299),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_259),
.B(n_280),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_150),
.B(n_236),
.C(n_258),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_136),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_88),
.B(n_136),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_121),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_105),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_90),
.B(n_105),
.C(n_121),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_91),
.B(n_96),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_93),
.B(n_179),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_100),
.B(n_101),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_97),
.A2(n_100),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_97),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_97),
.A2(n_204),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_97),
.A2(n_103),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_98),
.A2(n_102),
.B(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_98),
.A2(n_199),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_103),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_103),
.B(n_118),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_116),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_119),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_130),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_123),
.B(n_128),
.C(n_130),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_133),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_135),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_137),
.A2(n_138),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_142),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_147),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_148),
.B(n_198),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_235),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_228),
.B(n_234),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_180),
.B(n_227),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_170),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_154),
.B(n_170),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_163),
.C(n_166),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_155),
.A2(n_156),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_158),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_171),
.B(n_177),
.C(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_221),
.B(n_226),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_200),
.B(n_220),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_183),
.B(n_190),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_195),
.C(n_196),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

INVx11_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_208),
.B(n_219),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_206),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_214),
.B(n_218),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_210),
.B(n_211),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_223),
.Y(n_226)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_229),
.B(n_230),
.Y(n_234)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_237),
.B(n_238),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_256),
.B2(n_257),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_246),
.B2(n_247),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_247),
.C(n_257),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_250),
.C(n_254),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_261),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_279),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_272),
.B2(n_273),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_273),
.C(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_268),
.C(n_270),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_269),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_277),
.B2(n_278),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_275),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_277),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_275),
.A2(n_293),
.B(n_296),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_277),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_283),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_297),
.B2(n_298),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_292),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_292),
.C(n_298),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B(n_291),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_290),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_302),
.C(n_312),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_291),
.A2(n_302),
.B1(n_303),
.B2(n_327),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_291),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_297),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_314),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_314),
.Y(n_329)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_307),
.C(n_309),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_309),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_311),
.B1(n_316),
.B2(n_320),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_320),
.C(n_321),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_313),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_321),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_333),
.Y(n_335)
);


endmodule