module fake_jpeg_14652_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_0),
.B(n_31),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_58),
.Y(n_70)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_79),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_55),
.B1(n_46),
.B2(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_81),
.B1(n_75),
.B2(n_80),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_49),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_57),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_55),
.B1(n_45),
.B2(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_52),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_1),
.B(n_2),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_44),
.B1(n_54),
.B2(n_50),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_108)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_91),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_53),
.B1(n_48),
.B2(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_90),
.B1(n_96),
.B2(n_98),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_53),
.B1(n_23),
.B2(n_25),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_78),
.C(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_99),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_21),
.B1(n_39),
.B2(n_38),
.Y(n_98)
);

BUFx2_ASAP7_75t_SL g99 ( 
.A(n_78),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_5),
.Y(n_105)
);

OAI32xp33_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_19),
.A3(n_36),
.B1(n_35),
.B2(n_34),
.Y(n_101)
);

OR2x4_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_111),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_108),
.B(n_9),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_18),
.B1(n_33),
.B2(n_32),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_93),
.B1(n_96),
.B2(n_87),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_109),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_114),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_103),
.B(n_86),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_117),
.B(n_97),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_104),
.C(n_107),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_108),
.C(n_111),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_113),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_122),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_102),
.B(n_110),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_121),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_126),
.Y(n_131)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_106),
.C(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_130),
.Y(n_134)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_131),
.CI(n_129),
.CON(n_135),
.SN(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_127),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_135),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_133),
.B1(n_126),
.B2(n_12),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

OAI21x1_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_27),
.B(n_11),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_94),
.B1(n_92),
.B2(n_16),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_29),
.C(n_15),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_26),
.Y(n_143)
);


endmodule