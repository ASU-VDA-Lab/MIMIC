module real_jpeg_2407_n_19 (n_17, n_108, n_8, n_116, n_0, n_111, n_2, n_10, n_114, n_9, n_12, n_6, n_11, n_14, n_110, n_112, n_7, n_117, n_18, n_3, n_5, n_4, n_109, n_115, n_1, n_118, n_16, n_15, n_13, n_113, n_19);

input n_17;
input n_108;
input n_8;
input n_116;
input n_0;
input n_111;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_110;
input n_112;
input n_7;
input n_117;
input n_18;
input n_3;
input n_5;
input n_4;
input n_109;
input n_115;
input n_1;
input n_118;
input n_16;
input n_15;
input n_13;
input n_113;

output n_19;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx1_ASAP7_75t_L g91 ( 
.A(n_0),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_3),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_5),
.A2(n_21),
.B1(n_22),
.B2(n_27),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_7),
.B(n_48),
.C(n_63),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_9),
.A2(n_49),
.B1(n_51),
.B2(n_62),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_10),
.B(n_40),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_12),
.B(n_46),
.C(n_70),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_13),
.A2(n_44),
.B1(n_76),
.B2(n_79),
.Y(n_43)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_14),
.B(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_14),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_15),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_16),
.B(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_16),
.Y(n_98)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_18),
.A2(n_53),
.B(n_57),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_28),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_24),
.B(n_94),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_26),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_36),
.B(n_105),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_31),
.B(n_35),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_34),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_34),
.B(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI221xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B1(n_43),
.B2(n_81),
.C(n_95),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_72),
.C(n_73),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_65),
.C(n_66),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_60),
.C(n_61),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_60),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_90),
.Y(n_81)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_96),
.A3(n_97),
.B1(n_100),
.B2(n_101),
.C1(n_104),
.C2(n_118),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_84),
.C(n_87),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_108),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_109),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_110),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_111),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_112),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_113),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_114),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_115),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_116),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_117),
.Y(n_94)
);


endmodule