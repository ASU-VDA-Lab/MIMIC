module real_jpeg_28079_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_216;
wire n_128;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_0),
.A2(n_27),
.B1(n_30),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_0),
.A2(n_44),
.B1(n_81),
.B2(n_82),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_0),
.A2(n_33),
.B1(n_37),
.B2(n_44),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_0),
.A2(n_44),
.B1(n_50),
.B2(n_51),
.Y(n_102)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_1),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_81),
.B1(n_82),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_2),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_107),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_107),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_2),
.A2(n_33),
.B1(n_37),
.B2(n_107),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_3),
.A2(n_81),
.B1(n_82),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_3),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_152),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_3),
.A2(n_27),
.B1(n_30),
.B2(n_152),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_3),
.A2(n_33),
.B1(n_37),
.B2(n_152),
.Y(n_237)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_4),
.Y(n_80)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_5),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_5),
.B(n_84),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_5),
.B(n_50),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_5),
.A2(n_50),
.B(n_189),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_5),
.A2(n_27),
.B1(n_30),
.B2(n_150),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_5),
.A2(n_33),
.B(n_38),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_5),
.B(n_100),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_5),
.A2(n_65),
.B1(n_237),
.B2(n_238),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_7),
.A2(n_81),
.B1(n_82),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_7),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_132),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_7),
.A2(n_27),
.B1(n_30),
.B2(n_132),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_7),
.A2(n_33),
.B1(n_37),
.B2(n_132),
.Y(n_229)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_8),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_58),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_9),
.A2(n_33),
.B1(n_37),
.B2(n_58),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_10),
.A2(n_29),
.B1(n_33),
.B2(n_37),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_10),
.A2(n_29),
.B1(n_81),
.B2(n_82),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_10),
.A2(n_29),
.B1(n_50),
.B2(n_51),
.Y(n_127)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_36),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_12),
.A2(n_27),
.B1(n_30),
.B2(n_60),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_12),
.A2(n_33),
.B1(n_37),
.B2(n_60),
.Y(n_120)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_15),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_134),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_110),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_20),
.B(n_110),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_90),
.B2(n_109),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_62),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_45),
.B(n_61),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_24),
.B(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_25),
.A2(n_41),
.B(n_197),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_26),
.Y(n_143)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_27),
.A2(n_30),
.B1(n_49),
.B2(n_55),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_27),
.B(n_48),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_27),
.A2(n_36),
.B(n_150),
.C(n_216),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g187 ( 
.A1(n_30),
.A2(n_51),
.A3(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_31),
.B(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_32),
.A2(n_41),
.B1(n_73),
.B2(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_32),
.A2(n_39),
.B(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_32),
.A2(n_41),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_32),
.A2(n_41),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_32),
.A2(n_41),
.B1(n_196),
.B2(n_214),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_32),
.B(n_150),
.Y(n_235)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_37),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_73),
.B(n_74),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_41),
.A2(n_74),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_46),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_46),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_46),
.A2(n_54),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_46),
.A2(n_54),
.B1(n_146),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_46),
.A2(n_54),
.B1(n_175),
.B2(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_54),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_47)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_48),
.Y(n_188)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_51),
.B1(n_79),
.B2(n_80),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_50),
.B(n_79),
.Y(n_164)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_51),
.A2(n_83),
.B1(n_149),
.B2(n_164),
.Y(n_163)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_54),
.B(n_102),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_54),
.B(n_127),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_75),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_72),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_76),
.B1(n_77),
.B2(n_89),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_64),
.A2(n_72),
.B1(n_89),
.B2(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B(n_70),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_65),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_65),
.A2(n_68),
.B1(n_120),
.B2(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_65),
.A2(n_96),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_65),
.A2(n_229),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_94),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_66),
.A2(n_71),
.B(n_122),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_66),
.A2(n_67),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_71),
.Y(n_96)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_95),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_68),
.A2(n_93),
.B(n_166),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_72),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_85),
.B(n_86),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_78),
.A2(n_84),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B(n_83),
.C(n_84),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_81),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

HAxp5_ASAP7_75t_SL g149 ( 
.A(n_81),
.B(n_150),
.CON(n_149),
.SN(n_149)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_105),
.B1(n_106),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_87),
.A2(n_105),
.B1(n_131),
.B2(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_99),
.C(n_103),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_92),
.B(n_97),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_108),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_117),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_115),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_117),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.C(n_129),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_118),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_123),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_124),
.A2(n_129),
.B1(n_130),
.B2(n_271),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_124),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_128),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_160),
.B(n_161),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_275),
.B(n_280),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_179),
.B(n_261),
.C(n_274),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_167),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_137),
.B(n_167),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_153),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_139),
.B(n_140),
.C(n_153),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_148),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_150),
.B(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_162),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_155),
.B(n_159),
.C(n_162),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_165),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.C(n_173),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_168),
.A2(n_169),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_173),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_178),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_178),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_260),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_253),
.B(n_259),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_207),
.B(n_252),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_198),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_183),
.B(n_198),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_191),
.C(n_194),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_184),
.A2(n_185),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_187),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_199),
.B(n_205),
.C(n_206),
.Y(n_254)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_246),
.B(n_251),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_225),
.B(n_245),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_217),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_210),
.B(n_217),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_232),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_215),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_222),
.C(n_223),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_224),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_233),
.B(n_244),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_227),
.B(n_231),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_239),
.B(n_243),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_236),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_254),
.B(n_255),
.Y(n_259)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_262),
.B(n_263),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_272),
.B2(n_273),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_269),
.C(n_273),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);


endmodule