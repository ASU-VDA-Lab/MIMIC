module real_jpeg_29983_n_18 (n_17, n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_0),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_0),
.A2(n_45),
.B1(n_54),
.B2(n_55),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_1),
.Y(n_85)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_2),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_105),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_105),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_2),
.A2(n_48),
.B1(n_50),
.B2(n_105),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_3),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_28),
.B(n_32),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_115),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_3),
.B(n_30),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_3),
.A2(n_54),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_3),
.B(n_54),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_3),
.B(n_66),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_3),
.A2(n_83),
.B1(n_240),
.B2(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_3),
.A2(n_31),
.B(n_256),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_5),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_111),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_111),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_5),
.A2(n_48),
.B1(n_50),
.B2(n_111),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_6),
.A2(n_43),
.B1(n_54),
.B2(n_55),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_6),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_36),
.B1(n_54),
.B2(n_55),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_8),
.A2(n_36),
.B1(n_48),
.B2(n_50),
.Y(n_125)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_10),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_95),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_95),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_10),
.A2(n_48),
.B1(n_50),
.B2(n_95),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

OAI32xp33_ASAP7_75t_L g216 ( 
.A1(n_11),
.A2(n_50),
.A3(n_54),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_12),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_102),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_12),
.A2(n_48),
.B1(n_50),
.B2(n_102),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_102),
.Y(n_260)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_14),
.B(n_31),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_61),
.Y(n_63)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_14),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_15),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_15),
.A2(n_26),
.B1(n_48),
.B2(n_50),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_15),
.A2(n_26),
.B1(n_54),
.B2(n_55),
.Y(n_136)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_16),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_17),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g177 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_100),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_17),
.A2(n_54),
.B1(n_55),
.B2(n_100),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_17),
.A2(n_48),
.B1(n_50),
.B2(n_100),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_332),
.B(n_335),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_74),
.B(n_331),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_21),
.B(n_37),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_21),
.B(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_21),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_23),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_25),
.A2(n_34),
.B(n_115),
.C(n_116),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_30),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_27),
.A2(n_30),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_27),
.A2(n_30),
.B1(n_101),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_27),
.A2(n_30),
.B1(n_110),
.B2(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_27),
.A2(n_30),
.B(n_35),
.Y(n_334)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_31),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

OAI32xp33_ASAP7_75t_L g264 ( 
.A1(n_31),
.A2(n_55),
.A3(n_257),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_32),
.B(n_115),
.Y(n_257)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_67),
.C(n_69),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_38),
.A2(n_39),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_57),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_40),
.B(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_42),
.A2(n_71),
.B1(n_73),
.B2(n_163),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_46),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_46),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_46),
.A2(n_57),
.B1(n_309),
.B2(n_316),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_52),
.B(n_56),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_47),
.A2(n_52),
.B1(n_93),
.B2(n_96),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_47),
.A2(n_52),
.B1(n_96),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_47),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_47),
.A2(n_52),
.B1(n_56),
.B2(n_136),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_47),
.A2(n_52),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_47),
.A2(n_52),
.B1(n_214),
.B2(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_47),
.B(n_115),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_47),
.A2(n_52),
.B1(n_181),
.B2(n_284),
.Y(n_283)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_48),
.B(n_51),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_48),
.B(n_246),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_52),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_54),
.B(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_57),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_58),
.A2(n_66),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_58),
.A2(n_66),
.B1(n_106),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_58),
.A2(n_66),
.B1(n_177),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_58),
.A2(n_64),
.B1(n_66),
.B2(n_307),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_63),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_59),
.A2(n_63),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_59),
.A2(n_63),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_59),
.A2(n_63),
.B1(n_121),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_59),
.A2(n_63),
.B1(n_189),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_329),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_67),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_73),
.B1(n_109),
.B2(n_112),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_71),
.A2(n_73),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_324),
.B(n_330),
.Y(n_74)
);

OAI321xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_300),
.A3(n_319),
.B1(n_322),
.B2(n_323),
.C(n_341),
.Y(n_75)
);

AOI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_147),
.A3(n_169),
.B1(n_294),
.B2(n_299),
.C(n_342),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_78),
.A2(n_295),
.B(n_298),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_128),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_79),
.B(n_128),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_107),
.C(n_123),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_80),
.B(n_123),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_97),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_81),
.B(n_98),
.C(n_103),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_92),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_82),
.B(n_92),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_88),
.B2(n_91),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_90),
.B1(n_91),
.B2(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_83),
.A2(n_88),
.B(n_125),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_83),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_83),
.A2(n_90),
.B1(n_234),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_83),
.A2(n_228),
.B1(n_229),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_87),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_84),
.A2(n_89),
.B1(n_118),
.B2(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_84),
.A2(n_89),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g229 ( 
.A(n_89),
.Y(n_229)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_94),
.A2(n_134),
.B1(n_137),
.B2(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_104),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_107),
.B(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.C(n_120),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_108),
.B(n_120),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_113),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_114),
.B(n_117),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_115),
.B(n_244),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_126),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_127),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_146),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_140),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_140),
.C(n_146),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_138),
.B2(n_139),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_134),
.A2(n_137),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_139),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_138),
.A2(n_161),
.B(n_164),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_140),
.Y(n_340)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_143),
.CI(n_145),
.CON(n_140),
.SN(n_140)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_143),
.C(n_145),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_148),
.B(n_149),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_167),
.B2(n_168),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_158),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_152),
.B(n_158),
.C(n_168),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_156),
.B(n_157),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_156),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_155),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_157),
.B(n_302),
.C(n_311),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g321 ( 
.A(n_157),
.B(n_302),
.CI(n_311),
.CON(n_321),
.SN(n_321)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_167),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_199),
.C(n_204),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_193),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_171),
.B(n_193),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_184),
.C(n_185),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_172),
.B(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_182),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_179),
.C(n_182),
.Y(n_196)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_292),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_184),
.Y(n_292)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_187),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_190),
.B(n_192),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_191),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_196),
.C(n_197),
.Y(n_201)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_200),
.A2(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_201),
.B(n_202),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_288),
.B(n_293),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_274),
.B(n_287),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_250),
.B(n_273),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_230),
.B(n_249),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_219),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_209),
.B(n_219),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_210),
.A2(n_211),
.B1(n_215),
.B2(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_213),
.Y(n_217)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_226),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_224),
.C(n_226),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_225),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_227),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_237),
.B(n_248),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_236),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_242),
.B(n_247),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_241),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_252),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_263),
.B1(n_271),
.B2(n_272),
.Y(n_252)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_258),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_262),
.C(n_272),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_260),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_263),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_269),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_269),
.Y(n_282)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_275),
.B(n_276),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_283),
.C(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_312),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_312),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_310),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_304),
.B1(n_314),
.B2(n_317),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_306),
.C(n_309),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_317),
.C(n_318),
.Y(n_325)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_318),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_321),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_321),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_334),
.B(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_336),
.Y(n_335)
);


endmodule