module real_aes_8949_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_182;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g189 ( .A1(n_0), .A2(n_190), .B(n_191), .C(n_195), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_1), .B(n_185), .Y(n_196) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_3), .B(n_150), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_4), .A2(n_131), .B(n_480), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_5), .A2(n_136), .B(n_141), .C(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_6), .A2(n_131), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_7), .B(n_185), .Y(n_486) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_8), .A2(n_164), .B(n_214), .Y(n_213) );
AND2x6_ASAP7_75t_L g136 ( .A(n_9), .B(n_137), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_10), .A2(n_136), .B(n_141), .C(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g541 ( .A(n_11), .Y(n_541) );
INVx1_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_12), .B(n_39), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_13), .B(n_194), .Y(n_518) );
INVx1_ASAP7_75t_L g160 ( .A(n_14), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_15), .B(n_150), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_16), .A2(n_151), .B(n_526), .C(n_528), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_17), .B(n_185), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_18), .B(n_178), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_19), .A2(n_141), .B(n_172), .C(n_177), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_20), .A2(n_193), .B(n_208), .C(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_21), .B(n_194), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_22), .A2(n_76), .B1(n_735), .B2(n_736), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_22), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_23), .B(n_194), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_24), .Y(n_467) );
INVx1_ASAP7_75t_L g492 ( .A(n_25), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_26), .A2(n_141), .B(n_177), .C(n_217), .Y(n_216) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_27), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_28), .Y(n_514) );
INVx1_ASAP7_75t_L g568 ( .A(n_29), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_30), .A2(n_131), .B(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g134 ( .A(n_31), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_32), .A2(n_139), .B(n_144), .C(n_154), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_33), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_34), .A2(n_193), .B(n_483), .C(n_485), .Y(n_482) );
INVxp67_ASAP7_75t_L g569 ( .A(n_35), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_36), .B(n_219), .Y(n_218) );
CKINVDCx14_ASAP7_75t_R g481 ( .A(n_37), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_38), .A2(n_141), .B(n_177), .C(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_39), .B(n_107), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_40), .A2(n_195), .B(n_539), .C(n_540), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_41), .B(n_170), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_42), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_43), .B(n_150), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_44), .B(n_131), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_45), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_46), .Y(n_565) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_47), .A2(n_139), .B(n_154), .C(n_228), .Y(n_227) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_48), .A2(n_87), .B1(n_121), .B2(n_122), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_48), .Y(n_122) );
INVx1_ASAP7_75t_L g192 ( .A(n_49), .Y(n_192) );
INVx1_ASAP7_75t_L g229 ( .A(n_50), .Y(n_229) );
INVx1_ASAP7_75t_L g504 ( .A(n_51), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_52), .B(n_131), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_53), .Y(n_181) );
CKINVDCx14_ASAP7_75t_R g537 ( .A(n_54), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_55), .Y(n_448) );
INVx1_ASAP7_75t_L g137 ( .A(n_56), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_57), .B(n_131), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_58), .B(n_185), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_59), .A2(n_176), .B(n_239), .C(n_241), .Y(n_238) );
INVx1_ASAP7_75t_L g159 ( .A(n_60), .Y(n_159) );
INVx1_ASAP7_75t_SL g484 ( .A(n_61), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_62), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_63), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_64), .B(n_185), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_65), .B(n_151), .Y(n_205) );
INVx1_ASAP7_75t_L g470 ( .A(n_66), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g188 ( .A(n_67), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_68), .B(n_147), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_69), .A2(n_102), .B1(n_113), .B2(n_747), .Y(n_101) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_70), .A2(n_141), .B(n_154), .C(n_265), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_71), .Y(n_237) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_73), .A2(n_131), .B(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_74), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_75), .A2(n_131), .B(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_76), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_77), .A2(n_170), .B(n_564), .Y(n_563) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_78), .Y(n_489) );
INVx1_ASAP7_75t_L g524 ( .A(n_79), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_80), .B(n_146), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_81), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_82), .A2(n_131), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g527 ( .A(n_83), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_84), .Y(n_746) );
INVx2_ASAP7_75t_L g157 ( .A(n_85), .Y(n_157) );
INVx1_ASAP7_75t_L g517 ( .A(n_86), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_87), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_88), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_89), .B(n_194), .Y(n_206) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_90), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g443 ( .A(n_90), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g453 ( .A(n_90), .B(n_445), .Y(n_453) );
INVx2_ASAP7_75t_L g457 ( .A(n_90), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_91), .A2(n_141), .B(n_154), .C(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_92), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g145 ( .A(n_93), .Y(n_145) );
INVxp67_ASAP7_75t_L g242 ( .A(n_94), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_95), .B(n_164), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_96), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g201 ( .A(n_97), .Y(n_201) );
INVx1_ASAP7_75t_L g266 ( .A(n_98), .Y(n_266) );
INVx2_ASAP7_75t_L g507 ( .A(n_99), .Y(n_507) );
AND2x2_ASAP7_75t_L g231 ( .A(n_100), .B(n_156), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx5_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_105), .Y(n_748) );
OR2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
AND2x2_ASAP7_75t_L g445 ( .A(n_109), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OAI21x1_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_118), .B(n_449), .Y(n_113) );
OAI21xp5_ASAP7_75t_SL g449 ( .A1(n_114), .A2(n_447), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_441), .B(n_447), .Y(n_118) );
XOR2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
INVx2_ASAP7_75t_L g454 ( .A(n_123), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_123), .A2(n_738), .B1(n_741), .B2(n_742), .Y(n_737) );
OR3x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_355), .C(n_398), .Y(n_123) );
NAND5xp2_ASAP7_75t_L g124 ( .A(n_125), .B(n_282), .C(n_312), .D(n_329), .E(n_344), .Y(n_124) );
AOI221xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_197), .B1(n_244), .B2(n_250), .C(n_254), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_166), .Y(n_126) );
OR2x2_ASAP7_75t_L g259 ( .A(n_127), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g299 ( .A(n_127), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g317 ( .A(n_127), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_127), .B(n_252), .Y(n_334) );
OR2x2_ASAP7_75t_L g346 ( .A(n_127), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_127), .B(n_305), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_127), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_127), .B(n_283), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_127), .B(n_291), .Y(n_397) );
AND2x2_ASAP7_75t_L g429 ( .A(n_127), .B(n_183), .Y(n_429) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_127), .Y(n_437) );
INVx5_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_128), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g256 ( .A(n_128), .B(n_232), .Y(n_256) );
BUFx2_ASAP7_75t_L g279 ( .A(n_128), .Y(n_279) );
AND2x2_ASAP7_75t_L g308 ( .A(n_128), .B(n_167), .Y(n_308) );
AND2x2_ASAP7_75t_L g363 ( .A(n_128), .B(n_260), .Y(n_363) );
OR2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_161), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_138), .B(n_156), .Y(n_129) );
BUFx2_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
NAND2x1p5_ASAP7_75t_L g202 ( .A(n_132), .B(n_136), .Y(n_202) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g142 ( .A(n_134), .Y(n_142) );
INVx1_ASAP7_75t_L g209 ( .A(n_134), .Y(n_209) );
INVx1_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
INVx3_ASAP7_75t_L g151 ( .A(n_135), .Y(n_151) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_135), .Y(n_194) );
INVx1_ASAP7_75t_L g219 ( .A(n_135), .Y(n_219) );
INVx4_ASAP7_75t_SL g155 ( .A(n_136), .Y(n_155) );
BUFx3_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_SL g187 ( .A1(n_140), .A2(n_155), .B(n_188), .C(n_189), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_140), .A2(n_155), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_140), .A2(n_155), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g503 ( .A1(n_140), .A2(n_155), .B(n_504), .C(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g523 ( .A1(n_140), .A2(n_155), .B(n_524), .C(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_SL g536 ( .A1(n_140), .A2(n_155), .B(n_537), .C(n_538), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_SL g564 ( .A1(n_140), .A2(n_155), .B(n_565), .C(n_566), .Y(n_564) );
INVx5_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx3_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_142), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_149), .C(n_152), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_146), .A2(n_152), .B(n_229), .C(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_146), .A2(n_470), .B(n_471), .C(n_472), .Y(n_469) );
O2A1O1Ixp5_ASAP7_75t_L g516 ( .A1(n_146), .A2(n_472), .B(n_517), .C(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx4_ASAP7_75t_L g240 ( .A(n_148), .Y(n_240) );
INVx2_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_150), .B(n_242), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_150), .A2(n_175), .B(n_492), .C(n_493), .Y(n_491) );
OAI22xp33_ASAP7_75t_L g567 ( .A1(n_150), .A2(n_240), .B1(n_568), .B2(n_569), .Y(n_567) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_151), .B(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
INVx1_ASAP7_75t_L g528 ( .A(n_153), .Y(n_528) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
INVx1_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_156), .A2(n_226), .B(n_227), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_156), .A2(n_202), .B(n_489), .C(n_490), .Y(n_488) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_156), .A2(n_535), .B(n_542), .Y(n_534) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_157), .B(n_158), .Y(n_156) );
AND2x2_ASAP7_75t_L g165 ( .A(n_157), .B(n_158), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
INVx3_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_163), .A2(n_200), .B(n_210), .Y(n_199) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_163), .A2(n_263), .B(n_271), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_163), .B(n_272), .Y(n_271) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_163), .A2(n_466), .B(n_473), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_163), .B(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_163), .B(n_520), .Y(n_519) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_164), .A2(n_215), .B(n_216), .Y(n_214) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_164), .Y(n_234) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_166), .B(n_317), .Y(n_326) );
OAI32xp33_ASAP7_75t_L g340 ( .A1(n_166), .A2(n_276), .A3(n_341), .B1(n_342), .B2(n_343), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_166), .B(n_342), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_166), .B(n_259), .Y(n_383) );
INVx1_ASAP7_75t_SL g412 ( .A(n_166), .Y(n_412) );
NAND4xp25_ASAP7_75t_L g421 ( .A(n_166), .B(n_199), .C(n_363), .D(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_183), .Y(n_166) );
INVx5_ASAP7_75t_L g253 ( .A(n_167), .Y(n_253) );
AND2x2_ASAP7_75t_L g283 ( .A(n_167), .B(n_184), .Y(n_283) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_167), .Y(n_362) );
AND2x2_ASAP7_75t_L g432 ( .A(n_167), .B(n_379), .Y(n_432) );
OR2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_180), .Y(n_167) );
AOI21xp5_ASAP7_75t_SL g168 ( .A1(n_169), .A2(n_171), .B(n_178), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_175), .Y(n_172) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_176), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_179), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_182), .A2(n_513), .B(n_519), .Y(n_512) );
AND2x4_ASAP7_75t_L g305 ( .A(n_183), .B(n_253), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_183), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g339 ( .A(n_183), .B(n_260), .Y(n_339) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g252 ( .A(n_184), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g291 ( .A(n_184), .B(n_262), .Y(n_291) );
AND2x2_ASAP7_75t_L g300 ( .A(n_184), .B(n_261), .Y(n_300) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_196), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_193), .B(n_484), .Y(n_483) );
INVx4_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g539 ( .A(n_194), .Y(n_539) );
INVx2_ASAP7_75t_L g472 ( .A(n_195), .Y(n_472) );
AOI222xp33_ASAP7_75t_L g368 ( .A1(n_197), .A2(n_369), .B1(n_371), .B2(n_373), .C1(n_376), .C2(n_377), .Y(n_368) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_221), .Y(n_197) );
AND2x2_ASAP7_75t_L g301 ( .A(n_198), .B(n_302), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g418 ( .A(n_198), .B(n_279), .C(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_213), .Y(n_198) );
INVx5_ASAP7_75t_SL g249 ( .A(n_199), .Y(n_249) );
OAI322xp33_ASAP7_75t_L g254 ( .A1(n_199), .A2(n_255), .A3(n_257), .B1(n_258), .B2(n_273), .C1(n_276), .C2(n_278), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_199), .B(n_247), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_199), .B(n_233), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_203), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_202), .A2(n_467), .B(n_468), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_202), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_207), .A2(n_218), .B(n_220), .Y(n_217) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
INVx2_ASAP7_75t_L g562 ( .A(n_212), .Y(n_562) );
INVx2_ASAP7_75t_L g247 ( .A(n_213), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_213), .B(n_223), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_221), .B(n_286), .Y(n_341) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g320 ( .A(n_222), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_232), .Y(n_222) );
OR2x2_ASAP7_75t_L g248 ( .A(n_223), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_223), .B(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g288 ( .A(n_223), .B(n_233), .Y(n_288) );
AND2x2_ASAP7_75t_L g311 ( .A(n_223), .B(n_247), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_223), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g327 ( .A(n_223), .B(n_286), .Y(n_327) );
AND2x2_ASAP7_75t_L g335 ( .A(n_223), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_223), .B(n_295), .Y(n_385) );
INVx5_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g275 ( .A(n_224), .B(n_249), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_224), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g302 ( .A(n_224), .B(n_233), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_224), .B(n_349), .Y(n_390) );
OR2x2_ASAP7_75t_L g406 ( .A(n_224), .B(n_350), .Y(n_406) );
AND2x2_ASAP7_75t_SL g413 ( .A(n_224), .B(n_367), .Y(n_413) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_224), .Y(n_420) );
OR2x6_ASAP7_75t_L g224 ( .A(n_225), .B(n_231), .Y(n_224) );
AND2x2_ASAP7_75t_L g274 ( .A(n_232), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g324 ( .A(n_232), .B(n_247), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_232), .B(n_249), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_232), .B(n_286), .Y(n_408) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_233), .B(n_249), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_233), .B(n_247), .Y(n_296) );
OR2x2_ASAP7_75t_L g350 ( .A(n_233), .B(n_247), .Y(n_350) );
AND2x2_ASAP7_75t_L g367 ( .A(n_233), .B(n_246), .Y(n_367) );
INVxp67_ASAP7_75t_L g389 ( .A(n_233), .Y(n_389) );
AND2x2_ASAP7_75t_L g416 ( .A(n_233), .B(n_286), .Y(n_416) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_233), .Y(n_423) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_243), .Y(n_233) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_234), .A2(n_479), .B(n_486), .Y(n_478) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_234), .A2(n_502), .B(n_508), .Y(n_501) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_234), .A2(n_522), .B(n_529), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_239), .A2(n_266), .B(n_267), .C(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_240), .B(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_240), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_246), .B(n_297), .Y(n_370) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g286 ( .A(n_247), .B(n_249), .Y(n_286) );
OR2x2_ASAP7_75t_L g353 ( .A(n_247), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g297 ( .A(n_248), .Y(n_297) );
OR2x2_ASAP7_75t_L g358 ( .A(n_248), .B(n_350), .Y(n_358) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g257 ( .A(n_252), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_252), .B(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g258 ( .A(n_253), .B(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_253), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_253), .B(n_260), .Y(n_293) );
INVx2_ASAP7_75t_L g338 ( .A(n_253), .Y(n_338) );
AND2x2_ASAP7_75t_L g351 ( .A(n_253), .B(n_291), .Y(n_351) );
AND2x2_ASAP7_75t_L g376 ( .A(n_253), .B(n_300), .Y(n_376) );
INVx1_ASAP7_75t_L g328 ( .A(n_258), .Y(n_328) );
INVx2_ASAP7_75t_SL g315 ( .A(n_259), .Y(n_315) );
INVx1_ASAP7_75t_L g318 ( .A(n_260), .Y(n_318) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_261), .Y(n_281) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx2_ASAP7_75t_L g379 ( .A(n_262), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_270), .Y(n_263) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g485 ( .A(n_269), .Y(n_485) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g348 ( .A(n_275), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g354 ( .A(n_275), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_275), .A2(n_357), .B1(n_359), .B2(n_364), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_275), .B(n_367), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_276), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g310 ( .A(n_277), .Y(n_310) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
OR2x2_ASAP7_75t_L g292 ( .A(n_279), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_279), .B(n_283), .Y(n_343) );
AND2x2_ASAP7_75t_L g366 ( .A(n_279), .B(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g342 ( .A(n_281), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B(n_289), .C(n_303), .Y(n_282) );
INVx1_ASAP7_75t_L g306 ( .A(n_283), .Y(n_306) );
OAI221xp5_ASAP7_75t_SL g414 ( .A1(n_283), .A2(n_415), .B1(n_417), .B2(n_418), .C(n_421), .Y(n_414) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g433 ( .A(n_286), .Y(n_433) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g382 ( .A(n_288), .B(n_321), .Y(n_382) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_292), .B(n_294), .C(n_298), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OAI32xp33_ASAP7_75t_L g407 ( .A1(n_296), .A2(n_297), .A3(n_360), .B1(n_397), .B2(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x2_ASAP7_75t_L g439 ( .A(n_299), .B(n_338), .Y(n_439) );
AND2x2_ASAP7_75t_L g386 ( .A(n_300), .B(n_338), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_300), .B(n_308), .Y(n_404) );
AOI31xp33_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_306), .A3(n_307), .B(n_309), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_305), .B(n_317), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_305), .B(n_315), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_305), .A2(n_335), .B1(n_425), .B2(n_428), .C(n_430), .Y(n_424) );
CKINVDCx16_ASAP7_75t_R g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g330 ( .A(n_310), .B(n_331), .Y(n_330) );
AOI222xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_319), .B1(n_322), .B2(n_325), .C1(n_327), .C2(n_328), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g395 ( .A(n_314), .Y(n_395) );
INVx1_ASAP7_75t_L g417 ( .A(n_317), .Y(n_417) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_320), .A2(n_431), .B1(n_433), .B2(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g336 ( .A(n_321), .Y(n_336) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B1(n_335), .B2(n_337), .C(n_340), .Y(n_329) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g374 ( .A(n_332), .B(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g426 ( .A(n_332), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g401 ( .A(n_337), .Y(n_401) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g365 ( .A(n_338), .Y(n_365) );
INVx1_ASAP7_75t_L g347 ( .A(n_339), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_342), .B(n_429), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_348), .B1(n_351), .B2(n_352), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g438 ( .A(n_351), .Y(n_438) );
INVxp33_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_353), .B(n_397), .Y(n_396) );
OAI32xp33_ASAP7_75t_L g387 ( .A1(n_354), .A2(n_388), .A3(n_389), .B1(n_390), .B2(n_391), .Y(n_387) );
NAND4xp25_ASAP7_75t_L g355 ( .A(n_356), .B(n_368), .C(n_380), .D(n_392), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
NAND2xp33_ASAP7_75t_SL g359 ( .A(n_360), .B(n_361), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_363), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
CKINVDCx16_ASAP7_75t_R g373 ( .A(n_374), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_377), .A2(n_393), .B1(n_410), .B2(n_413), .C(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g428 ( .A(n_379), .B(n_429), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B1(n_384), .B2(n_386), .C(n_387), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_389), .B(n_420), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B(n_396), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND4xp25_ASAP7_75t_L g398 ( .A(n_399), .B(n_409), .C(n_424), .D(n_435), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_403), .B(n_405), .C(n_407), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g440 ( .A(n_427), .Y(n_440) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .B(n_440), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
NOR2xp33_ASAP7_75t_SL g447 ( .A(n_443), .B(n_448), .Y(n_447) );
NOR2x2_ASAP7_75t_L g745 ( .A(n_444), .B(n_457), .Y(n_745) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g456 ( .A(n_445), .B(n_457), .Y(n_456) );
OAI222xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_734), .B1(n_737), .B2(n_743), .C1(n_744), .C2(n_746), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_454), .B1(n_455), .B2(n_458), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g740 ( .A(n_453), .Y(n_740) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx6_ASAP7_75t_L g741 ( .A(n_456), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_458), .Y(n_742) );
AND2x2_ASAP7_75t_SL g458 ( .A(n_459), .B(n_689), .Y(n_458) );
NOR4xp25_ASAP7_75t_L g459 ( .A(n_460), .B(n_626), .C(n_660), .D(n_676), .Y(n_459) );
NAND4xp25_ASAP7_75t_SL g460 ( .A(n_461), .B(n_555), .C(n_590), .D(n_606), .Y(n_460) );
AOI222xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_496), .B1(n_530), .B2(n_543), .C1(n_548), .C2(n_554), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI31xp33_ASAP7_75t_L g722 ( .A1(n_463), .A2(n_723), .A3(n_724), .B(n_726), .Y(n_722) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_475), .Y(n_463) );
AND2x2_ASAP7_75t_L g697 ( .A(n_464), .B(n_477), .Y(n_697) );
BUFx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_SL g547 ( .A(n_465), .Y(n_547) );
AND2x2_ASAP7_75t_L g554 ( .A(n_465), .B(n_487), .Y(n_554) );
AND2x2_ASAP7_75t_L g611 ( .A(n_465), .B(n_478), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_475), .B(n_641), .Y(n_640) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_476), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_476), .B(n_558), .Y(n_601) );
AND2x2_ASAP7_75t_L g694 ( .A(n_476), .B(n_634), .Y(n_694) );
OAI321xp33_ASAP7_75t_L g728 ( .A1(n_476), .A2(n_547), .A3(n_701), .B1(n_729), .B2(n_731), .C(n_732), .Y(n_728) );
NAND4xp25_ASAP7_75t_L g732 ( .A(n_476), .B(n_533), .C(n_641), .D(n_733), .Y(n_732) );
AND2x4_ASAP7_75t_L g476 ( .A(n_477), .B(n_487), .Y(n_476) );
AND2x2_ASAP7_75t_L g596 ( .A(n_477), .B(n_545), .Y(n_596) );
AND2x2_ASAP7_75t_L g615 ( .A(n_477), .B(n_547), .Y(n_615) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g546 ( .A(n_478), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g571 ( .A(n_478), .B(n_487), .Y(n_571) );
AND2x2_ASAP7_75t_L g657 ( .A(n_478), .B(n_545), .Y(n_657) );
INVx3_ASAP7_75t_SL g545 ( .A(n_487), .Y(n_545) );
AND2x2_ASAP7_75t_L g589 ( .A(n_487), .B(n_576), .Y(n_589) );
OR2x2_ASAP7_75t_L g622 ( .A(n_487), .B(n_547), .Y(n_622) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_487), .Y(n_629) );
AND2x2_ASAP7_75t_L g658 ( .A(n_487), .B(n_546), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_487), .B(n_631), .Y(n_673) );
AND2x2_ASAP7_75t_L g705 ( .A(n_487), .B(n_697), .Y(n_705) );
AND2x2_ASAP7_75t_L g714 ( .A(n_487), .B(n_559), .Y(n_714) );
OR2x6_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .Y(n_487) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_509), .Y(n_497) );
INVx1_ASAP7_75t_SL g682 ( .A(n_498), .Y(n_682) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g550 ( .A(n_499), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g532 ( .A(n_500), .B(n_511), .Y(n_532) );
AND2x2_ASAP7_75t_L g618 ( .A(n_500), .B(n_534), .Y(n_618) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g588 ( .A(n_501), .B(n_521), .Y(n_588) );
OR2x2_ASAP7_75t_L g599 ( .A(n_501), .B(n_534), .Y(n_599) );
AND2x2_ASAP7_75t_L g625 ( .A(n_501), .B(n_534), .Y(n_625) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_501), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_509), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_509), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g598 ( .A(n_510), .B(n_599), .Y(n_598) );
AOI322xp5_ASAP7_75t_L g684 ( .A1(n_510), .A2(n_588), .A3(n_594), .B1(n_625), .B2(n_675), .C1(n_685), .C2(n_687), .Y(n_684) );
OR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_521), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_511), .B(n_533), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_511), .B(n_534), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_511), .B(n_551), .Y(n_605) );
AND2x2_ASAP7_75t_L g659 ( .A(n_511), .B(n_625), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_511), .Y(n_663) );
AND2x2_ASAP7_75t_L g675 ( .A(n_511), .B(n_521), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_511), .B(n_550), .Y(n_707) );
INVx4_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g572 ( .A(n_512), .B(n_521), .Y(n_572) );
BUFx3_ASAP7_75t_L g586 ( .A(n_512), .Y(n_586) );
AND3x2_ASAP7_75t_L g668 ( .A(n_512), .B(n_648), .C(n_669), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_521), .B(n_532), .C(n_533), .Y(n_531) );
INVx1_ASAP7_75t_SL g551 ( .A(n_521), .Y(n_551) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_521), .Y(n_653) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g647 ( .A(n_532), .B(n_648), .Y(n_647) );
INVxp67_ASAP7_75t_L g654 ( .A(n_532), .Y(n_654) );
AND2x2_ASAP7_75t_L g692 ( .A(n_533), .B(n_670), .Y(n_692) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx3_ASAP7_75t_L g573 ( .A(n_534), .Y(n_573) );
AND2x2_ASAP7_75t_L g648 ( .A(n_534), .B(n_551), .Y(n_648) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
OR2x2_ASAP7_75t_L g592 ( .A(n_545), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g711 ( .A(n_545), .B(n_611), .Y(n_711) );
AND2x2_ASAP7_75t_L g725 ( .A(n_545), .B(n_547), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_546), .B(n_559), .Y(n_666) );
AND2x2_ASAP7_75t_L g713 ( .A(n_546), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g576 ( .A(n_547), .B(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g593 ( .A(n_547), .B(n_559), .Y(n_593) );
INVx1_ASAP7_75t_L g603 ( .A(n_547), .Y(n_603) );
AND2x2_ASAP7_75t_L g634 ( .A(n_547), .B(n_559), .Y(n_634) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_549), .A2(n_677), .B1(n_681), .B2(n_683), .C(n_684), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_550), .B(n_552), .Y(n_549) );
AND2x2_ASAP7_75t_L g580 ( .A(n_550), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_553), .B(n_587), .Y(n_730) );
AOI322xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_572), .A3(n_573), .B1(n_574), .B2(n_580), .C1(n_582), .C2(n_589), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_571), .Y(n_557) );
NAND2x1p5_ASAP7_75t_L g610 ( .A(n_558), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_558), .B(n_621), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_558), .A2(n_571), .B(n_645), .C(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_558), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_558), .B(n_615), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_558), .B(n_697), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_558), .B(n_725), .Y(n_724) );
BUFx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_559), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_559), .B(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g686 ( .A(n_559), .B(n_573), .Y(n_686) );
OA21x2_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_563), .B(n_570), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_561), .A2(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g578 ( .A(n_563), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_570), .Y(n_579) );
INVx1_ASAP7_75t_L g661 ( .A(n_571), .Y(n_661) );
OAI31xp33_ASAP7_75t_L g671 ( .A1(n_571), .A2(n_596), .A3(n_672), .B(n_674), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_571), .B(n_577), .Y(n_723) );
INVx1_ASAP7_75t_SL g584 ( .A(n_572), .Y(n_584) );
AND2x2_ASAP7_75t_L g617 ( .A(n_572), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g698 ( .A(n_572), .B(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g583 ( .A(n_573), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g608 ( .A(n_573), .Y(n_608) );
AND2x2_ASAP7_75t_L g635 ( .A(n_573), .B(n_588), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_573), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g727 ( .A(n_573), .B(n_675), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_575), .B(n_645), .Y(n_718) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g614 ( .A(n_577), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g632 ( .A(n_577), .Y(n_632) );
NAND2xp33_ASAP7_75t_SL g582 ( .A(n_583), .B(n_585), .Y(n_582) );
OAI211xp5_ASAP7_75t_SL g626 ( .A1(n_584), .A2(n_627), .B(n_633), .C(n_649), .Y(n_626) );
OR2x2_ASAP7_75t_L g701 ( .A(n_584), .B(n_682), .Y(n_701) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
CKINVDCx16_ASAP7_75t_R g638 ( .A(n_586), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_586), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g607 ( .A(n_588), .B(n_608), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_594), .B(n_597), .C(n_600), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_SL g641 ( .A(n_593), .Y(n_641) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_596), .B(n_634), .Y(n_639) );
INVx1_ASAP7_75t_L g645 ( .A(n_596), .Y(n_645) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g604 ( .A(n_599), .B(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g637 ( .A(n_599), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g699 ( .A(n_599), .Y(n_699) );
AOI21xp33_ASAP7_75t_SL g600 ( .A1(n_601), .A2(n_602), .B(n_604), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_602), .A2(n_613), .B(n_616), .Y(n_612) );
AOI211xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_609), .B(n_612), .C(n_619), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_607), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_610), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g623 ( .A(n_611), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_613), .A2(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_618), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g643 ( .A(n_618), .Y(n_643) );
AOI21xp33_ASAP7_75t_SL g619 ( .A1(n_620), .A2(n_623), .B(n_624), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g674 ( .A(n_625), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_631), .B(n_657), .Y(n_683) );
AND2x2_ASAP7_75t_L g696 ( .A(n_631), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g710 ( .A(n_631), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g720 ( .A(n_631), .B(n_658), .Y(n_720) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI211xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B(n_636), .C(n_644), .Y(n_633) );
INVx1_ASAP7_75t_L g680 ( .A(n_634), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B1(n_640), .B2(n_642), .Y(n_636) );
OR2x2_ASAP7_75t_L g642 ( .A(n_638), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_638), .B(n_699), .Y(n_721) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g715 ( .A(n_648), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_655), .B1(n_658), .B2(n_659), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g733 ( .A(n_653), .Y(n_733) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g679 ( .A(n_657), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_662), .B(n_664), .C(n_671), .Y(n_660) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVx2_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_679), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR5xp2_ASAP7_75t_L g689 ( .A(n_690), .B(n_708), .C(n_716), .D(n_722), .E(n_728), .Y(n_689) );
OAI211xp5_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_693), .B(n_695), .C(n_702), .Y(n_690) );
INVxp67_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B(n_700), .Y(n_695) );
OAI21xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .B(n_706), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_705), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_712), .B(n_715), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g731 ( .A(n_711), .Y(n_731) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_719), .B(n_721), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
CKINVDCx16_ASAP7_75t_R g743 ( .A(n_734), .Y(n_743) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx3_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
endmodule