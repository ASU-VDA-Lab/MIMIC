module real_aes_1249_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_503;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_564;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_0), .A2(n_67), .B1(n_120), .B2(n_123), .Y(n_119) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_1), .A2(n_55), .B1(n_90), .B2(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g170 ( .A(n_2), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g153 ( .A1(n_3), .A2(n_13), .B1(n_154), .B2(n_155), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_3), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_4), .B(n_197), .Y(n_220) );
INVx1_ASAP7_75t_L g242 ( .A(n_5), .Y(n_242) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_6), .A2(n_19), .B1(n_90), .B2(n_98), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_7), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_8), .A2(n_39), .B1(n_133), .B2(n_137), .Y(n_132) );
INVx2_ASAP7_75t_L g196 ( .A(n_9), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g140 ( .A1(n_10), .A2(n_24), .B1(n_141), .B2(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g230 ( .A(n_11), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_12), .A2(n_76), .B1(n_146), .B2(n_147), .Y(n_145) );
INVx1_ASAP7_75t_L g155 ( .A(n_13), .Y(n_155) );
INVx1_ASAP7_75t_L g227 ( .A(n_14), .Y(n_227) );
INVx1_ASAP7_75t_SL g302 ( .A(n_15), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_16), .B(n_207), .Y(n_206) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_17), .Y(n_151) );
AOI33xp33_ASAP7_75t_L g279 ( .A1(n_17), .A2(n_36), .A3(n_187), .B1(n_202), .B2(n_280), .B3(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g251 ( .A(n_18), .Y(n_251) );
OAI221xp5_ASAP7_75t_L g162 ( .A1(n_19), .A2(n_55), .B1(n_57), .B2(n_163), .C(n_165), .Y(n_162) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_20), .A2(n_69), .B(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_L g198 ( .A(n_20), .B(n_69), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_21), .B(n_240), .Y(n_299) );
INVx3_ASAP7_75t_L g90 ( .A(n_22), .Y(n_90) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_23), .A2(n_150), .B1(n_157), .B2(n_158), .Y(n_149) );
INVx1_ASAP7_75t_L g157 ( .A(n_23), .Y(n_157) );
INVx1_ASAP7_75t_SL g91 ( .A(n_25), .Y(n_91) );
INVx1_ASAP7_75t_L g172 ( .A(n_26), .Y(n_172) );
AND2x2_ASAP7_75t_L g191 ( .A(n_26), .B(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g216 ( .A(n_26), .B(n_170), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_27), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_28), .B(n_240), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_29), .A2(n_184), .B1(n_194), .B2(n_197), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_30), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_31), .B(n_207), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_32), .B(n_218), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_33), .B(n_207), .Y(n_243) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_34), .A2(n_57), .B1(n_90), .B2(n_94), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_35), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_37), .B(n_207), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_38), .A2(n_64), .B1(n_104), .B2(n_108), .Y(n_103) );
INVx1_ASAP7_75t_L g188 ( .A(n_40), .Y(n_188) );
INVx1_ASAP7_75t_L g209 ( .A(n_40), .Y(n_209) );
AND2x2_ASAP7_75t_L g271 ( .A(n_41), .B(n_272), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g239 ( .A1(n_42), .A2(n_60), .B1(n_200), .B2(n_240), .C(n_241), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_43), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_44), .B(n_240), .Y(n_294) );
INVx1_ASAP7_75t_L g92 ( .A(n_45), .Y(n_92) );
AOI22xp33_ASAP7_75t_SL g127 ( .A1(n_46), .A2(n_59), .B1(n_128), .B2(n_130), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_47), .B(n_194), .Y(n_260) );
AOI21xp5_ASAP7_75t_SL g290 ( .A1(n_48), .A2(n_200), .B(n_291), .Y(n_290) );
AOI22xp33_ASAP7_75t_SL g112 ( .A1(n_49), .A2(n_72), .B1(n_113), .B2(n_116), .Y(n_112) );
INVx1_ASAP7_75t_L g223 ( .A(n_50), .Y(n_223) );
OAI22xp5_ASAP7_75t_SL g556 ( .A1(n_51), .A2(n_80), .B1(n_81), .B2(n_557), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_51), .Y(n_557) );
INVx1_ASAP7_75t_L g269 ( .A(n_52), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_53), .A2(n_80), .B1(n_81), .B2(n_148), .Y(n_79) );
INVx1_ASAP7_75t_L g148 ( .A(n_53), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_54), .A2(n_200), .B(n_268), .Y(n_267) );
INVxp33_ASAP7_75t_L g167 ( .A(n_55), .Y(n_167) );
INVx1_ASAP7_75t_L g192 ( .A(n_56), .Y(n_192) );
INVx1_ASAP7_75t_L g211 ( .A(n_56), .Y(n_211) );
INVxp67_ASAP7_75t_L g166 ( .A(n_57), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_58), .B(n_240), .Y(n_282) );
AND2x2_ASAP7_75t_L g304 ( .A(n_61), .B(n_247), .Y(n_304) );
INVx1_ASAP7_75t_L g224 ( .A(n_62), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_63), .A2(n_200), .B(n_301), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_65), .A2(n_200), .B(n_205), .C(n_217), .Y(n_199) );
AND2x2_ASAP7_75t_SL g288 ( .A(n_66), .B(n_247), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_68), .A2(n_200), .B1(n_277), .B2(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g292 ( .A(n_70), .Y(n_292) );
AND2x2_ASAP7_75t_L g283 ( .A(n_71), .B(n_247), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_73), .A2(n_249), .B(n_250), .C(n_252), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_73), .A2(n_80), .B1(n_81), .B2(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_73), .Y(n_548) );
BUFx2_ASAP7_75t_SL g164 ( .A(n_74), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_75), .B(n_207), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_159), .B1(n_173), .B2(n_544), .C(n_546), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_149), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND2x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_125), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_111), .Y(n_83) );
OAI21xp5_ASAP7_75t_SL g84 ( .A1(n_85), .A2(n_102), .B(n_103), .Y(n_84) );
INVx2_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
AND2x4_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
AND2x2_ASAP7_75t_L g116 ( .A(n_87), .B(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g123 ( .A(n_87), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
AND2x2_ASAP7_75t_L g106 ( .A(n_88), .B(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_88), .Y(n_109) );
INVx2_ASAP7_75t_L g122 ( .A(n_88), .Y(n_122) );
OAI22x1_ASAP7_75t_L g88 ( .A1(n_89), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g94 ( .A(n_90), .Y(n_94) );
INVx2_ASAP7_75t_L g98 ( .A(n_90), .Y(n_98) );
INVx1_ASAP7_75t_L g101 ( .A(n_90), .Y(n_101) );
INVx2_ASAP7_75t_L g107 ( .A(n_93), .Y(n_107) );
AND2x2_ASAP7_75t_L g121 ( .A(n_93), .B(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g131 ( .A(n_93), .Y(n_131) );
AND2x4_ASAP7_75t_L g135 ( .A(n_95), .B(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g142 ( .A(n_95), .B(n_106), .Y(n_142) );
AND2x6_ASAP7_75t_L g146 ( .A(n_95), .B(n_121), .Y(n_146) );
AND2x4_ASAP7_75t_L g95 ( .A(n_96), .B(n_99), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x4_ASAP7_75t_L g105 ( .A(n_97), .B(n_99), .Y(n_105) );
AND2x2_ASAP7_75t_L g110 ( .A(n_97), .B(n_100), .Y(n_110) );
INVx1_ASAP7_75t_L g115 ( .A(n_97), .Y(n_115) );
INVxp67_ASAP7_75t_L g124 ( .A(n_99), .Y(n_124) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g114 ( .A(n_100), .B(n_115), .Y(n_114) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g120 ( .A(n_105), .B(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g138 ( .A(n_105), .B(n_136), .Y(n_138) );
AND2x4_ASAP7_75t_L g113 ( .A(n_106), .B(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g136 ( .A(n_107), .B(n_122), .Y(n_136) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x4_ASAP7_75t_L g130 ( .A(n_110), .B(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g144 ( .A(n_110), .B(n_136), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_119), .Y(n_111) );
AND2x2_ASAP7_75t_L g129 ( .A(n_114), .B(n_121), .Y(n_129) );
AND2x6_ASAP7_75t_L g147 ( .A(n_114), .B(n_136), .Y(n_147) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_115), .Y(n_118) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NOR2x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_139), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_132), .Y(n_126) );
BUFx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx3_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
INVx8_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_145), .Y(n_139) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_150), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B1(n_153), .B2(n_156), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_151), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_161), .Y(n_160) );
AND3x1_ASAP7_75t_SL g161 ( .A(n_162), .B(n_168), .C(n_171), .Y(n_161) );
INVxp67_ASAP7_75t_L g554 ( .A(n_162), .Y(n_554) );
CKINVDCx8_ASAP7_75t_R g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
CKINVDCx16_ASAP7_75t_R g552 ( .A(n_168), .Y(n_552) );
AO21x1_ASAP7_75t_SL g563 ( .A1(n_168), .A2(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g186 ( .A(n_169), .B(n_187), .Y(n_186) );
OR2x2_ASAP7_75t_SL g560 ( .A(n_169), .B(n_171), .Y(n_560) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g204 ( .A(n_170), .B(n_188), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_171), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2x1p5_ASAP7_75t_L g201 ( .A(n_172), .B(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_478), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_401), .Y(n_176) );
NAND3xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_348), .C(n_381), .Y(n_177) );
AOI211xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_305), .B(n_314), .C(n_338), .Y(n_178) );
OAI21xp33_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_234), .B(n_284), .Y(n_179) );
OR2x2_ASAP7_75t_L g358 ( .A(n_180), .B(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g513 ( .A(n_180), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_181), .A2(n_404), .B1(n_408), .B2(n_410), .Y(n_403) );
AND2x2_ASAP7_75t_L g440 ( .A(n_181), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_219), .Y(n_181) );
INVx1_ASAP7_75t_L g337 ( .A(n_182), .Y(n_337) );
AND2x4_ASAP7_75t_L g354 ( .A(n_182), .B(n_335), .Y(n_354) );
INVx2_ASAP7_75t_L g376 ( .A(n_182), .Y(n_376) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_182), .Y(n_459) );
AND2x2_ASAP7_75t_L g530 ( .A(n_182), .B(n_287), .Y(n_530) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_199), .Y(n_182) );
NOR3xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_189), .C(n_193), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x4_ASAP7_75t_L g240 ( .A(n_186), .B(n_190), .Y(n_240) );
OR2x6_ASAP7_75t_L g214 ( .A(n_187), .B(n_203), .Y(n_214) );
INVxp33_ASAP7_75t_L g280 ( .A(n_187), .Y(n_280) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_187), .Y(n_565) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x4_ASAP7_75t_L g232 ( .A(n_188), .B(n_210), .Y(n_232) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g203 ( .A(n_192), .Y(n_203) );
AND2x6_ASAP7_75t_L g229 ( .A(n_192), .B(n_208), .Y(n_229) );
INVx4_ASAP7_75t_L g247 ( .A(n_194), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_194), .B(n_257), .Y(n_256) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
BUFx4f_ASAP7_75t_L g218 ( .A(n_195), .Y(n_218) );
AND2x4_ASAP7_75t_L g197 ( .A(n_196), .B(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_SL g273 ( .A(n_196), .B(n_198), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_197), .B(n_215), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_197), .A2(n_290), .B(n_294), .Y(n_289) );
INVxp67_ASAP7_75t_L g259 ( .A(n_200), .Y(n_259) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_204), .Y(n_200) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_201), .Y(n_564) );
INVx1_ASAP7_75t_L g281 ( .A(n_202), .Y(n_281) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_212), .B(n_215), .Y(n_205) );
INVx1_ASAP7_75t_L g225 ( .A(n_207), .Y(n_225) );
AND2x4_ASAP7_75t_L g545 ( .A(n_207), .B(n_216), .Y(n_545) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_210), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_214), .A2(n_223), .B1(n_224), .B2(n_225), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_SL g241 ( .A1(n_214), .A2(n_215), .B(n_242), .C(n_243), .Y(n_241) );
INVxp67_ASAP7_75t_L g249 ( .A(n_214), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_214), .A2(n_215), .B(n_269), .C(n_270), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g291 ( .A1(n_214), .A2(n_215), .B(n_292), .C(n_293), .Y(n_291) );
O2A1O1Ixp33_ASAP7_75t_SL g301 ( .A1(n_214), .A2(n_215), .B(n_302), .C(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g277 ( .A(n_215), .Y(n_277) );
INVx5_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_216), .Y(n_252) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_217), .A2(n_275), .B(n_283), .Y(n_274) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_217), .A2(n_275), .B(n_283), .Y(n_319) );
INVx2_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_218), .A2(n_239), .B(n_244), .Y(n_238) );
AND2x2_ASAP7_75t_L g295 ( .A(n_219), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g324 ( .A(n_219), .Y(n_324) );
INVx3_ASAP7_75t_L g335 ( .A(n_219), .Y(n_335) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_226), .B(n_233), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_225), .B(n_251), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B1(n_230), .B2(n_231), .Y(n_226) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVxp67_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_234), .A2(n_525), .B1(n_527), .B2(n_529), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_234), .B(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_262), .Y(n_235) );
INVx3_ASAP7_75t_L g308 ( .A(n_236), .Y(n_308) );
AND2x2_ASAP7_75t_L g316 ( .A(n_236), .B(n_317), .Y(n_316) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_236), .Y(n_346) );
NAND2x1_ASAP7_75t_SL g540 ( .A(n_236), .B(n_307), .Y(n_540) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_245), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g313 ( .A(n_238), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_238), .B(n_319), .Y(n_331) );
AND2x2_ASAP7_75t_L g344 ( .A(n_238), .B(n_245), .Y(n_344) );
AND2x4_ASAP7_75t_L g351 ( .A(n_238), .B(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_238), .Y(n_400) );
INVxp67_ASAP7_75t_L g407 ( .A(n_238), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_238), .Y(n_412) );
INVx1_ASAP7_75t_L g261 ( .A(n_240), .Y(n_261) );
INVx1_ASAP7_75t_L g311 ( .A(n_245), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_245), .B(n_321), .Y(n_330) );
INVx2_ASAP7_75t_L g398 ( .A(n_245), .Y(n_398) );
INVx1_ASAP7_75t_L g437 ( .A(n_245), .Y(n_437) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_255), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B1(n_253), .B2(n_254), .Y(n_246) );
INVx3_ASAP7_75t_L g254 ( .A(n_247), .Y(n_254) );
OAI222xp33_ASAP7_75t_L g546 ( .A1(n_251), .A2(n_547), .B1(n_549), .B2(n_555), .C1(n_558), .C2(n_561), .Y(n_546) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_254), .A2(n_265), .B(n_271), .Y(n_264) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_254), .A2(n_265), .B(n_271), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_259), .B1(n_260), .B2(n_261), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g367 ( .A(n_262), .B(n_344), .Y(n_367) );
AND2x2_ASAP7_75t_L g435 ( .A(n_262), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g449 ( .A(n_262), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_262), .B(n_464), .Y(n_463) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_274), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NOR2x1_ASAP7_75t_L g312 ( .A(n_264), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g405 ( .A(n_264), .B(n_398), .Y(n_405) );
AND2x2_ASAP7_75t_L g496 ( .A(n_264), .B(n_318), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_272), .Y(n_297) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g307 ( .A(n_274), .Y(n_307) );
INVx2_ASAP7_75t_L g352 ( .A(n_274), .Y(n_352) );
AND2x2_ASAP7_75t_L g397 ( .A(n_274), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_276), .B(n_282), .Y(n_275) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_295), .Y(n_285) );
AND2x2_ASAP7_75t_L g439 ( .A(n_286), .B(n_440), .Y(n_439) );
OR2x6_ASAP7_75t_L g498 ( .A(n_286), .B(n_499), .Y(n_498) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx4_ASAP7_75t_L g328 ( .A(n_287), .Y(n_328) );
AND2x4_ASAP7_75t_L g336 ( .A(n_287), .B(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g371 ( .A(n_287), .B(n_296), .Y(n_371) );
INVx2_ASAP7_75t_L g420 ( .A(n_287), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_287), .B(n_394), .Y(n_469) );
AND2x2_ASAP7_75t_L g506 ( .A(n_287), .B(n_324), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_287), .B(n_389), .Y(n_514) );
OR2x6_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AND2x2_ASAP7_75t_L g347 ( .A(n_295), .B(n_336), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_295), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_SL g486 ( .A(n_295), .B(n_374), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_295), .B(n_387), .Y(n_508) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
AND2x2_ASAP7_75t_L g334 ( .A(n_296), .B(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_296), .Y(n_357) );
INVx2_ASAP7_75t_L g360 ( .A(n_296), .Y(n_360) );
INVx1_ASAP7_75t_L g393 ( .A(n_296), .Y(n_393) );
INVx1_ASAP7_75t_L g441 ( .A(n_296), .Y(n_441) );
AO21x2_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B(n_304), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NAND2xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_307), .B(n_310), .Y(n_383) );
OR2x2_ASAP7_75t_L g455 ( .A(n_307), .B(n_456), .Y(n_455) );
AND4x1_ASAP7_75t_SL g501 ( .A(n_307), .B(n_483), .C(n_502), .D(n_503), .Y(n_501) );
OR2x2_ASAP7_75t_L g525 ( .A(n_308), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g362 ( .A(n_311), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_311), .B(n_320), .Y(n_512) );
AND2x2_ASAP7_75t_L g537 ( .A(n_312), .B(n_397), .Y(n_537) );
OAI32xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_322), .A3(n_327), .B1(n_329), .B2(n_332), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g410 ( .A(n_317), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g510 ( .A(n_317), .B(n_464), .Y(n_510) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
AND2x2_ASAP7_75t_L g406 ( .A(n_318), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g492 ( .A(n_318), .Y(n_492) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_319), .B(n_321), .Y(n_526) );
INVx3_ASAP7_75t_L g343 ( .A(n_320), .Y(n_343) );
NAND2x1p5_ASAP7_75t_L g521 ( .A(n_320), .B(n_448), .Y(n_521) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_321), .Y(n_380) );
AND2x2_ASAP7_75t_L g399 ( .A(n_321), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g533 ( .A(n_323), .Y(n_533) );
NAND2x1_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g373 ( .A(n_324), .Y(n_373) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_324), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_327), .B(n_433), .Y(n_432) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g365 ( .A(n_328), .B(n_333), .Y(n_365) );
AND2x4_ASAP7_75t_L g387 ( .A(n_328), .B(n_337), .Y(n_387) );
AND2x4_ASAP7_75t_SL g458 ( .A(n_328), .B(n_459), .Y(n_458) );
NOR2x1_ASAP7_75t_L g484 ( .A(n_328), .B(n_409), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_329), .A2(n_452), .B1(n_455), .B2(n_457), .Y(n_451) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx2_ASAP7_75t_SL g471 ( .A(n_330), .Y(n_471) );
INVx2_ASAP7_75t_L g363 ( .A(n_331), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_336), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_334), .B(n_340), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_334), .A2(n_470), .B1(n_473), .B2(n_476), .Y(n_472) );
INVx1_ASAP7_75t_L g394 ( .A(n_335), .Y(n_394) );
AND2x2_ASAP7_75t_L g417 ( .A(n_335), .B(n_376), .Y(n_417) );
INVx2_ASAP7_75t_L g340 ( .A(n_336), .Y(n_340) );
OAI21xp5_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_341), .B(n_345), .Y(n_338) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_342), .A2(n_414), .B1(n_418), .B2(n_419), .Y(n_413) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_343), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_343), .B(n_411), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_343), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
NOR3xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_364), .C(n_368), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_353), .B1(n_358), .B2(n_361), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g378 ( .A(n_351), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g418 ( .A(n_351), .B(n_405), .Y(n_418) );
AND2x2_ASAP7_75t_L g470 ( .A(n_351), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g487 ( .A(n_351), .B(n_437), .Y(n_487) );
AND2x2_ASAP7_75t_L g542 ( .A(n_351), .B(n_436), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx4_ASAP7_75t_L g409 ( .A(n_354), .Y(n_409) );
AND2x2_ASAP7_75t_L g419 ( .A(n_354), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g424 ( .A(n_357), .Y(n_424) );
AND2x2_ASAP7_75t_L g433 ( .A(n_357), .B(n_417), .Y(n_433) );
INVx1_ASAP7_75t_L g468 ( .A(n_359), .Y(n_468) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g389 ( .A(n_360), .Y(n_389) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_362), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_363), .B(n_431), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B(n_377), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_370), .B(n_409), .Y(n_518) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
AOI21xp33_ASAP7_75t_SL g381 ( .A1(n_373), .A2(n_382), .B(n_384), .Y(n_381) );
AND2x2_ASAP7_75t_L g528 ( .A(n_373), .B(n_387), .Y(n_528) );
AND2x4_ASAP7_75t_L g391 ( .A(n_374), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_SL g425 ( .A(n_374), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_374), .B(n_441), .Y(n_507) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI21xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_390), .B(n_395), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_387), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_387), .B(n_392), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_388), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g450 ( .A(n_388), .Y(n_450) );
INVx1_ASAP7_75t_L g454 ( .A(n_388), .Y(n_454) );
AND2x2_ASAP7_75t_L g538 ( .A(n_388), .B(n_506), .Y(n_538) );
AND2x2_ASAP7_75t_L g541 ( .A(n_388), .B(n_458), .Y(n_541) );
INVx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_SL g392 ( .A(n_393), .B(n_394), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_393), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
INVx1_ASAP7_75t_L g520 ( .A(n_397), .Y(n_520) );
AND2x2_ASAP7_75t_L g411 ( .A(n_398), .B(n_412), .Y(n_411) );
NAND4xp75_ASAP7_75t_L g401 ( .A(n_402), .B(n_421), .C(n_442), .D(n_460), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_413), .Y(n_402) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
NAND2x1p5_ASAP7_75t_L g491 ( .A(n_405), .B(n_492), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g477 ( .A(n_406), .B(n_471), .Y(n_477) );
NAND2xp5_ASAP7_75t_R g493 ( .A(n_409), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g543 ( .A(n_409), .Y(n_543) );
INVx2_ASAP7_75t_L g456 ( .A(n_411), .Y(n_456) );
BUFx3_ASAP7_75t_L g448 ( .A(n_412), .Y(n_448) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g499 ( .A(n_417), .Y(n_499) );
AND2x2_ASAP7_75t_L g453 ( .A(n_419), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g475 ( .A(n_420), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_426), .B(n_428), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_424), .B(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_425), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_427), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_432), .B1(n_434), .B2(n_438), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_436), .A2(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g464 ( .A(n_436), .Y(n_464) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g495 ( .A(n_437), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g503 ( .A(n_437), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_438), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g473 ( .A(n_441), .B(n_474), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_449), .B(n_451), .Y(n_442) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g490 ( .A(n_447), .B(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_454), .Y(n_502) );
INVx2_ASAP7_75t_SL g494 ( .A(n_458), .Y(n_494) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_472), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_465), .B1(n_467), .B2(n_470), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g523 ( .A(n_467), .Y(n_523) );
NOR2x1_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_515), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_488), .C(n_500), .Y(n_479) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_481), .B(n_485), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g488 ( .A1(n_489), .A2(n_493), .B1(n_495), .B2(n_497), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_504), .C(n_511), .Y(n_500) );
AOI21xp33_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_508), .B(n_509), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_534), .Y(n_515) );
NOR3xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_524), .C(n_531), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_522), .B2(n_523), .Y(n_517) );
OR2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g531 ( .A(n_525), .B(n_530), .C(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVxp67_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AOI222xp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_538), .B1(n_539), .B2(n_541), .C1(n_542), .C2(n_543), .Y(n_534) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_550), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVxp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_562), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_563), .Y(n_562) );
endmodule