module fake_jpeg_2263_n_160 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_53),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_43),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_49),
.B1(n_64),
.B2(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_46),
.C(n_55),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_87),
.Y(n_99)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_52),
.C(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_51),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_0),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_22),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_1),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_1),
.CI(n_2),
.CON(n_93),
.SN(n_93)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_96),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_76),
.Y(n_96)
);

NOR2x1_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_109),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_45),
.B(n_56),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_6),
.B(n_7),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_2),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_108),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_69),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_34),
.C(n_33),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_108),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_113),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_80),
.B1(n_45),
.B2(n_5),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_112),
.B1(n_117),
.B2(n_127),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_16),
.B1(n_37),
.B2(n_35),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_15),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_121),
.C(n_122),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_39),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_3),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_128),
.A2(n_8),
.B(n_9),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_104),
.Y(n_129)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_135),
.A3(n_123),
.B1(n_120),
.B2(n_122),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_12),
.B(n_28),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_8),
.C(n_9),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_112),
.B1(n_117),
.B2(n_13),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_144),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_27),
.B(n_30),
.C(n_29),
.D(n_23),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_146),
.A2(n_147),
.B1(n_131),
.B2(n_133),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_129),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_143),
.B1(n_141),
.B2(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_151),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_152),
.B1(n_148),
.B2(n_149),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_145),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_141),
.B(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_135),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_157),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_140),
.B(n_32),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_140),
.Y(n_160)
);


endmodule