module fake_jpeg_1466_n_529 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_529);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_529;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_SL g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_57),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_26),
.A2(n_10),
.B(n_16),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_61),
.B(n_0),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_10),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_64),
.B(n_74),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_67),
.Y(n_202)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_69),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_9),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_73),
.B(n_101),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_11),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_76),
.B(n_77),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_18),
.B(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_34),
.B(n_8),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_78),
.B(n_84),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_81),
.Y(n_167)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_35),
.B(n_8),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_85),
.Y(n_147)
);

BUFx16f_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_88),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_90),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_91),
.Y(n_204)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_21),
.B(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_116),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_100),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_21),
.B(n_8),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

BUFx8_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_120),
.Y(n_137)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_39),
.Y(n_109)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_111),
.Y(n_193)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_46),
.B(n_7),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_22),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_118),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_22),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_22),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_25),
.Y(n_170)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_121),
.B(n_122),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_26),
.B1(n_42),
.B2(n_27),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_128),
.A2(n_143),
.B1(n_149),
.B2(n_161),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_73),
.A2(n_25),
.B1(n_27),
.B2(n_54),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_129),
.A2(n_199),
.B1(n_90),
.B2(n_91),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_55),
.C(n_46),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_133),
.B(n_155),
.C(n_174),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_26),
.B1(n_42),
.B2(n_55),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_107),
.A2(n_43),
.B1(n_54),
.B2(n_24),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_24),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_152),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_53),
.B1(n_41),
.B2(n_45),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_163),
.B(n_168),
.Y(n_228)
);

AO22x1_ASAP7_75t_SL g168 ( 
.A1(n_121),
.A2(n_54),
.B1(n_36),
.B2(n_45),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_72),
.A2(n_54),
.B1(n_53),
.B2(n_41),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_169),
.A2(n_175),
.B1(n_180),
.B2(n_181),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_200),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_85),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_171),
.B(n_189),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_122),
.A2(n_45),
.B1(n_36),
.B2(n_25),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_60),
.A2(n_32),
.B1(n_30),
.B2(n_45),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_112),
.A2(n_45),
.B1(n_36),
.B2(n_32),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_70),
.A2(n_36),
.B1(n_30),
.B2(n_2),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_194),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_100),
.A2(n_36),
.B1(n_13),
.B2(n_2),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_184),
.A2(n_197),
.B1(n_201),
.B2(n_16),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_58),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_185),
.A2(n_192),
.B1(n_201),
.B2(n_197),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_61),
.B(n_7),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_62),
.A2(n_69),
.B1(n_105),
.B2(n_103),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_81),
.B(n_13),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_99),
.B(n_14),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_195),
.B(n_147),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_108),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_65),
.A2(n_0),
.B1(n_1),
.B2(n_14),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_87),
.B(n_15),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_109),
.A2(n_15),
.B1(n_16),
.B2(n_0),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_110),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_205),
.B(n_212),
.Y(n_273)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_206),
.Y(n_279)
);

OR2x2_ASAP7_75t_SL g208 ( 
.A(n_130),
.B(n_102),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_208),
.B(n_220),
.Y(n_297)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_209),
.Y(n_306)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_210),
.Y(n_274)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_211),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_1),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_214),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_159),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_215),
.B(n_237),
.Y(n_304)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_147),
.Y(n_216)
);

INVx4_ASAP7_75t_SL g276 ( 
.A(n_216),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_124),
.B(n_89),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_217),
.B(n_219),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_83),
.B1(n_94),
.B2(n_67),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_218),
.A2(n_221),
.B1(n_225),
.B2(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_79),
.Y(n_219)
);

OR2x2_ASAP7_75t_SL g220 ( 
.A(n_148),
.B(n_15),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_222),
.Y(n_289)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_134),
.Y(n_223)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_223),
.Y(n_292)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_145),
.Y(n_224)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_224),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_168),
.A2(n_161),
.B1(n_200),
.B2(n_156),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_226),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_150),
.B(n_95),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_227),
.B(n_232),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_152),
.A2(n_169),
.B(n_137),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_229),
.A2(n_245),
.B(n_264),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_127),
.Y(n_230)
);

INVx3_ASAP7_75t_SL g318 ( 
.A(n_230),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_151),
.B(n_157),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_231),
.B(n_249),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_131),
.B(n_146),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_127),
.Y(n_235)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_175),
.A2(n_143),
.B1(n_180),
.B2(n_185),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_236),
.A2(n_247),
.B1(n_258),
.B2(n_265),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_131),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_160),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_240),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_142),
.Y(n_239)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_239),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_141),
.B(n_158),
.Y(n_240)
);

AO22x1_ASAP7_75t_L g242 ( 
.A1(n_194),
.A2(n_136),
.B1(n_135),
.B2(n_126),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g298 ( 
.A1(n_242),
.A2(n_228),
.B(n_244),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_254),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_138),
.B(n_123),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_246),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_149),
.A2(n_128),
.B(n_184),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_142),
.Y(n_248)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_248),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_139),
.B(n_144),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_191),
.Y(n_250)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_250),
.Y(n_321)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_125),
.Y(n_251)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_251),
.Y(n_323)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_125),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_259),
.Y(n_290)
);

OAI32xp33_ASAP7_75t_L g253 ( 
.A1(n_138),
.A2(n_198),
.A3(n_193),
.B1(n_162),
.B2(n_186),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_242),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_155),
.B(n_173),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_255),
.B(n_256),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_132),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_205),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_132),
.A2(n_140),
.B1(n_179),
.B2(n_204),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_164),
.B(n_140),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_167),
.B(n_173),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_260),
.B(n_266),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_167),
.A2(n_164),
.B1(n_183),
.B2(n_187),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_261),
.A2(n_267),
.B1(n_216),
.B2(n_252),
.Y(n_322)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_183),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_268),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_179),
.A2(n_187),
.B(n_154),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_153),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_153),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_267),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_203),
.B(n_154),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_202),
.B(n_145),
.C(n_134),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_229),
.C(n_228),
.Y(n_295)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_202),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_271),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_203),
.B(n_124),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_199),
.A2(n_181),
.B1(n_129),
.B2(n_195),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g332 ( 
.A(n_277),
.B(n_295),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_280),
.A2(n_287),
.B1(n_307),
.B2(n_317),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_225),
.A2(n_234),
.B1(n_272),
.B2(n_221),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_212),
.B(n_217),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_291),
.B(n_293),
.C(n_273),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_219),
.B(n_231),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_301),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_262),
.A2(n_228),
.B(n_213),
.C(n_241),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_299),
.A2(n_263),
.B(n_239),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_207),
.B(n_269),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_308),
.Y(n_345)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_208),
.B(n_257),
.CI(n_220),
.CON(n_303),
.SN(n_303)
);

XNOR2x1_ASAP7_75t_SL g355 ( 
.A(n_303),
.B(n_299),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_234),
.A2(n_245),
.B1(n_247),
.B2(n_268),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_249),
.B(n_242),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_259),
.A2(n_258),
.B1(n_264),
.B2(n_211),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_251),
.B1(n_210),
.B2(n_209),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_223),
.B(n_224),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_273),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_237),
.A2(n_244),
.B1(n_266),
.B2(n_270),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_322),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_280),
.A2(n_267),
.B1(n_253),
.B2(n_206),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_324),
.A2(n_327),
.B1(n_333),
.B2(n_335),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_275),
.B(n_250),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_330),
.Y(n_363)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_328),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_281),
.B(n_214),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_283),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_336),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_296),
.A2(n_235),
.B1(n_230),
.B2(n_255),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_334),
.A2(n_306),
.B(n_276),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_281),
.A2(n_248),
.B1(n_246),
.B2(n_233),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_283),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_308),
.A2(n_222),
.B1(n_246),
.B2(n_285),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_338),
.A2(n_343),
.B1(n_347),
.B2(n_356),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_294),
.Y(n_339)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_339),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_340),
.B(n_352),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_277),
.B(n_246),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_341),
.B(n_361),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_316),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_344),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_301),
.A2(n_295),
.B1(n_285),
.B2(n_298),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_292),
.B(n_311),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_346),
.B(n_355),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_298),
.A2(n_293),
.B1(n_315),
.B2(n_300),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_310),
.A2(n_300),
.B1(n_290),
.B2(n_291),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_348),
.A2(n_360),
.B1(n_288),
.B2(n_274),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_351),
.Y(n_386)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_294),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_290),
.B(n_302),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_282),
.B(n_278),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_303),
.C(n_297),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_354),
.C(n_362),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_297),
.B(n_303),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_313),
.A2(n_312),
.B1(n_309),
.B2(n_311),
.Y(n_356)
);

OAI21xp33_ASAP7_75t_L g357 ( 
.A1(n_313),
.A2(n_305),
.B(n_317),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_357),
.A2(n_289),
.B(n_279),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_279),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_358),
.Y(n_373)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_286),
.Y(n_359)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_359),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_284),
.A2(n_286),
.B1(n_321),
.B2(n_314),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_321),
.B(n_323),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_288),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_334),
.A2(n_320),
.B(n_319),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_366),
.A2(n_377),
.B(n_335),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_367),
.B(n_389),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_329),
.A2(n_320),
.B(n_319),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_368),
.A2(n_376),
.B(n_336),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_337),
.A2(n_314),
.B1(n_318),
.B2(n_274),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_369),
.A2(n_384),
.B1(n_387),
.B2(n_367),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_SL g397 ( 
.A(n_374),
.B(n_375),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_355),
.A2(n_289),
.B(n_306),
.Y(n_375)
);

NAND2x1_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_318),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_326),
.A2(n_276),
.B1(n_333),
.B2(n_327),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_380),
.A2(n_391),
.B1(n_348),
.B2(n_342),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_326),
.A2(n_329),
.B1(n_324),
.B2(n_338),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_381),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_337),
.A2(n_329),
.B1(n_345),
.B2(n_326),
.Y(n_384)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_387),
.Y(n_394)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_388),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_344),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_390),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_347),
.A2(n_343),
.B1(n_345),
.B2(n_349),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_393),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_395),
.A2(n_400),
.B(n_412),
.Y(n_433)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_377),
.A2(n_353),
.B(n_351),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_399),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_332),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_402),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_385),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_332),
.C(n_341),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_403),
.C(n_419),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_379),
.C(n_392),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_330),
.Y(n_405)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_405),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_385),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_406),
.B(n_378),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_407),
.A2(n_415),
.B1(n_383),
.B2(n_369),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_325),
.Y(n_409)
);

NAND3xp33_ASAP7_75t_L g429 ( 
.A(n_409),
.B(n_410),
.C(n_411),
.Y(n_429)
);

NOR3xp33_ASAP7_75t_SL g410 ( 
.A(n_386),
.B(n_354),
.C(n_346),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_350),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_368),
.A2(n_362),
.B(n_366),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_365),
.Y(n_413)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_413),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_384),
.Y(n_416)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_416),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_372),
.Y(n_417)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_417),
.Y(n_442)
);

OAI21xp33_ASAP7_75t_L g418 ( 
.A1(n_382),
.A2(n_372),
.B(n_368),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_382),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_392),
.B(n_379),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_419),
.B(n_392),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_376),
.A2(n_375),
.B(n_377),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_420),
.A2(n_388),
.B(n_390),
.Y(n_445)
);

XOR2x1_ASAP7_75t_SL g422 ( 
.A(n_397),
.B(n_377),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_422),
.A2(n_426),
.B(n_445),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_424),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_383),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_425),
.B(n_432),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_428),
.A2(n_430),
.B1(n_431),
.B2(n_415),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_416),
.A2(n_371),
.B1(n_381),
.B2(n_374),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_401),
.A2(n_371),
.B1(n_363),
.B2(n_373),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_363),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_435),
.B(n_437),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_411),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_436),
.B(n_399),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_364),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_396),
.B(n_364),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_407),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_396),
.B(n_378),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_446),
.C(n_412),
.Y(n_458)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_443),
.Y(n_465)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_404),
.Y(n_444)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_444),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_396),
.B(n_365),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_406),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_450),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_443),
.B(n_414),
.Y(n_449)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_449),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_414),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_451),
.A2(n_456),
.B1(n_457),
.B2(n_460),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_452),
.A2(n_461),
.B1(n_462),
.B2(n_464),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_427),
.B(n_417),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_455),
.B(n_465),
.Y(n_479)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_442),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_434),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_435),
.Y(n_468)
);

MAJx2_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_433),
.C(n_445),
.Y(n_475)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_431),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_428),
.A2(n_401),
.B1(n_420),
.B2(n_395),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_430),
.A2(n_421),
.B1(n_394),
.B2(n_400),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_440),
.A2(n_427),
.B1(n_441),
.B2(n_446),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_463),
.B(n_425),
.C(n_423),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_467),
.B(n_471),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_475),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_432),
.C(n_437),
.Y(n_471)
);

NOR3xp33_ASAP7_75t_SL g472 ( 
.A(n_457),
.B(n_410),
.C(n_409),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_410),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_439),
.C(n_433),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_474),
.B(n_476),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_466),
.B(n_424),
.C(n_422),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_447),
.B(n_397),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_477),
.B(n_478),
.C(n_458),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_405),
.Y(n_478)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_479),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_464),
.A2(n_394),
.B(n_408),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_480),
.A2(n_449),
.B(n_465),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_481),
.Y(n_482)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_482),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_478),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_469),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_486),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_468),
.C(n_471),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_476),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_490),
.A2(n_480),
.B(n_453),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_473),
.A2(n_460),
.B1(n_454),
.B2(n_450),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_491),
.A2(n_461),
.B1(n_462),
.B2(n_459),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_470),
.Y(n_492)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_492),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_493),
.B(n_456),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_498),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_497),
.B(n_502),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_493),
.B(n_452),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_482),
.A2(n_472),
.B1(n_475),
.B2(n_454),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_501),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_503),
.B(n_504),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_453),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_496),
.A2(n_484),
.B(n_489),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_506),
.A2(n_490),
.B(n_438),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_502),
.A2(n_488),
.B(n_487),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_508),
.A2(n_509),
.B(n_504),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_501),
.A2(n_487),
.B(n_483),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_486),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_510),
.B(n_513),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_500),
.C(n_497),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_515),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_491),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_516),
.B(n_507),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_512),
.B(n_413),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_517),
.B(n_518),
.Y(n_523)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_512),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_519),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_520),
.Y(n_525)
);

NAND4xp25_ASAP7_75t_SL g524 ( 
.A(n_521),
.B(n_511),
.C(n_507),
.D(n_474),
.Y(n_524)
);

AO21x1_ASAP7_75t_L g526 ( 
.A1(n_524),
.A2(n_522),
.B(n_523),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_525),
.B(n_408),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_527),
.B(n_404),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_528),
.Y(n_529)
);


endmodule