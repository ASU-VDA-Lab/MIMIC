module fake_netlist_6_437_n_1921 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1921);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1921;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1669;
wire n_1403;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_87),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_93),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_38),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_39),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_138),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_72),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_27),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_70),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_1),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_106),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_28),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_82),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_110),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_153),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_167),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_183),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_20),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_101),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_49),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_76),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_156),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_22),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_114),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_50),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_103),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_78),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_149),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_20),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_49),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_27),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_141),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_68),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_71),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_120),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_118),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_104),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_173),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_85),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_91),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_44),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_0),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_109),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_19),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_124),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_163),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_65),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_102),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_99),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_151),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_144),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_92),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_111),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_42),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_121),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_142),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_26),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_136),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_79),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_107),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_152),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_143),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_28),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_50),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_16),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_39),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_95),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_42),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_7),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_59),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_6),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_64),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_8),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_112),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_53),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_35),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_97),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_113),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_90),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_73),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_122),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_58),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_17),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_69),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_62),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_31),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_177),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_14),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_137),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_135),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_32),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_66),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_19),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_179),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_37),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_54),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_36),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_2),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_51),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_96),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_133),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_89),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_159),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_11),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_11),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_174),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_115),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_158),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_17),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_29),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_105),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_176),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_15),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_160),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_32),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_40),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_22),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_58),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_43),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_12),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_59),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_148),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_86),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_8),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_48),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_77),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_80),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_10),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_36),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_4),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_84),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_2),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_147),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_139),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_154),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_62),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_161),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_94),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_61),
.Y(n_336)
);

BUFx2_ASAP7_75t_SL g337 ( 
.A(n_116),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_117),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_63),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_169),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_164),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_15),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_21),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_132),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_56),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_24),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_53),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_23),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_38),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_126),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_10),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_26),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_6),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_51),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_67),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_166),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_157),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_74),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_134),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_33),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_45),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_47),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_5),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_5),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_150),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_3),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_57),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_234),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_211),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_235),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_212),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_249),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_312),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_222),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_259),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_367),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_218),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_248),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_262),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_0),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_264),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_188),
.B(n_1),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_188),
.B(n_3),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_286),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_367),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_265),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_267),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_278),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_287),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_227),
.B(n_7),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_282),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_292),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_187),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_208),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_240),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_294),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_190),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_242),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_227),
.B(n_9),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_213),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_291),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_215),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_220),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_238),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_260),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_293),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_198),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_302),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_260),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_307),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_243),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_331),
.B(n_217),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_252),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_310),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_314),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_246),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_186),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_261),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_266),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_271),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_247),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_272),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_186),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_192),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_281),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_201),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_290),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_192),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_295),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_217),
.B(n_9),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_296),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_197),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_306),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_322),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_250),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_201),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_329),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_197),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_206),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_346),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_347),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_349),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_198),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_206),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_209),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_351),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_245),
.B(n_12),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_209),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_291),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_207),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_291),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_221),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_233),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_245),
.B(n_13),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_364),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_458),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_369),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_399),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_400),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_458),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_433),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_403),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_458),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_416),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_458),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_381),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_458),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_372),
.A2(n_313),
.B1(n_342),
.B2(n_279),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_412),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_422),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_R g477 ( 
.A(n_421),
.B(n_253),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_378),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_426),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_440),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_417),
.B(n_184),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_448),
.B(n_207),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_382),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_368),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_393),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_371),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_371),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

CKINVDCx8_ASAP7_75t_R g490 ( 
.A(n_431),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_374),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_406),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_454),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_454),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_441),
.B(n_201),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_456),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_422),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_433),
.Y(n_498)
);

AND2x2_ASAP7_75t_SL g499 ( 
.A(n_452),
.B(n_273),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_455),
.B(n_244),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_455),
.B(n_184),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_374),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_398),
.Y(n_503)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_446),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_456),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

CKINVDCx8_ASAP7_75t_R g508 ( 
.A(n_410),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_459),
.A2(n_284),
.B(n_219),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_R g510 ( 
.A(n_377),
.B(n_383),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_377),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_455),
.B(n_244),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_373),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_408),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_386),
.B(n_185),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_387),
.B(n_185),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_412),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_379),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_384),
.B(n_311),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_380),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_395),
.B(n_404),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_383),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_385),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_418),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_423),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_385),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_424),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_390),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_390),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_425),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_411),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_391),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_430),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_432),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_478),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_504),
.B(n_392),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_499),
.B(n_273),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_523),
.B(n_376),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_503),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_475),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_475),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_521),
.A2(n_388),
.B1(n_394),
.B2(n_392),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_475),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_521),
.B(n_523),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_481),
.B(n_396),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_503),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_468),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_478),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_519),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_519),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_499),
.B(n_299),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_481),
.B(n_396),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_505),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_478),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_477),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_533),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_499),
.B(n_397),
.Y(n_560)
);

BUFx6f_ASAP7_75t_SL g561 ( 
.A(n_519),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_462),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_513),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_517),
.B(n_397),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_500),
.B(n_401),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_505),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_493),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_533),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_483),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_507),
.Y(n_570)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_466),
.B(n_420),
.C(n_413),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_513),
.B(n_299),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_509),
.A2(n_435),
.B1(n_366),
.B2(n_325),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_513),
.B(n_233),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_507),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_493),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_500),
.B(n_401),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_493),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_517),
.A2(n_429),
.B1(n_457),
.B2(n_453),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_493),
.Y(n_580)
);

INVx4_ASAP7_75t_SL g581 ( 
.A(n_493),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_468),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_514),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_513),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_500),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_518),
.B(n_233),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_482),
.B(n_285),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_468),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_482),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_483),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_482),
.B(n_370),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_518),
.B(n_413),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_468),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_466),
.B(n_415),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_501),
.B(n_415),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_501),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_512),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_509),
.A2(n_366),
.B1(n_325),
.B2(n_219),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_SL g599 ( 
.A(n_495),
.B(n_221),
.Y(n_599)
);

INVx4_ASAP7_75t_SL g600 ( 
.A(n_493),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_468),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_512),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_468),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_468),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_469),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_515),
.B(n_375),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_465),
.B(n_419),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_520),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_494),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_483),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_498),
.B(n_337),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_509),
.A2(n_288),
.B1(n_284),
.B2(n_338),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_484),
.B(n_233),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_465),
.B(n_285),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_509),
.A2(n_288),
.B1(n_297),
.B2(n_334),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_494),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_485),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_476),
.B(n_428),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_487),
.B(n_428),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_494),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_515),
.B(n_434),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_516),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_522),
.Y(n_624)
);

BUFx10_ASAP7_75t_L g625 ( 
.A(n_488),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_485),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_465),
.B(n_297),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_494),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_485),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_489),
.Y(n_630)
);

BUFx10_ASAP7_75t_L g631 ( 
.A(n_491),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_526),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_465),
.B(n_339),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_526),
.B(n_529),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_476),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_529),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_489),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_532),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_502),
.B(n_233),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_471),
.B(n_255),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_532),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_486),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_489),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_471),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_492),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_511),
.B(n_304),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_492),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_527),
.B(n_436),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_524),
.B(n_429),
.Y(n_649)
);

CKINVDCx16_ASAP7_75t_R g650 ( 
.A(n_510),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_525),
.B(n_437),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_528),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_497),
.A2(n_444),
.B1(n_457),
.B2(n_453),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_461),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_530),
.B(n_304),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_486),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_473),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_496),
.B(n_304),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_496),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_527),
.B(n_438),
.Y(n_660)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_461),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_531),
.A2(n_420),
.B1(n_450),
.B2(n_449),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_497),
.B(n_437),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_461),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_473),
.Y(n_665)
);

INVxp67_ASAP7_75t_SL g666 ( 
.A(n_470),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_527),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_534),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_534),
.B(n_439),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_535),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_474),
.B(n_317),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_496),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_506),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_506),
.B(n_256),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_470),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_534),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_536),
.A2(n_460),
.B1(n_451),
.B2(n_447),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_506),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_536),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_536),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_470),
.B(n_257),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_537),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_537),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_SL g684 ( 
.A1(n_474),
.A2(n_277),
.B1(n_318),
.B2(n_326),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_472),
.B(n_258),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_559),
.B(n_443),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_547),
.B(n_443),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_543),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_543),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_585),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_585),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_544),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_596),
.B(n_589),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_540),
.A2(n_269),
.B1(n_321),
.B2(n_304),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_558),
.B(n_464),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_596),
.B(n_472),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_637),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_563),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_563),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_541),
.B(n_490),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_584),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_592),
.B(n_490),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_589),
.B(n_472),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_564),
.B(n_193),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_548),
.B(n_194),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_555),
.B(n_196),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_560),
.B(n_490),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_595),
.B(n_565),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_577),
.B(n_199),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_584),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_644),
.B(n_200),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_568),
.B(n_304),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_591),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_637),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_635),
.B(n_414),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_540),
.B(n_291),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_558),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_644),
.B(n_210),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_579),
.A2(n_309),
.B1(n_274),
.B2(n_275),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_637),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_616),
.B(n_216),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_635),
.B(n_650),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_591),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_554),
.A2(n_283),
.B1(n_276),
.B2(n_289),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_554),
.B(n_291),
.Y(n_725)
);

OR2x6_ASAP7_75t_L g726 ( 
.A(n_583),
.B(n_670),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_632),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_587),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_632),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_613),
.B(n_225),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_542),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_587),
.B(n_228),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_549),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_587),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_562),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_539),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_657),
.B(n_231),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_556),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_594),
.B(n_508),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_622),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_634),
.B(n_601),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_665),
.B(n_236),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_546),
.B(n_237),
.Y(n_743)
);

NOR2xp67_ASAP7_75t_L g744 ( 
.A(n_571),
.B(n_467),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_544),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_634),
.B(n_291),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_672),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_634),
.B(n_291),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_546),
.B(n_239),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_553),
.B(n_659),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_601),
.B(n_617),
.Y(n_751)
);

OAI221xp5_ASAP7_75t_L g752 ( 
.A1(n_684),
.A2(n_537),
.B1(n_445),
.B2(n_442),
.C(n_365),
.Y(n_752)
);

NOR3xp33_ASAP7_75t_L g753 ( 
.A(n_653),
.B(n_241),
.C(n_251),
.Y(n_753)
);

BUFx4f_ASAP7_75t_L g754 ( 
.A(n_612),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_620),
.B(n_479),
.C(n_480),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_601),
.B(n_291),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_553),
.B(n_659),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_566),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_570),
.Y(n_759)
);

OAI22xp33_ASAP7_75t_L g760 ( 
.A1(n_671),
.A2(n_352),
.B1(n_363),
.B2(n_362),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_575),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_630),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_630),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_659),
.B(n_254),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_678),
.B(n_263),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_678),
.B(n_268),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_599),
.A2(n_300),
.B1(n_303),
.B2(n_305),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_597),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_552),
.B(n_270),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_603),
.Y(n_770)
);

BUFx5_ASAP7_75t_L g771 ( 
.A(n_658),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_670),
.B(n_508),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_573),
.A2(n_598),
.B1(n_586),
.B2(n_671),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_586),
.A2(n_280),
.B(n_355),
.C(n_298),
.Y(n_774)
);

CKINVDCx6p67_ASAP7_75t_R g775 ( 
.A(n_625),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_617),
.B(n_508),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_678),
.B(n_308),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_612),
.B(n_324),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_672),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_623),
.B(n_335),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_675),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_672),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_614),
.B(n_189),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_L g784 ( 
.A1(n_671),
.A2(n_327),
.B1(n_363),
.B2(n_362),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_578),
.A2(n_666),
.B(n_661),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_608),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_614),
.B(n_189),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_636),
.B(n_341),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_619),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_638),
.B(n_359),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_617),
.B(n_191),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_639),
.B(n_646),
.Y(n_792)
);

OAI22xp33_ASAP7_75t_L g793 ( 
.A1(n_671),
.A2(n_326),
.B1(n_361),
.B2(n_360),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_610),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_562),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_641),
.B(n_191),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_621),
.B(n_195),
.Y(n_797)
);

BUFx8_ASAP7_75t_L g798 ( 
.A(n_561),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_621),
.B(n_195),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_622),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_612),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_660),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_621),
.B(n_674),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_660),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_642),
.B(n_202),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_610),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_607),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_599),
.A2(n_327),
.B(n_361),
.C(n_360),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_656),
.B(n_202),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_649),
.B(n_463),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_619),
.B(n_315),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_572),
.A2(n_318),
.B1(n_315),
.B2(n_316),
.Y(n_812)
);

INVx4_ASAP7_75t_L g813 ( 
.A(n_628),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_607),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_572),
.A2(n_358),
.B(n_357),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_663),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_663),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_648),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_633),
.B(n_203),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_640),
.B(n_204),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_643),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_667),
.B(n_204),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_668),
.B(n_205),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_676),
.B(n_205),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_648),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_639),
.B(n_214),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_679),
.B(n_214),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_680),
.B(n_223),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_612),
.A2(n_358),
.B1(n_357),
.B2(n_356),
.Y(n_829)
);

AND2x6_ASAP7_75t_L g830 ( 
.A(n_645),
.B(n_277),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_682),
.B(n_223),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_683),
.B(n_224),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_545),
.B(n_662),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_648),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_646),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_675),
.B(n_224),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_654),
.B(n_664),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_681),
.B(n_226),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_685),
.B(n_226),
.Y(n_839)
);

BUFx8_ASAP7_75t_L g840 ( 
.A(n_561),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_645),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_574),
.B(n_229),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_651),
.B(n_316),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_647),
.Y(n_844)
);

INVx8_ASAP7_75t_L g845 ( 
.A(n_561),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_669),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_654),
.Y(n_847)
);

NOR2xp67_ASAP7_75t_SL g848 ( 
.A(n_582),
.B(n_229),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_574),
.B(n_230),
.Y(n_849)
);

BUFx6f_ASAP7_75t_SL g850 ( 
.A(n_625),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_655),
.A2(n_356),
.B(n_232),
.C(n_319),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_567),
.B(n_230),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_647),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_687),
.A2(n_615),
.B(n_627),
.C(n_669),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_701),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_818),
.Y(n_856)
);

BUFx12f_ASAP7_75t_L g857 ( 
.A(n_798),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_785),
.A2(n_602),
.B(n_593),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_837),
.A2(n_602),
.B(n_593),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_708),
.A2(n_590),
.B(n_557),
.C(n_551),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_740),
.B(n_669),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_750),
.A2(n_576),
.B(n_580),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_715),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_701),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_773),
.A2(n_580),
.B1(n_567),
.B2(n_576),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_756),
.A2(n_673),
.B(n_567),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_762),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_757),
.A2(n_580),
.B(n_576),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_707),
.A2(n_624),
.B1(n_609),
.B2(n_631),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_800),
.B(n_625),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_800),
.B(n_550),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_741),
.A2(n_602),
.B(n_593),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_686),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_687),
.A2(n_323),
.B1(n_350),
.B2(n_320),
.Y(n_874)
);

BUFx12f_ASAP7_75t_L g875 ( 
.A(n_798),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_816),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_792),
.A2(n_557),
.B(n_569),
.C(n_551),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_803),
.A2(n_741),
.B(n_837),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_693),
.B(n_550),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_704),
.B(n_705),
.Y(n_880)
);

OAI321xp33_ASAP7_75t_L g881 ( 
.A1(n_760),
.A2(n_677),
.A3(n_354),
.B1(n_353),
.B2(n_333),
.C(n_336),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_792),
.A2(n_330),
.B1(n_320),
.B2(n_323),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_781),
.A2(n_582),
.B(n_588),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_781),
.A2(n_582),
.B(n_588),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_835),
.A2(n_340),
.B1(n_328),
.B2(n_344),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_716),
.A2(n_550),
.B(n_590),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_762),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_730),
.A2(n_588),
.B(n_604),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_688),
.B(n_606),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_L g890 ( 
.A(n_760),
.B(n_340),
.C(n_350),
.Y(n_890)
);

AND3x2_ASAP7_75t_L g891 ( 
.A(n_801),
.B(n_652),
.C(n_631),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_745),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_736),
.B(n_631),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_736),
.B(n_652),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_716),
.A2(n_569),
.B(n_611),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_703),
.A2(n_604),
.B(n_605),
.Y(n_896)
);

NOR2x1p5_ASAP7_75t_L g897 ( 
.A(n_775),
.B(n_333),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_706),
.B(n_654),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_700),
.B(n_652),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_789),
.B(n_654),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_721),
.A2(n_605),
.B(n_628),
.Y(n_901)
);

OAI21xp33_ASAP7_75t_L g902 ( 
.A1(n_700),
.A2(n_352),
.B(n_336),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_825),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_786),
.B(n_664),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_728),
.A2(n_734),
.B1(n_707),
.B2(n_694),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_763),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_690),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_SL g908 ( 
.A1(n_725),
.A2(n_748),
.B(n_746),
.C(n_791),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_745),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_802),
.A2(n_538),
.B(n_629),
.C(n_626),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_696),
.A2(n_605),
.B(n_628),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_753),
.A2(n_538),
.B1(n_611),
.B2(n_618),
.Y(n_912)
);

BUFx12f_ASAP7_75t_L g913 ( 
.A(n_840),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_804),
.A2(n_626),
.B(n_658),
.C(n_277),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_732),
.A2(n_605),
.B(n_628),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_799),
.A2(n_605),
.B(n_628),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_691),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_745),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_764),
.A2(n_664),
.B(n_581),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_709),
.B(n_664),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_783),
.A2(n_328),
.B(n_344),
.C(n_354),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_765),
.A2(n_600),
.B(n_581),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_SL g923 ( 
.A1(n_746),
.A2(n_748),
.B(n_797),
.C(n_791),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_766),
.A2(n_600),
.B(n_581),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_713),
.B(n_600),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_834),
.Y(n_926)
);

CKINVDCx10_ASAP7_75t_R g927 ( 
.A(n_850),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_777),
.A2(n_658),
.B(n_353),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_847),
.A2(n_600),
.B(n_581),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_847),
.A2(n_852),
.B(n_806),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_845),
.B(n_13),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_723),
.B(n_731),
.Y(n_932)
);

NOR3xp33_ASAP7_75t_L g933 ( 
.A(n_784),
.B(n_348),
.C(n_345),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_821),
.Y(n_934)
);

AOI21x1_ASAP7_75t_L g935 ( 
.A1(n_743),
.A2(n_658),
.B(n_129),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_783),
.A2(n_348),
.B(n_345),
.C(n_343),
.Y(n_936)
);

AO22x1_ASAP7_75t_L g937 ( 
.A1(n_753),
.A2(n_343),
.B1(n_658),
.B2(n_18),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_846),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_694),
.A2(n_658),
.B1(n_16),
.B2(n_18),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_745),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_733),
.B(n_14),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_738),
.B(n_21),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_847),
.A2(n_181),
.B(n_172),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_759),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_789),
.B(n_23),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_L g946 ( 
.A(n_784),
.B(n_24),
.C(n_25),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_847),
.A2(n_168),
.B(n_146),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_787),
.A2(n_25),
.B(n_29),
.C(n_30),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_768),
.B(n_30),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_770),
.B(n_31),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_819),
.B(n_33),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_794),
.A2(n_145),
.B(n_140),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_807),
.B(n_34),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_814),
.B(n_34),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_769),
.B(n_35),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_749),
.A2(n_838),
.B(n_839),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_722),
.B(n_128),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_833),
.A2(n_125),
.B1(n_119),
.B2(n_100),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_836),
.A2(n_88),
.B(n_83),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_702),
.A2(n_81),
.B1(n_75),
.B2(n_41),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_SL g961 ( 
.A1(n_752),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_698),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_845),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_817),
.B(n_702),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_SL g965 ( 
.A1(n_797),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_820),
.A2(n_46),
.B(n_47),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_769),
.B(n_46),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_787),
.B(n_48),
.Y(n_968)
);

AO22x1_ASAP7_75t_L g969 ( 
.A1(n_826),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_969)
);

CKINVDCx11_ASAP7_75t_R g970 ( 
.A(n_726),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_699),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_697),
.A2(n_57),
.B(n_60),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_714),
.A2(n_60),
.B(n_61),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_739),
.B(n_754),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_808),
.A2(n_793),
.B(n_718),
.C(n_711),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_735),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_720),
.A2(n_779),
.B(n_747),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_795),
.Y(n_978)
);

OAI321xp33_ASAP7_75t_L g979 ( 
.A1(n_793),
.A2(n_812),
.A3(n_826),
.B1(n_808),
.B2(n_843),
.C(n_811),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_754),
.B(n_758),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_841),
.A2(n_853),
.B(n_844),
.Y(n_981)
);

NAND2x1p5_ASAP7_75t_L g982 ( 
.A(n_688),
.B(n_689),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_782),
.A2(n_710),
.B(n_727),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_729),
.B(n_758),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_761),
.B(n_776),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_761),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_737),
.A2(n_742),
.B(n_780),
.C(n_790),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_689),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_L g989 ( 
.A(n_755),
.B(n_772),
.C(n_801),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_813),
.A2(n_831),
.B(n_828),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_842),
.A2(n_849),
.B(n_815),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_692),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_692),
.A2(n_776),
.B1(n_724),
.B2(n_829),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_813),
.A2(n_824),
.B(n_822),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_796),
.A2(n_809),
.B(n_805),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_827),
.A2(n_832),
.B(n_788),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_823),
.A2(n_712),
.B(n_851),
.C(n_774),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_712),
.B(n_823),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_719),
.A2(n_767),
.B(n_744),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_717),
.B(n_778),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_778),
.A2(n_810),
.B(n_726),
.C(n_695),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_845),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_778),
.A2(n_726),
.B1(n_850),
.B2(n_848),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_830),
.A2(n_547),
.B(n_554),
.C(n_540),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_771),
.A2(n_830),
.B(n_840),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_771),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_771),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_771),
.A2(n_757),
.B(n_750),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_771),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_830),
.Y(n_1010)
);

AO22x1_ASAP7_75t_L g1011 ( 
.A1(n_687),
.A2(n_547),
.B1(n_700),
.B2(n_707),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_762),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_708),
.A2(n_547),
.B1(n_707),
.B2(n_792),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_708),
.B(n_559),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_687),
.A2(n_547),
.B(n_792),
.C(n_564),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_750),
.A2(n_757),
.B(n_751),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_818),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_708),
.B(n_547),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_750),
.A2(n_757),
.B(n_751),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_708),
.B(n_547),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_686),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_687),
.B(n_547),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_708),
.B(n_547),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_701),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_750),
.A2(n_757),
.B(n_751),
.Y(n_1025)
);

INVx11_ASAP7_75t_L g1026 ( 
.A(n_798),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_SL g1027 ( 
.A(n_717),
.B(n_559),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_773),
.A2(n_547),
.B1(n_800),
.B2(n_740),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_687),
.B(n_547),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_708),
.B(n_547),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_750),
.A2(n_757),
.B(n_751),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_708),
.B(n_547),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_750),
.A2(n_757),
.B(n_751),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_740),
.B(n_559),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_762),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_SL g1036 ( 
.A(n_889),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1034),
.B(n_1022),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_1022),
.B(n_1029),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_988),
.B(n_980),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_1029),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_867),
.Y(n_1041)
);

AOI21x1_ASAP7_75t_L g1042 ( 
.A1(n_865),
.A2(n_1019),
.B(n_1016),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_SL g1043 ( 
.A1(n_961),
.A2(n_976),
.B1(n_931),
.B2(n_869),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_859),
.A2(n_858),
.B(n_981),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_983),
.A2(n_878),
.B(n_1025),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_887),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_892),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1018),
.B(n_1020),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1031),
.A2(n_1033),
.B(n_923),
.Y(n_1049)
);

NOR2x1_ASAP7_75t_SL g1050 ( 
.A(n_892),
.B(n_909),
.Y(n_1050)
);

OAI22x1_ASAP7_75t_L g1051 ( 
.A1(n_1013),
.A2(n_964),
.B1(n_945),
.B2(n_870),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1023),
.B(n_1030),
.Y(n_1052)
);

AOI21xp33_ASAP7_75t_L g1053 ( 
.A1(n_999),
.A2(n_979),
.B(n_1028),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_1032),
.A2(n_1004),
.B(n_939),
.C(n_968),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_939),
.A2(n_881),
.B(n_975),
.C(n_880),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_876),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_1008),
.A2(n_930),
.B(n_910),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_SL g1058 ( 
.A1(n_854),
.A2(n_861),
.B(n_993),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1011),
.B(n_964),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_1014),
.A2(n_936),
.B(n_948),
.C(n_921),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_905),
.A2(n_991),
.B1(n_863),
.B2(n_998),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_876),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_892),
.Y(n_1063)
);

OAI22x1_ASAP7_75t_L g1064 ( 
.A1(n_945),
.A2(n_894),
.B1(n_974),
.B2(n_899),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_975),
.A2(n_961),
.B(n_890),
.C(n_933),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_906),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_908),
.A2(n_898),
.B(n_920),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_SL g1068 ( 
.A1(n_951),
.A2(n_967),
.B(n_955),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_890),
.A2(n_933),
.B(n_946),
.C(n_902),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_863),
.B(n_995),
.Y(n_1070)
);

AND2x4_ASAP7_75t_SL g1071 ( 
.A(n_1002),
.B(n_963),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_855),
.B(n_864),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_889),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_873),
.B(n_1021),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_895),
.A2(n_886),
.B(n_872),
.Y(n_1075)
);

AO21x1_ASAP7_75t_L g1076 ( 
.A1(n_997),
.A2(n_985),
.B(n_960),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_892),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_988),
.B(n_963),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_1002),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1012),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_944),
.B(n_900),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_978),
.B(n_932),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_907),
.B(n_917),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_1002),
.B(n_986),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_1027),
.B(n_984),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_856),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_903),
.B(n_926),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_877),
.A2(n_860),
.B(n_996),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_938),
.B(n_1017),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_990),
.A2(n_994),
.B(n_868),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_871),
.A2(n_855),
.B1(n_1024),
.B2(n_864),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_909),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_866),
.A2(n_862),
.B(n_860),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_879),
.A2(n_987),
.B(n_997),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1035),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_919),
.A2(n_888),
.B(n_916),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_989),
.B(n_894),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_989),
.B(n_1000),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_946),
.A2(n_966),
.B(n_954),
.C(n_953),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_904),
.B(n_962),
.Y(n_1100)
);

AND2x2_ASAP7_75t_SL g1101 ( 
.A(n_909),
.B(n_918),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_896),
.A2(n_1010),
.B(n_924),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1010),
.A2(n_922),
.B(n_977),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1024),
.B(n_942),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_883),
.A2(n_884),
.B(n_987),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_911),
.A2(n_929),
.B(n_901),
.Y(n_1106)
);

AOI221x1_ASAP7_75t_L g1107 ( 
.A1(n_972),
.A2(n_973),
.B1(n_941),
.B2(n_950),
.C(n_949),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_934),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_909),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_SL g1110 ( 
.A1(n_918),
.A2(n_1005),
.B(n_957),
.Y(n_1110)
);

OAI22x1_ASAP7_75t_L g1111 ( 
.A1(n_893),
.A2(n_1000),
.B1(n_992),
.B2(n_982),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_935),
.A2(n_915),
.B(n_956),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1006),
.A2(n_1007),
.B(n_1009),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_912),
.A2(n_928),
.B(n_925),
.Y(n_1114)
);

NAND2xp33_ASAP7_75t_SL g1115 ( 
.A(n_1002),
.B(n_918),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_940),
.A2(n_918),
.B(n_959),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_882),
.A2(n_914),
.B(n_940),
.Y(n_1117)
);

OAI22x1_ASAP7_75t_L g1118 ( 
.A1(n_982),
.A2(n_897),
.B1(n_969),
.B2(n_970),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_958),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_914),
.A2(n_952),
.B(n_947),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_943),
.A2(n_1001),
.B(n_965),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_931),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_874),
.B(n_885),
.Y(n_1123)
);

OAI211xp5_ASAP7_75t_L g1124 ( 
.A1(n_1001),
.A2(n_971),
.B(n_1003),
.C(n_937),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_931),
.B(n_891),
.Y(n_1125)
);

BUFx12f_ASAP7_75t_L g1126 ( 
.A(n_857),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_891),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1026),
.A2(n_875),
.B(n_913),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_927),
.A2(n_859),
.B(n_983),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1022),
.B(n_1029),
.Y(n_1130)
);

AOI21x1_ASAP7_75t_L g1131 ( 
.A1(n_865),
.A2(n_756),
.B(n_1016),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_859),
.A2(n_983),
.B(n_878),
.Y(n_1132)
);

BUFx8_ASAP7_75t_SL g1133 ( 
.A(n_857),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_859),
.A2(n_983),
.B(n_878),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1016),
.A2(n_751),
.B(n_1031),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_1022),
.Y(n_1136)
);

OA21x2_ASAP7_75t_L g1137 ( 
.A1(n_983),
.A2(n_877),
.B(n_878),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1022),
.B(n_1029),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_892),
.Y(n_1139)
);

BUFx4f_ASAP7_75t_L g1140 ( 
.A(n_1002),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_SL g1141 ( 
.A(n_1027),
.B(n_559),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_1022),
.Y(n_1142)
);

NAND2x1p5_ASAP7_75t_L g1143 ( 
.A(n_892),
.B(n_909),
.Y(n_1143)
);

AO21x2_ASAP7_75t_L g1144 ( 
.A1(n_1015),
.A2(n_878),
.B(n_1016),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_SL g1145 ( 
.A1(n_1005),
.A2(n_999),
.B(n_1001),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1016),
.A2(n_751),
.B(n_1031),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1022),
.B(n_1029),
.Y(n_1147)
);

AOI21x1_ASAP7_75t_L g1148 ( 
.A1(n_865),
.A2(n_756),
.B(n_1016),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1016),
.A2(n_751),
.B(n_1031),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_SL g1150 ( 
.A1(n_1005),
.A2(n_999),
.B(n_1001),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_988),
.B(n_728),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_859),
.A2(n_983),
.B(n_878),
.Y(n_1152)
);

AOI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_1022),
.A2(n_1029),
.B(n_547),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1034),
.B(n_559),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_1022),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_1022),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1022),
.A2(n_1029),
.B(n_547),
.C(n_1015),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_859),
.A2(n_983),
.B(n_878),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_859),
.A2(n_858),
.B(n_981),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_944),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1034),
.B(n_559),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_859),
.A2(n_983),
.B(n_878),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_867),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_859),
.A2(n_983),
.B(n_878),
.Y(n_1164)
);

AO21x2_ASAP7_75t_L g1165 ( 
.A1(n_1015),
.A2(n_878),
.B(n_1016),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_1015),
.A2(n_1028),
.A3(n_1029),
.B(n_1022),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_859),
.A2(n_983),
.B(n_878),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_1022),
.Y(n_1168)
);

BUFx2_ASAP7_75t_SL g1169 ( 
.A(n_1002),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1015),
.A2(n_1028),
.A3(n_1029),
.B(n_1022),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1022),
.B(n_1029),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_859),
.A2(n_983),
.B(n_878),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_944),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_859),
.A2(n_983),
.B(n_878),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_1022),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_859),
.A2(n_983),
.B(n_878),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1022),
.A2(n_1029),
.B(n_547),
.C(n_1015),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1034),
.B(n_559),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_1022),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1022),
.A2(n_1029),
.B1(n_1015),
.B2(n_1020),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1016),
.A2(n_751),
.B(n_1031),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1016),
.A2(n_751),
.B(n_1031),
.Y(n_1182)
);

NAND3xp33_ASAP7_75t_L g1183 ( 
.A(n_1022),
.B(n_1029),
.C(n_547),
.Y(n_1183)
);

OAI21xp33_ASAP7_75t_L g1184 ( 
.A1(n_1022),
.A2(n_1029),
.B(n_547),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_1027),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_867),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_859),
.A2(n_983),
.B(n_878),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1022),
.B(n_1029),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1016),
.A2(n_751),
.B(n_1031),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1022),
.A2(n_1029),
.B1(n_1015),
.B2(n_1020),
.Y(n_1190)
);

OAI22x1_ASAP7_75t_L g1191 ( 
.A1(n_1022),
.A2(n_1029),
.B1(n_687),
.B2(n_1013),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_867),
.Y(n_1192)
);

OA22x2_ASAP7_75t_L g1193 ( 
.A1(n_1013),
.A2(n_671),
.B1(n_789),
.B2(n_816),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1038),
.B(n_1130),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1049),
.A2(n_1058),
.B(n_1135),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1038),
.A2(n_1184),
.B1(n_1141),
.B2(n_1183),
.Y(n_1196)
);

NOR2x1_ASAP7_75t_R g1197 ( 
.A(n_1126),
.B(n_1169),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1154),
.B(n_1161),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1062),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1178),
.B(n_1037),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1041),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1160),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1062),
.Y(n_1203)
);

OAI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1138),
.A2(n_1171),
.B1(n_1188),
.B2(n_1147),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1173),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1048),
.B(n_1052),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1059),
.B(n_1070),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1056),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1071),
.B(n_1079),
.Y(n_1209)
);

CKINVDCx11_ASAP7_75t_R g1210 ( 
.A(n_1126),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1146),
.A2(n_1181),
.B(n_1149),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1086),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1133),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1074),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1087),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1153),
.B(n_1157),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1133),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1078),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1157),
.B(n_1177),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1182),
.A2(n_1189),
.B(n_1090),
.Y(n_1220)
);

AOI21xp33_ASAP7_75t_L g1221 ( 
.A1(n_1191),
.A2(n_1180),
.B(n_1190),
.Y(n_1221)
);

AOI222xp33_ASAP7_75t_L g1222 ( 
.A1(n_1043),
.A2(n_1177),
.B1(n_1065),
.B2(n_1040),
.C1(n_1155),
.C2(n_1179),
.Y(n_1222)
);

AOI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1131),
.A2(n_1148),
.B(n_1105),
.Y(n_1223)
);

AO21x2_ASAP7_75t_L g1224 ( 
.A1(n_1053),
.A2(n_1150),
.B(n_1145),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1140),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1071),
.B(n_1079),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1166),
.B(n_1170),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1067),
.A2(n_1094),
.B(n_1088),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1082),
.B(n_1073),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1098),
.B(n_1185),
.Y(n_1230)
);

BUFx12f_ASAP7_75t_L g1231 ( 
.A(n_1122),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1089),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1136),
.A2(n_1156),
.B(n_1168),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1046),
.Y(n_1234)
);

NOR2x1_ASAP7_75t_SL g1235 ( 
.A(n_1109),
.B(n_1081),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1085),
.A2(n_1097),
.B1(n_1193),
.B2(n_1051),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1166),
.B(n_1170),
.Y(n_1237)
);

OR2x6_ASAP7_75t_L g1238 ( 
.A(n_1039),
.B(n_1078),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1193),
.A2(n_1123),
.B1(n_1175),
.B2(n_1142),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1085),
.B(n_1039),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1166),
.B(n_1170),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1066),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1101),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1144),
.A2(n_1165),
.B(n_1114),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1140),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1166),
.B(n_1170),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1066),
.Y(n_1247)
);

AOI222xp33_ASAP7_75t_L g1248 ( 
.A1(n_1065),
.A2(n_1055),
.B1(n_1069),
.B2(n_1118),
.C1(n_1061),
.C2(n_1054),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1116),
.A2(n_1110),
.B(n_1144),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1080),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1039),
.B(n_1083),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1151),
.B(n_1069),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1119),
.A2(n_1076),
.B1(n_1064),
.B2(n_1036),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1100),
.B(n_1108),
.Y(n_1254)
);

BUFx12f_ASAP7_75t_L g1255 ( 
.A(n_1125),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1165),
.A2(n_1054),
.B(n_1093),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1080),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1055),
.A2(n_1119),
.B1(n_1101),
.B2(n_1099),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1151),
.A2(n_1111),
.B1(n_1104),
.B2(n_1095),
.Y(n_1259)
);

INVx5_ASAP7_75t_L g1260 ( 
.A(n_1063),
.Y(n_1260)
);

BUFx12f_ASAP7_75t_L g1261 ( 
.A(n_1084),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1163),
.Y(n_1262)
);

AOI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1121),
.A2(n_1042),
.B(n_1044),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1084),
.B(n_1151),
.Y(n_1264)
);

CKINVDCx11_ASAP7_75t_R g1265 ( 
.A(n_1127),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1093),
.A2(n_1045),
.B(n_1057),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1127),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1092),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1084),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1072),
.A2(n_1192),
.B1(n_1186),
.B2(n_1163),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1063),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1099),
.A2(n_1060),
.B(n_1124),
.C(n_1117),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1186),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1192),
.B(n_1092),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1063),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1109),
.B(n_1139),
.Y(n_1276)
);

AO21x2_ASAP7_75t_L g1277 ( 
.A1(n_1045),
.A2(n_1112),
.B(n_1158),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1063),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1072),
.A2(n_1091),
.B1(n_1139),
.B2(n_1047),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1047),
.B(n_1077),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1077),
.B(n_1107),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1143),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1143),
.B(n_1050),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1109),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1113),
.B(n_1109),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1115),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1129),
.Y(n_1287)
);

AOI21xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1129),
.A2(n_1120),
.B(n_1128),
.Y(n_1288)
);

AND2x6_ASAP7_75t_L g1289 ( 
.A(n_1115),
.B(n_1068),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1137),
.A2(n_1075),
.B1(n_1057),
.B2(n_1120),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1137),
.B(n_1102),
.Y(n_1291)
);

INVx5_ASAP7_75t_L g1292 ( 
.A(n_1102),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1106),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1103),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1103),
.Y(n_1295)
);

AOI221xp5_ASAP7_75t_L g1296 ( 
.A1(n_1132),
.A2(n_1162),
.B1(n_1176),
.B2(n_1174),
.C(n_1134),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1106),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1112),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1096),
.A2(n_1134),
.B1(n_1152),
.B2(n_1187),
.Y(n_1299)
);

OR2x6_ASAP7_75t_SL g1300 ( 
.A(n_1096),
.B(n_1152),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1162),
.A2(n_1164),
.B(n_1167),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1164),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1167),
.B(n_1172),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1187),
.B(n_1172),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1174),
.B(n_1176),
.Y(n_1305)
);

BUFx10_ASAP7_75t_L g1306 ( 
.A(n_1159),
.Y(n_1306)
);

INVx4_ASAP7_75t_L g1307 ( 
.A(n_1140),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1154),
.B(n_1161),
.Y(n_1308)
);

BUFx12f_ASAP7_75t_L g1309 ( 
.A(n_1126),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1153),
.B(n_1022),
.Y(n_1310)
);

CKINVDCx8_ASAP7_75t_R g1311 ( 
.A(n_1169),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1154),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1049),
.A2(n_1058),
.B(n_1135),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1038),
.B(n_1130),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1056),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1154),
.B(n_1161),
.Y(n_1316)
);

OAI321xp33_ASAP7_75t_L g1317 ( 
.A1(n_1184),
.A2(n_1029),
.A3(n_1022),
.B1(n_1183),
.B2(n_1038),
.C(n_1138),
.Y(n_1317)
);

NAND2x1p5_ASAP7_75t_L g1318 ( 
.A(n_1109),
.B(n_1101),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1160),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1049),
.A2(n_1058),
.B(n_1135),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1154),
.B(n_1161),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_SL g1322 ( 
.A(n_1184),
.B(n_1029),
.Y(n_1322)
);

NAND2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1109),
.B(n_1101),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1154),
.B(n_1161),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1160),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1071),
.B(n_1079),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1056),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1154),
.B(n_1161),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1078),
.Y(n_1329)
);

OR2x6_ASAP7_75t_L g1330 ( 
.A(n_1169),
.B(n_1002),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1062),
.Y(n_1331)
);

AND2x6_ASAP7_75t_L g1332 ( 
.A(n_1119),
.B(n_1063),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1038),
.B(n_1130),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1038),
.A2(n_1029),
.B(n_1022),
.C(n_1015),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1038),
.A2(n_1029),
.B1(n_1022),
.B2(n_1130),
.Y(n_1335)
);

AO32x2_ASAP7_75t_L g1336 ( 
.A1(n_1180),
.A2(n_1190),
.A3(n_1061),
.B1(n_1028),
.B2(n_1043),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1038),
.B(n_1130),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1041),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1049),
.A2(n_1058),
.B(n_1135),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1038),
.B(n_1130),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1056),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1038),
.A2(n_1029),
.B(n_1022),
.C(n_1015),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1038),
.A2(n_1029),
.B1(n_1022),
.B2(n_1153),
.Y(n_1343)
);

INVx3_ASAP7_75t_SL g1344 ( 
.A(n_1082),
.Y(n_1344)
);

INVx1_ASAP7_75t_SL g1345 ( 
.A(n_1154),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1056),
.Y(n_1346)
);

CKINVDCx12_ASAP7_75t_R g1347 ( 
.A(n_1154),
.Y(n_1347)
);

OR2x6_ASAP7_75t_L g1348 ( 
.A(n_1169),
.B(n_1002),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1310),
.A2(n_1222),
.B1(n_1343),
.B2(n_1335),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1252),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1281),
.Y(n_1351)
);

INVx5_ASAP7_75t_L g1352 ( 
.A(n_1332),
.Y(n_1352)
);

BUFx2_ASAP7_75t_R g1353 ( 
.A(n_1213),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1210),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1332),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1335),
.A2(n_1322),
.B1(n_1347),
.B2(n_1196),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1222),
.A2(n_1248),
.B1(n_1322),
.B2(n_1233),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1312),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1202),
.Y(n_1359)
);

INVx4_ASAP7_75t_L g1360 ( 
.A(n_1225),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1205),
.Y(n_1361)
);

INVx8_ASAP7_75t_L g1362 ( 
.A(n_1330),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_1225),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1292),
.B(n_1302),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1281),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1332),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1312),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1332),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1227),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1212),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1238),
.B(n_1264),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1250),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1345),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1273),
.Y(n_1374)
);

NAND2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1292),
.B(n_1287),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1228),
.A2(n_1256),
.B(n_1244),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1237),
.B(n_1241),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1292),
.B(n_1297),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1345),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1206),
.B(n_1204),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1230),
.A2(n_1194),
.B1(n_1333),
.B2(n_1314),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1338),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1234),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1242),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1237),
.Y(n_1385)
);

AOI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1301),
.A2(n_1263),
.B(n_1266),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1241),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1194),
.A2(n_1337),
.B1(n_1333),
.B2(n_1340),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1256),
.A2(n_1244),
.B(n_1220),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1199),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1301),
.A2(n_1249),
.B(n_1223),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1334),
.B(n_1342),
.Y(n_1392)
);

AO21x1_ASAP7_75t_SL g1393 ( 
.A1(n_1221),
.A2(n_1219),
.B(n_1246),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1247),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1311),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1314),
.B(n_1337),
.Y(n_1396)
);

CKINVDCx6p67_ASAP7_75t_R g1397 ( 
.A(n_1309),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1257),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1262),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1319),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1217),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1207),
.A2(n_1216),
.B1(n_1340),
.B2(n_1258),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1225),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1323),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1245),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1308),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1240),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1248),
.A2(n_1233),
.B1(n_1221),
.B2(n_1239),
.Y(n_1408)
);

NAND2x1_ASAP7_75t_L g1409 ( 
.A(n_1289),
.B(n_1294),
.Y(n_1409)
);

BUFx2_ASAP7_75t_SL g1410 ( 
.A(n_1260),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1218),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1325),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1195),
.A2(n_1320),
.B(n_1313),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1258),
.A2(n_1216),
.B1(n_1200),
.B2(n_1286),
.Y(n_1414)
);

INVx4_ASAP7_75t_L g1415 ( 
.A(n_1245),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1245),
.Y(n_1416)
);

BUFx2_ASAP7_75t_R g1417 ( 
.A(n_1344),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1316),
.A2(n_1321),
.B1(n_1328),
.B2(n_1324),
.Y(n_1418)
);

AO21x1_ASAP7_75t_SL g1419 ( 
.A1(n_1219),
.A2(n_1253),
.B(n_1236),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1251),
.A2(n_1198),
.B1(n_1259),
.B2(n_1224),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1224),
.A2(n_1264),
.B1(n_1232),
.B2(n_1215),
.Y(n_1421)
);

AO21x1_ASAP7_75t_L g1422 ( 
.A1(n_1272),
.A2(n_1339),
.B(n_1320),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1254),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1274),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1238),
.B(n_1218),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1331),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1268),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1268),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1289),
.A2(n_1243),
.B1(n_1214),
.B2(n_1229),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1336),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1267),
.A2(n_1203),
.B1(n_1208),
.B2(n_1315),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1291),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1280),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1327),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1291),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1329),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1220),
.A2(n_1211),
.B(n_1339),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1282),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1278),
.Y(n_1439)
);

BUFx2_ASAP7_75t_R g1440 ( 
.A(n_1269),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1278),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1284),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1270),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1271),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1265),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1341),
.B(n_1346),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1271),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1289),
.A2(n_1255),
.B1(n_1261),
.B2(n_1231),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1260),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1275),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1306),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1283),
.B(n_1279),
.Y(n_1452)
);

AOI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1303),
.A2(n_1304),
.B(n_1305),
.Y(n_1453)
);

BUFx2_ASAP7_75t_SL g1454 ( 
.A(n_1260),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1298),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1306),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_SL g1457 ( 
.A1(n_1235),
.A2(n_1288),
.B(n_1285),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1209),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1209),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1304),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1299),
.A2(n_1277),
.B(n_1285),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1226),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1197),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1226),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1307),
.A2(n_1317),
.B1(n_1326),
.B2(n_1348),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1317),
.A2(n_1300),
.B(n_1296),
.Y(n_1466)
);

OR2x6_ASAP7_75t_L g1467 ( 
.A(n_1293),
.B(n_1348),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1307),
.A2(n_1348),
.B1(n_1330),
.B2(n_1294),
.Y(n_1468)
);

NAND2x1_ASAP7_75t_L g1469 ( 
.A(n_1295),
.B(n_1293),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1326),
.A2(n_1330),
.B1(n_1276),
.B2(n_1271),
.Y(n_1470)
);

AO21x2_ASAP7_75t_L g1471 ( 
.A1(n_1296),
.A2(n_1053),
.B(n_1228),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1290),
.B(n_1022),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1201),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1206),
.B(n_1022),
.Y(n_1474)
);

AO21x1_ASAP7_75t_L g1475 ( 
.A1(n_1233),
.A2(n_1053),
.B(n_1272),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1318),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1301),
.A2(n_1263),
.B(n_1249),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1201),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1396),
.B(n_1474),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1369),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1460),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1350),
.B(n_1430),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1377),
.B(n_1369),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1349),
.B(n_1357),
.C(n_1408),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1428),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1455),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1386),
.A2(n_1391),
.B(n_1477),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1377),
.B(n_1385),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1428),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1387),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1355),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1350),
.B(n_1430),
.Y(n_1492)
);

BUFx4f_ASAP7_75t_SL g1493 ( 
.A(n_1450),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1413),
.B(n_1422),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1427),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1409),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1358),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1380),
.B(n_1388),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1351),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1367),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1401),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1381),
.B(n_1423),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1373),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1409),
.A2(n_1469),
.B(n_1453),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1355),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1365),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1365),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1375),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1392),
.A2(n_1419),
.B1(n_1414),
.B2(n_1356),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1352),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1453),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1383),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1457),
.A2(n_1375),
.B(n_1422),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1392),
.A2(n_1472),
.B(n_1402),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1455),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1475),
.A2(n_1471),
.B(n_1466),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1383),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1419),
.A2(n_1475),
.B1(n_1452),
.B2(n_1418),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1420),
.A2(n_1421),
.B(n_1443),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1471),
.B(n_1466),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1384),
.Y(n_1521)
);

AO21x2_ASAP7_75t_L g1522 ( 
.A1(n_1471),
.A2(n_1466),
.B(n_1461),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1451),
.B(n_1467),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1379),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1384),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1394),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1451),
.B(n_1467),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1432),
.A2(n_1435),
.B(n_1456),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1393),
.B(n_1407),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1406),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1452),
.B(n_1424),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1465),
.A2(n_1431),
.B(n_1429),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1394),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1467),
.B(n_1456),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1398),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1390),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1399),
.Y(n_1537)
);

AO21x2_ASAP7_75t_L g1538 ( 
.A1(n_1461),
.A2(n_1412),
.B(n_1361),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1399),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1352),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1364),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1433),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1458),
.B(n_1459),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1359),
.B(n_1370),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1378),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1378),
.Y(n_1546)
);

AOI21xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1445),
.A2(n_1448),
.B(n_1463),
.Y(n_1547)
);

NOR2x1_ASAP7_75t_L g1548 ( 
.A(n_1467),
.B(n_1368),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1426),
.B(n_1464),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1400),
.B(n_1478),
.Y(n_1550)
);

AO21x2_ASAP7_75t_L g1551 ( 
.A1(n_1442),
.A2(n_1439),
.B(n_1441),
.Y(n_1551)
);

AO21x2_ASAP7_75t_L g1552 ( 
.A1(n_1438),
.A2(n_1437),
.B(n_1389),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1434),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1437),
.A2(n_1389),
.B(n_1376),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1366),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1389),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1366),
.Y(n_1557)
);

NAND2x1p5_ASAP7_75t_L g1558 ( 
.A(n_1352),
.B(n_1368),
.Y(n_1558)
);

AOI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1425),
.A2(n_1478),
.B(n_1374),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_SL g1560 ( 
.A(n_1353),
.B(n_1417),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1504),
.B(n_1425),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1486),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1486),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1528),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1482),
.B(n_1382),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1520),
.B(n_1372),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1482),
.B(n_1382),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1504),
.B(n_1508),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1528),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1510),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1492),
.B(n_1473),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1496),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1485),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1556),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1484),
.A2(n_1509),
.B1(n_1498),
.B2(n_1514),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1489),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1520),
.B(n_1476),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1538),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1484),
.A2(n_1532),
.B1(n_1519),
.B2(n_1518),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1483),
.B(n_1488),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1511),
.B(n_1476),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1483),
.B(n_1468),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1552),
.B(n_1411),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1508),
.B(n_1476),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1552),
.B(n_1411),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1516),
.B(n_1436),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1488),
.B(n_1476),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1516),
.B(n_1476),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1516),
.B(n_1436),
.Y(n_1589)
);

CKINVDCx12_ASAP7_75t_R g1590 ( 
.A(n_1493),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1494),
.B(n_1371),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1559),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1494),
.B(n_1371),
.Y(n_1593)
);

NOR2x1_ASAP7_75t_SL g1594 ( 
.A(n_1510),
.B(n_1454),
.Y(n_1594)
);

INVx4_ASAP7_75t_R g1595 ( 
.A(n_1491),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1515),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1515),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1497),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1494),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1499),
.B(n_1404),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1501),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_L g1602 ( 
.A(n_1551),
.B(n_1410),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1494),
.B(n_1371),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1579),
.B(n_1502),
.C(n_1479),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1574),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1598),
.B(n_1500),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1598),
.B(n_1503),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1579),
.A2(n_1547),
.B(n_1513),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_SL g1609 ( 
.A(n_1601),
.B(n_1560),
.Y(n_1609)
);

NAND4xp25_ASAP7_75t_L g1610 ( 
.A(n_1575),
.B(n_1549),
.C(n_1530),
.D(n_1553),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1580),
.B(n_1524),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1580),
.B(n_1495),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1575),
.A2(n_1547),
.B1(n_1536),
.B2(n_1531),
.C(n_1542),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_SL g1614 ( 
.A1(n_1590),
.A2(n_1354),
.B1(n_1445),
.B2(n_1401),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1582),
.A2(n_1440),
.B1(n_1558),
.B2(n_1450),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_R g1616 ( 
.A(n_1562),
.B(n_1354),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1582),
.A2(n_1558),
.B1(n_1548),
.B2(n_1470),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1594),
.A2(n_1494),
.B(n_1592),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1573),
.B(n_1495),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1562),
.A2(n_1529),
.B1(n_1531),
.B2(n_1534),
.Y(n_1620)
);

AOI221xp5_ASAP7_75t_L g1621 ( 
.A1(n_1573),
.A2(n_1543),
.B1(n_1544),
.B2(n_1529),
.C(n_1499),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1576),
.A2(n_1544),
.B1(n_1507),
.B2(n_1506),
.C(n_1550),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1591),
.B(n_1481),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1576),
.B(n_1506),
.Y(n_1624)
);

OA211x2_ASAP7_75t_L g1625 ( 
.A1(n_1600),
.A2(n_1548),
.B(n_1446),
.C(n_1558),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1587),
.B(n_1507),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1587),
.B(n_1512),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1593),
.B(n_1481),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1597),
.B(n_1512),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1597),
.B(n_1517),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1562),
.B(n_1517),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1563),
.B(n_1521),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1563),
.B(n_1521),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1563),
.B(n_1525),
.Y(n_1634)
);

NAND3xp33_ASAP7_75t_L g1635 ( 
.A(n_1588),
.B(n_1602),
.C(n_1581),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1596),
.B(n_1525),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1596),
.B(n_1526),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1596),
.B(n_1526),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_L g1639 ( 
.A(n_1588),
.B(n_1557),
.C(n_1555),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1565),
.B(n_1533),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1577),
.A2(n_1510),
.B1(n_1540),
.B2(n_1462),
.Y(n_1641)
);

NAND2xp33_ASAP7_75t_SL g1642 ( 
.A(n_1570),
.B(n_1540),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1565),
.B(n_1533),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1603),
.A2(n_1534),
.B1(n_1523),
.B2(n_1527),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1565),
.B(n_1535),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1578),
.A2(n_1554),
.B(n_1487),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1577),
.A2(n_1540),
.B1(n_1462),
.B2(n_1505),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1567),
.B(n_1571),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1571),
.B(n_1537),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1561),
.B(n_1523),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1603),
.B(n_1522),
.Y(n_1651)
);

AOI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1586),
.A2(n_1550),
.B1(n_1539),
.B2(n_1480),
.C(n_1490),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1603),
.B(n_1522),
.Y(n_1653)
);

OAI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1588),
.A2(n_1395),
.B1(n_1541),
.B2(n_1546),
.C(n_1545),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1586),
.B(n_1522),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_L g1656 ( 
.A(n_1602),
.B(n_1581),
.C(n_1577),
.Y(n_1656)
);

OA211x2_ASAP7_75t_L g1657 ( 
.A1(n_1600),
.A2(n_1594),
.B(n_1595),
.C(n_1540),
.Y(n_1657)
);

OAI221xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1599),
.A2(n_1397),
.B1(n_1395),
.B2(n_1505),
.C(n_1491),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1584),
.A2(n_1534),
.B1(n_1527),
.B2(n_1523),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1605),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1650),
.B(n_1568),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1605),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1655),
.B(n_1564),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1650),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1642),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1646),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1646),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1612),
.B(n_1652),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1626),
.B(n_1586),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1656),
.B(n_1568),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1629),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1630),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1624),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1635),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1646),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1640),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1651),
.B(n_1561),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1651),
.B(n_1653),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1646),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1611),
.B(n_1569),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1643),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1653),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1631),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1623),
.B(n_1568),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1623),
.B(n_1561),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1645),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1648),
.B(n_1569),
.Y(n_1687)
);

NOR2xp67_ASAP7_75t_L g1688 ( 
.A(n_1618),
.B(n_1639),
.Y(n_1688)
);

NAND2x1p5_ASAP7_75t_L g1689 ( 
.A(n_1628),
.B(n_1570),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1649),
.B(n_1566),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1627),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1632),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1633),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1634),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1644),
.B(n_1583),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_R g1696 ( 
.A(n_1609),
.B(n_1397),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1636),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1668),
.B(n_1606),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1668),
.B(n_1607),
.Y(n_1699)
);

NOR3x1_ASAP7_75t_L g1700 ( 
.A(n_1665),
.B(n_1604),
.C(n_1610),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1680),
.B(n_1619),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1674),
.A2(n_1604),
.B1(n_1613),
.B2(n_1608),
.C(n_1621),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1660),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1680),
.B(n_1637),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1693),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1660),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1662),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1662),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1693),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1677),
.B(n_1568),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1692),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1661),
.B(n_1568),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1692),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1697),
.Y(n_1714)
);

INVx2_ASAP7_75t_SL g1715 ( 
.A(n_1661),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1677),
.B(n_1616),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1673),
.B(n_1622),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1678),
.B(n_1585),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1673),
.B(n_1614),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1697),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1678),
.B(n_1585),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1691),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1661),
.B(n_1572),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1663),
.B(n_1638),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1691),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1683),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1674),
.B(n_1589),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1683),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1690),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1690),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1678),
.B(n_1585),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1671),
.B(n_1589),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1671),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1684),
.B(n_1620),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1672),
.B(n_1589),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1684),
.B(n_1659),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1672),
.B(n_1614),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1722),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1717),
.B(n_1694),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_SL g1740 ( 
.A(n_1737),
.B(n_1658),
.Y(n_1740)
);

OR2x6_ASAP7_75t_L g1741 ( 
.A(n_1716),
.B(n_1665),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1733),
.B(n_1694),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1716),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1701),
.B(n_1687),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1701),
.B(n_1687),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1722),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1736),
.B(n_1734),
.Y(n_1747)
);

NOR2xp67_ASAP7_75t_SL g1748 ( 
.A(n_1705),
.B(n_1540),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1719),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1733),
.B(n_1694),
.Y(n_1750)
);

NAND2x1_ASAP7_75t_L g1751 ( 
.A(n_1723),
.B(n_1664),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1698),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1729),
.B(n_1669),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1709),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1725),
.B(n_1676),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1709),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1725),
.Y(n_1757)
);

OAI21xp5_ASAP7_75t_SL g1758 ( 
.A1(n_1702),
.A2(n_1615),
.B(n_1617),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1714),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1736),
.B(n_1685),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1714),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1699),
.B(n_1676),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1720),
.Y(n_1763)
);

NOR2x1_ASAP7_75t_L g1764 ( 
.A(n_1711),
.B(n_1688),
.Y(n_1764)
);

OR2x6_ASAP7_75t_L g1765 ( 
.A(n_1715),
.B(n_1688),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1720),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1704),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1715),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1703),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1711),
.B(n_1681),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1703),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1713),
.B(n_1681),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1734),
.B(n_1685),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1723),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1713),
.B(n_1686),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1700),
.B(n_1686),
.Y(n_1776)
);

NAND2x1p5_ASAP7_75t_L g1777 ( 
.A(n_1723),
.B(n_1664),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1729),
.B(n_1683),
.Y(n_1778)
);

NAND2x1_ASAP7_75t_SL g1779 ( 
.A(n_1712),
.B(n_1670),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1706),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1739),
.B(n_1727),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1747),
.B(n_1730),
.Y(n_1782)
);

INVx1_ASAP7_75t_SL g1783 ( 
.A(n_1764),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1741),
.B(n_1712),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1741),
.B(n_1712),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1769),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1771),
.Y(n_1787)
);

OA21x2_ASAP7_75t_L g1788 ( 
.A1(n_1758),
.A2(n_1675),
.B(n_1666),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1741),
.B(n_1730),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1760),
.B(n_1710),
.Y(n_1790)
);

INVx3_ASAP7_75t_SL g1791 ( 
.A(n_1765),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1773),
.B(n_1710),
.Y(n_1792)
);

OAI21x1_ASAP7_75t_L g1793 ( 
.A1(n_1779),
.A2(n_1679),
.B(n_1667),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1740),
.A2(n_1625),
.B1(n_1654),
.B2(n_1641),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1739),
.B(n_1704),
.Y(n_1795)
);

INVxp67_ASAP7_75t_L g1796 ( 
.A(n_1754),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1752),
.B(n_1706),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1780),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1767),
.B(n_1724),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1776),
.B(n_1708),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1756),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1738),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1765),
.B(n_1712),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1777),
.B(n_1718),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1777),
.B(n_1718),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1749),
.B(n_1724),
.Y(n_1806)
);

INVx2_ASAP7_75t_SL g1807 ( 
.A(n_1751),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1746),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1765),
.B(n_1721),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1743),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1762),
.B(n_1708),
.Y(n_1811)
);

NOR2x1_ASAP7_75t_L g1812 ( 
.A(n_1757),
.B(n_1726),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1774),
.A2(n_1670),
.B1(n_1664),
.B2(n_1695),
.Y(n_1813)
);

CKINVDCx16_ASAP7_75t_R g1814 ( 
.A(n_1768),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1759),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1778),
.B(n_1721),
.Y(n_1816)
);

OAI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1794),
.A2(n_1744),
.B1(n_1745),
.B2(n_1753),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1783),
.A2(n_1772),
.B(n_1770),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1808),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1808),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1815),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1796),
.B(n_1761),
.Y(n_1822)
);

AOI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1794),
.A2(n_1748),
.B1(n_1670),
.B2(n_1775),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1783),
.A2(n_1670),
.B1(n_1772),
.B2(n_1770),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1815),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1810),
.A2(n_1775),
.B1(n_1766),
.B2(n_1763),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1814),
.B(n_1731),
.Y(n_1827)
);

NAND3xp33_ASAP7_75t_L g1828 ( 
.A(n_1796),
.B(n_1750),
.C(n_1742),
.Y(n_1828)
);

AOI221xp5_ASAP7_75t_L g1829 ( 
.A1(n_1806),
.A2(n_1750),
.B1(n_1742),
.B2(n_1755),
.C(n_1696),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1807),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1807),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1791),
.Y(n_1832)
);

O2A1O1Ixp33_ASAP7_75t_L g1833 ( 
.A1(n_1791),
.A2(n_1800),
.B(n_1801),
.C(n_1810),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1814),
.A2(n_1661),
.B1(n_1682),
.B2(n_1689),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1782),
.A2(n_1625),
.B1(n_1696),
.B2(n_1695),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1801),
.B(n_1782),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1807),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1791),
.A2(n_1755),
.B1(n_1642),
.B2(n_1726),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1800),
.B(n_1731),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1788),
.A2(n_1728),
.B(n_1732),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1788),
.A2(n_1728),
.B(n_1735),
.Y(n_1841)
);

CKINVDCx8_ASAP7_75t_R g1842 ( 
.A(n_1788),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1842),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1832),
.B(n_1833),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1827),
.B(n_1789),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1836),
.B(n_1799),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1819),
.Y(n_1847)
);

INVx1_ASAP7_75t_SL g1848 ( 
.A(n_1836),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1820),
.Y(n_1849)
);

INVx1_ASAP7_75t_SL g1850 ( 
.A(n_1830),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1839),
.B(n_1799),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1823),
.A2(n_1817),
.B1(n_1835),
.B2(n_1829),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1829),
.A2(n_1788),
.B1(n_1784),
.B2(n_1785),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1831),
.Y(n_1854)
);

NOR2x1_ASAP7_75t_L g1855 ( 
.A(n_1837),
.B(n_1812),
.Y(n_1855)
);

OAI21xp33_ASAP7_75t_SL g1856 ( 
.A1(n_1818),
.A2(n_1785),
.B(n_1784),
.Y(n_1856)
);

INVxp67_ASAP7_75t_L g1857 ( 
.A(n_1821),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1825),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1826),
.B(n_1789),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1828),
.A2(n_1788),
.B(n_1797),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1822),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1822),
.B(n_1816),
.Y(n_1862)
);

O2A1O1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1843),
.A2(n_1841),
.B(n_1797),
.C(n_1840),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1850),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1843),
.A2(n_1812),
.B(n_1838),
.Y(n_1865)
);

NOR3xp33_ASAP7_75t_L g1866 ( 
.A(n_1844),
.B(n_1839),
.C(n_1824),
.Y(n_1866)
);

NOR3xp33_ASAP7_75t_L g1867 ( 
.A(n_1852),
.B(n_1834),
.C(n_1785),
.Y(n_1867)
);

OAI322xp33_ASAP7_75t_L g1868 ( 
.A1(n_1860),
.A2(n_1787),
.A3(n_1798),
.B1(n_1786),
.B2(n_1781),
.C1(n_1802),
.C2(n_1795),
.Y(n_1868)
);

AOI221xp5_ASAP7_75t_L g1869 ( 
.A1(n_1859),
.A2(n_1853),
.B1(n_1846),
.B2(n_1848),
.C(n_1857),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1854),
.B(n_1816),
.Y(n_1870)
);

O2A1O1Ixp5_ASAP7_75t_L g1871 ( 
.A1(n_1862),
.A2(n_1784),
.B(n_1803),
.C(n_1802),
.Y(n_1871)
);

A2O1A1Ixp33_ASAP7_75t_L g1872 ( 
.A1(n_1856),
.A2(n_1793),
.B(n_1813),
.C(n_1803),
.Y(n_1872)
);

AOI211xp5_ASAP7_75t_L g1873 ( 
.A1(n_1861),
.A2(n_1803),
.B(n_1809),
.C(n_1795),
.Y(n_1873)
);

AOI221xp5_ASAP7_75t_L g1874 ( 
.A1(n_1857),
.A2(n_1787),
.B1(n_1798),
.B2(n_1786),
.C(n_1802),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1845),
.B(n_1816),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1869),
.B(n_1858),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1870),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1875),
.Y(n_1878)
);

NOR2x1_ASAP7_75t_SL g1879 ( 
.A(n_1864),
.B(n_1847),
.Y(n_1879)
);

NAND4xp75_ASAP7_75t_L g1880 ( 
.A(n_1865),
.B(n_1855),
.C(n_1849),
.D(n_1809),
.Y(n_1880)
);

NOR2x1_ASAP7_75t_L g1881 ( 
.A(n_1868),
.B(n_1851),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1866),
.B(n_1858),
.Y(n_1882)
);

NOR4xp25_ASAP7_75t_L g1883 ( 
.A(n_1863),
.B(n_1781),
.C(n_1811),
.D(n_1804),
.Y(n_1883)
);

NOR4xp25_ASAP7_75t_L g1884 ( 
.A(n_1874),
.B(n_1872),
.C(n_1873),
.D(n_1867),
.Y(n_1884)
);

AND5x1_ASAP7_75t_L g1885 ( 
.A(n_1871),
.B(n_1793),
.C(n_1805),
.D(n_1804),
.E(n_1792),
.Y(n_1885)
);

NAND3xp33_ASAP7_75t_SL g1886 ( 
.A(n_1869),
.B(n_1805),
.C(n_1811),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1864),
.B(n_1790),
.Y(n_1887)
);

NAND2x1p5_ASAP7_75t_L g1888 ( 
.A(n_1885),
.B(n_1360),
.Y(n_1888)
);

NOR2x1_ASAP7_75t_L g1889 ( 
.A(n_1880),
.B(n_1405),
.Y(n_1889)
);

NAND4xp25_ASAP7_75t_L g1890 ( 
.A(n_1887),
.B(n_1881),
.C(n_1876),
.D(n_1882),
.Y(n_1890)
);

XNOR2xp5_ASAP7_75t_L g1891 ( 
.A(n_1884),
.B(n_1790),
.Y(n_1891)
);

NAND4xp25_ASAP7_75t_SL g1892 ( 
.A(n_1876),
.B(n_1792),
.C(n_1793),
.D(n_1663),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1879),
.B(n_1707),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1893),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1889),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1890),
.A2(n_1886),
.B1(n_1878),
.B2(n_1877),
.Y(n_1896)
);

NOR3xp33_ASAP7_75t_L g1897 ( 
.A(n_1892),
.B(n_1883),
.C(n_1363),
.Y(n_1897)
);

AOI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1891),
.A2(n_1682),
.B1(n_1657),
.B2(n_1683),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1888),
.Y(n_1899)
);

CKINVDCx20_ASAP7_75t_R g1900 ( 
.A(n_1891),
.Y(n_1900)
);

NOR3xp33_ASAP7_75t_L g1901 ( 
.A(n_1894),
.B(n_1896),
.C(n_1899),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1895),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1900),
.Y(n_1903)
);

XNOR2x1_ASAP7_75t_L g1904 ( 
.A(n_1898),
.B(n_1405),
.Y(n_1904)
);

NOR3xp33_ASAP7_75t_SL g1905 ( 
.A(n_1897),
.B(n_1647),
.C(n_1669),
.Y(n_1905)
);

XNOR2xp5_ASAP7_75t_L g1906 ( 
.A(n_1900),
.B(n_1416),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1903),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1902),
.Y(n_1908)
);

NAND4xp25_ASAP7_75t_L g1909 ( 
.A(n_1901),
.B(n_1416),
.C(n_1363),
.D(n_1403),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1907),
.Y(n_1910)
);

NOR3xp33_ASAP7_75t_L g1911 ( 
.A(n_1910),
.B(n_1908),
.C(n_1909),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1911),
.A2(n_1906),
.B1(n_1904),
.B2(n_1905),
.Y(n_1912)
);

AOI22xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1911),
.A2(n_1360),
.B1(n_1363),
.B2(n_1403),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_SL g1914 ( 
.A1(n_1912),
.A2(n_1360),
.B1(n_1415),
.B2(n_1403),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1913),
.Y(n_1915)
);

AOI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1707),
.B1(n_1415),
.B2(n_1683),
.C(n_1679),
.Y(n_1916)
);

OA21x2_ASAP7_75t_L g1917 ( 
.A1(n_1914),
.A2(n_1675),
.B(n_1666),
.Y(n_1917)
);

OAI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1916),
.A2(n_1415),
.B(n_1444),
.Y(n_1918)
);

OAI221xp5_ASAP7_75t_R g1919 ( 
.A1(n_1918),
.A2(n_1917),
.B1(n_1362),
.B2(n_1657),
.C(n_1679),
.Y(n_1919)
);

AOI221xp5_ASAP7_75t_L g1920 ( 
.A1(n_1919),
.A2(n_1683),
.B1(n_1682),
.B2(n_1667),
.C(n_1679),
.Y(n_1920)
);

AOI211xp5_ASAP7_75t_L g1921 ( 
.A1(n_1920),
.A2(n_1449),
.B(n_1540),
.C(n_1447),
.Y(n_1921)
);


endmodule