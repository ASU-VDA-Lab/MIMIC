module fake_jpeg_7798_n_285 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_285);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_28),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_27),
.B1(n_31),
.B2(n_16),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_25),
.B1(n_33),
.B2(n_19),
.Y(n_77)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_48),
.Y(n_87)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_31),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_27),
.B1(n_16),
.B2(n_30),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_21),
.B1(n_33),
.B2(n_19),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_27),
.B1(n_16),
.B2(n_33),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_61),
.B1(n_28),
.B2(n_24),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_23),
.B1(n_32),
.B2(n_18),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_29),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_20),
.C(n_17),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_63),
.B(n_78),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_64),
.A2(n_8),
.B1(n_14),
.B2(n_3),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_32),
.B1(n_18),
.B2(n_26),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_65),
.A2(n_85),
.B1(n_22),
.B2(n_21),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_70),
.B1(n_74),
.B2(n_77),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_20),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_79),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_10),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_54),
.B1(n_59),
.B2(n_55),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_48),
.B1(n_20),
.B2(n_17),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_59),
.B1(n_55),
.B2(n_47),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_48),
.B(n_21),
.C(n_20),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_86),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_29),
.B1(n_22),
.B2(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_47),
.B(n_10),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_22),
.B1(n_29),
.B2(n_21),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_49),
.B(n_10),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_8),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_93),
.B(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_90),
.B(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_98),
.B(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_115),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_100),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_63),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_118),
.B1(n_72),
.B2(n_90),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_108),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_0),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_0),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_0),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_20),
.B1(n_8),
.B2(n_2),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_63),
.B1(n_83),
.B2(n_67),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_11),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_119),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_120),
.A2(n_124),
.B1(n_133),
.B2(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_123),
.B(n_12),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_80),
.B1(n_67),
.B2(n_81),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_62),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_136),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_69),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_139),
.B(n_145),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_80),
.B1(n_67),
.B2(n_69),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_73),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_82),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_143),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_95),
.B(n_66),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_146),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_94),
.A2(n_72),
.B(n_84),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_107),
.B(n_92),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_153),
.Y(n_192)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_97),
.B(n_106),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_159),
.A2(n_167),
.B(n_169),
.Y(n_179)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_161),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_133),
.B1(n_124),
.B2(n_128),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_98),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_92),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_113),
.B1(n_103),
.B2(n_118),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_125),
.B1(n_119),
.B2(n_143),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_101),
.B(n_105),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_172),
.B(n_176),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_116),
.B(n_101),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_173),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_112),
.C(n_100),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_1),
.C(n_5),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_121),
.A2(n_112),
.B(n_76),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_0),
.B(n_1),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_120),
.C(n_135),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_196),
.C(n_201),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_121),
.B(n_130),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_197),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_183),
.B(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_135),
.C(n_125),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_129),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_156),
.B1(n_154),
.B2(n_153),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_12),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_177),
.C(n_159),
.Y(n_212)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_204),
.B(n_207),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_162),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_208),
.C(n_211),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_192),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_175),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_180),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_218),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_213),
.B(n_217),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_164),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_202),
.C(n_191),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_178),
.B(n_172),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

OAI21x1_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_171),
.B(n_168),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_185),
.B(n_167),
.Y(n_222)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_223),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_233),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_210),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_195),
.B1(n_194),
.B2(n_193),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_228),
.A2(n_229),
.B1(n_236),
.B2(n_219),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_188),
.B1(n_186),
.B2(n_181),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_203),
.A2(n_188),
.B1(n_186),
.B2(n_189),
.Y(n_231)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_215),
.A2(n_182),
.B1(n_174),
.B2(n_149),
.Y(n_234)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_160),
.B1(n_187),
.B2(n_170),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_208),
.C(n_209),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_248),
.Y(n_254)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_151),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_245),
.Y(n_257)
);

AOI221xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_231),
.B1(n_226),
.B2(n_239),
.C(n_228),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_211),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_250),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_150),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_209),
.C(n_214),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_251),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_206),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_229),
.B(n_219),
.CI(n_212),
.CON(n_252),
.SN(n_252)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_252),
.B(n_233),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_244),
.A2(n_237),
.B(n_230),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_261),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_262),
.B(n_161),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_257),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_232),
.B(n_151),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_201),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_241),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_250),
.B1(n_241),
.B2(n_173),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_267),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_266),
.B(n_270),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_249),
.C(n_240),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_253),
.A3(n_263),
.B1(n_262),
.B2(n_259),
.C1(n_161),
.C2(n_129),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_155),
.C(n_129),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_1),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_155),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_271),
.A2(n_6),
.B(n_7),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_276),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_274),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_275),
.A2(n_264),
.B1(n_269),
.B2(n_267),
.Y(n_278)
);

AOI321xp33_ASAP7_75t_SL g280 ( 
.A1(n_278),
.A2(n_264),
.A3(n_272),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_281),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_SL g281 ( 
.A(n_279),
.B(n_7),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_282),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_277),
.B(n_9),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_7),
.B1(n_9),
.B2(n_13),
.Y(n_285)
);


endmodule