module fake_jpeg_1061_n_160 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_61),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_0),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_72),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_55),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_47),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_53),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_56),
.B1(n_55),
.B2(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_81),
.B1(n_42),
.B2(n_43),
.Y(n_100)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_59),
.B1(n_41),
.B2(n_49),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_83),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_77),
.B(n_50),
.Y(n_101)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_46),
.B(n_19),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_44),
.B1(n_42),
.B2(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_65),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_87),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_41),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_63),
.B1(n_40),
.B2(n_48),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_100),
.B1(n_90),
.B2(n_93),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_97),
.Y(n_107)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_15),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_81),
.B1(n_45),
.B2(n_4),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_101),
.B(n_102),
.Y(n_111)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_104),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_111),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_80),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_120),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_121),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_2),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_119),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_3),
.B(n_5),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_21),
.C(n_38),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_6),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_7),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_130),
.Y(n_139)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_17),
.A3(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_133),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_8),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_120),
.C(n_13),
.Y(n_143)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_137),
.A2(n_118),
.B1(n_113),
.B2(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_132),
.B(n_136),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_144),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_12),
.C(n_28),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_SL g146 ( 
.A(n_139),
.B(n_125),
.C(n_142),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_149),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_128),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_148),
.A2(n_136),
.B1(n_132),
.B2(n_134),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_151),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_138),
.B1(n_137),
.B2(n_131),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_145),
.Y(n_155)
);

AOI21x1_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_152),
.B(n_129),
.Y(n_156)
);

AOI321xp33_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_147),
.A3(n_22),
.B1(n_24),
.B2(n_39),
.C(n_25),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_157),
.A2(n_8),
.B(n_9),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_10),
.B(n_11),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_11),
.Y(n_160)
);


endmodule