module fake_jpeg_30257_n_152 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_152);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_40),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_17),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_16),
.B1(n_23),
.B2(n_17),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_23),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_28),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_59),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_56),
.B1(n_61),
.B2(n_0),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_15),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_63),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_53),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_21),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_13),
.B1(n_23),
.B2(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_31),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_5),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_51),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_19),
.B1(n_18),
.B2(n_27),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_27),
.B(n_21),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_70),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_74),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_53),
.B(n_43),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_64),
.B1(n_45),
.B2(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_89),
.B1(n_85),
.B2(n_84),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_43),
.B1(n_49),
.B2(n_45),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_49),
.B(n_59),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_67),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_69),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_50),
.A3(n_64),
.B1(n_5),
.B2(n_6),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_75),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_50),
.C(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_104),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_116),
.B(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_77),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_84),
.B1(n_85),
.B2(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_85),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_80),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_97),
.C(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_115),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_88),
.A2(n_66),
.B1(n_64),
.B2(n_7),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_97),
.B1(n_88),
.B2(n_102),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_118),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_94),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_92),
.C(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_105),
.B1(n_110),
.B2(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

AOI21x1_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_130),
.B(n_133),
.Y(n_136)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_116),
.B1(n_114),
.B2(n_111),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_132),
.A2(n_125),
.B1(n_118),
.B2(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_131),
.C(n_127),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_120),
.C(n_126),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_139),
.B(n_140),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_136),
.A2(n_100),
.B(n_131),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_142),
.B(n_144),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_139),
.B(n_108),
.CI(n_101),
.CON(n_144),
.SN(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_143),
.A2(n_140),
.B(n_138),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.Y(n_148)
);

AOI211xp5_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_135),
.B(n_137),
.C(n_142),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_101),
.C(n_93),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_148),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_93),
.Y(n_152)
);


endmodule