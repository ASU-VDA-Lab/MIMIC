module fake_jpeg_12439_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_2),
.Y(n_6)
);

INVx13_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_0),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_10),
.A2(n_9),
.B1(n_11),
.B2(n_8),
.Y(n_13)
);

OAI21xp33_ASAP7_75t_SL g20 ( 
.A1(n_13),
.A2(n_7),
.B(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_18),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_16),
.A2(n_17),
.B1(n_19),
.B2(n_11),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_3),
.C(n_7),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_22),
.B1(n_14),
.B2(n_19),
.Y(n_24)
);

AO22x1_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_26),
.B1(n_21),
.B2(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_16),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_30),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_30),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_32),
.B(n_27),
.Y(n_33)
);


endmodule