module fake_jpeg_29501_n_70 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_70);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_70;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx24_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_10),
.B(n_2),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_17),
.C(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_9),
.B(n_5),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_25),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_16),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_24),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_20),
.B1(n_25),
.B2(n_23),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR3xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_24),
.C(n_19),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_27),
.B(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_44),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_25),
.A3(n_38),
.B1(n_40),
.B2(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_19),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_50),
.B1(n_19),
.B2(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_53),
.B(n_42),
.Y(n_54)
);

AND2x6_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_13),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_8),
.B(n_5),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_41),
.B1(n_17),
.B2(n_18),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_55),
.A2(n_58),
.B1(n_21),
.B2(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_13),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_21),
.C(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_62),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_61),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_13),
.C(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_58),
.B1(n_57),
.B2(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_67),
.Y(n_68)
);

OAI21x1_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_6),
.B(n_7),
.Y(n_67)
);

AOI322xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_63),
.A3(n_7),
.B1(n_16),
.B2(n_4),
.C1(n_3),
.C2(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_16),
.Y(n_70)
);


endmodule