module fake_jpeg_815_n_343 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_46),
.Y(n_118)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_47),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_53),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_55),
.Y(n_151)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_20),
.B(n_0),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_57),
.B(n_2),
.C(n_3),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_59),
.B(n_61),
.Y(n_112)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_33),
.B(n_6),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_5),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_62),
.B(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_31),
.B(n_8),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_67),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_8),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_17),
.B(n_9),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_11),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_82),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_80),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

CKINVDCx9p33_ASAP7_75t_R g131 ( 
.A(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_19),
.B(n_11),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_87),
.Y(n_128)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g154 ( 
.A(n_85),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_29),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_15),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_91),
.Y(n_130)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_25),
.B(n_1),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_1),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_28),
.B(n_1),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_41),
.B(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_98),
.Y(n_145)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_100),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_27),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_41),
.B(n_2),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_2),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_100),
.B(n_95),
.Y(n_108)
);

AND2x4_ASAP7_75t_L g191 ( 
.A(n_108),
.B(n_129),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_62),
.A2(n_37),
.B1(n_39),
.B2(n_43),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_78),
.B1(n_83),
.B2(n_55),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_66),
.A2(n_39),
.B1(n_27),
.B2(n_42),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_120),
.A2(n_133),
.B1(n_53),
.B2(n_48),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_67),
.A2(n_42),
.B1(n_34),
.B2(n_43),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_138),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_73),
.A2(n_21),
.B1(n_34),
.B2(n_29),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_129),
.A2(n_107),
.B1(n_151),
.B2(n_132),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_87),
.A2(n_21),
.B1(n_29),
.B2(n_45),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_139),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_69),
.B(n_2),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_3),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_142),
.B(n_147),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_52),
.A2(n_29),
.B(n_45),
.C(n_4),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_4),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_159),
.B1(n_192),
.B2(n_119),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_154),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_157),
.B(n_167),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_166),
.B1(n_172),
.B2(n_179),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_58),
.B1(n_64),
.B2(n_80),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_81),
.B1(n_88),
.B2(n_45),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_4),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_164),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_45),
.B1(n_145),
.B2(n_137),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_108),
.B(n_122),
.C(n_105),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_171),
.A2(n_191),
.B(n_141),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_124),
.B1(n_107),
.B2(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_110),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_181),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_114),
.B(n_106),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_186),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_111),
.A2(n_103),
.B1(n_125),
.B2(n_117),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_180),
.A2(n_184),
.B1(n_140),
.B2(n_148),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_188),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_112),
.A2(n_109),
.B1(n_134),
.B2(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_146),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_115),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_190),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_105),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_118),
.A2(n_102),
.B1(n_113),
.B2(n_119),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_191),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_SL g195 ( 
.A(n_178),
.B(n_123),
.C(n_140),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_206),
.B(n_210),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_118),
.C(n_126),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_165),
.C(n_169),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_176),
.A2(n_113),
.B1(n_102),
.B2(n_153),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_201),
.A2(n_215),
.B1(n_219),
.B2(n_165),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_123),
.B(n_104),
.C(n_126),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_153),
.B1(n_104),
.B2(n_141),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_203),
.B(n_164),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_221),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_164),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_191),
.B(n_172),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_234),
.B(n_193),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_212),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_237),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_185),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_210),
.B(n_185),
.Y(n_226)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

O2A1O1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_206),
.A2(n_180),
.B(n_187),
.C(n_186),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_223),
.B(n_229),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_214),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_236),
.C(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_238),
.B1(n_201),
.B2(n_219),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_190),
.B(n_155),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_200),
.A2(n_155),
.B1(n_170),
.B2(n_173),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_177),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_211),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_200),
.A2(n_155),
.B1(n_168),
.B2(n_183),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_240),
.A2(n_193),
.B1(n_216),
.B2(n_211),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_242),
.B1(n_251),
.B2(n_234),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_230),
.C(n_236),
.Y(n_261)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_195),
.B1(n_197),
.B2(n_216),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_256),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_202),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_254),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_225),
.B(n_199),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_205),
.B(n_209),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_228),
.Y(n_275)
);

CKINVDCx12_ASAP7_75t_R g259 ( 
.A(n_239),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_259),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_265),
.C(n_268),
.Y(n_285)
);

A2O1A1O1Ixp25_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_221),
.B(n_226),
.C(n_228),
.D(n_227),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_262),
.A2(n_252),
.B(n_253),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_263),
.A2(n_264),
.B1(n_241),
.B2(n_251),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_238),
.B1(n_233),
.B2(n_240),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_230),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_220),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_231),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_273),
.C(n_259),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_256),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_276),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_253),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_222),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_254),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_252),
.B(n_246),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_250),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_287),
.B1(n_257),
.B2(n_267),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_272),
.Y(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_289),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_245),
.B(n_243),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_250),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_266),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_284),
.B(n_286),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_267),
.A2(n_258),
.B1(n_251),
.B2(n_257),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_244),
.Y(n_288)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_295),
.B1(n_303),
.B2(n_282),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_273),
.B1(n_242),
.B2(n_262),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_278),
.A2(n_243),
.B1(n_245),
.B2(n_244),
.Y(n_296)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_265),
.C(n_261),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_301),
.C(n_293),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_287),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_268),
.C(n_237),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_235),
.B1(n_249),
.B2(n_208),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_305),
.Y(n_316)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_281),
.C(n_289),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_209),
.C(n_208),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_309),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_286),
.C(n_291),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_313),
.C(n_298),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_300),
.Y(n_311)
);

OAI22x1_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_312),
.B1(n_303),
.B2(n_290),
.Y(n_315)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_288),
.C(n_280),
.Y(n_313)
);

OAI321xp33_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_299),
.A3(n_300),
.B1(n_295),
.B2(n_292),
.C(n_294),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_314),
.A2(n_315),
.B1(n_208),
.B2(n_174),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_175),
.C(n_212),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_306),
.A2(n_279),
.B(n_249),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_321),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_304),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_205),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_313),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_198),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_310),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_325),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_309),
.C(n_212),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_328),
.A2(n_198),
.B(n_161),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_163),
.B1(n_198),
.B2(n_189),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_332),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_331),
.B(n_181),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_329),
.B(n_322),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_337),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_325),
.C(n_181),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_331),
.C(n_330),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_336),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_339),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_181),
.B(n_148),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_104),
.Y(n_343)
);


endmodule