module real_aes_204_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_287;
wire n_503;
wire n_357;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g295 ( .A(n_0), .B(n_212), .Y(n_295) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_1), .A2(n_58), .B1(n_90), .B2(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g177 ( .A(n_2), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_3), .B(n_197), .Y(n_196) );
NAND2xp33_ASAP7_75t_SL g280 ( .A(n_4), .B(n_203), .Y(n_280) );
AOI22xp33_ASAP7_75t_SL g111 ( .A1(n_5), .A2(n_26), .B1(n_112), .B2(n_117), .Y(n_111) );
INVx1_ASAP7_75t_L g271 ( .A(n_6), .Y(n_271) );
AOI222xp33_ASAP7_75t_L g83 ( .A1(n_7), .A2(n_16), .B1(n_65), .B2(n_84), .C1(n_102), .C2(n_106), .Y(n_83) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_8), .A2(n_21), .B1(n_90), .B2(n_98), .Y(n_97) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_9), .A2(n_80), .B1(n_81), .B2(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_9), .Y(n_503) );
AND2x2_ASAP7_75t_L g191 ( .A(n_10), .B(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g193 ( .A(n_11), .Y(n_193) );
AOI221x1_ASAP7_75t_L g274 ( .A1(n_12), .A2(n_205), .B1(n_275), .B2(n_277), .C(n_279), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_13), .B(n_197), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_14), .A2(n_160), .B1(n_161), .B2(n_164), .Y(n_159) );
INVx1_ASAP7_75t_L g164 ( .A(n_14), .Y(n_164) );
AOI22xp33_ASAP7_75t_SL g123 ( .A1(n_15), .A2(n_34), .B1(n_124), .B2(n_128), .Y(n_123) );
AOI221xp5_ASAP7_75t_SL g285 ( .A1(n_17), .A2(n_35), .B1(n_197), .B2(n_205), .C(n_286), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_18), .A2(n_75), .B1(n_140), .B2(n_142), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_19), .A2(n_205), .B(n_210), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_20), .B(n_212), .Y(n_211) );
OAI221xp5_ASAP7_75t_L g169 ( .A1(n_21), .A2(n_58), .B1(n_60), .B2(n_170), .C(n_172), .Y(n_169) );
OR2x2_ASAP7_75t_L g194 ( .A(n_22), .B(n_69), .Y(n_194) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_22), .A2(n_69), .B(n_193), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_23), .B(n_214), .Y(n_265) );
INVxp67_ASAP7_75t_L g273 ( .A(n_24), .Y(n_273) );
AND2x2_ASAP7_75t_L g236 ( .A(n_25), .B(n_226), .Y(n_236) );
INVx3_ASAP7_75t_L g90 ( .A(n_27), .Y(n_90) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_28), .A2(n_57), .B1(n_132), .B2(n_136), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_29), .A2(n_205), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_30), .B(n_214), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_31), .A2(n_80), .B1(n_81), .B2(n_156), .Y(n_79) );
INVx1_ASAP7_75t_L g156 ( .A(n_31), .Y(n_156) );
INVx1_ASAP7_75t_SL g91 ( .A(n_32), .Y(n_91) );
INVx1_ASAP7_75t_L g179 ( .A(n_33), .Y(n_179) );
AND2x2_ASAP7_75t_L g203 ( .A(n_33), .B(n_177), .Y(n_203) );
AND2x2_ASAP7_75t_L g206 ( .A(n_33), .B(n_207), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_36), .A2(n_63), .B1(n_205), .B2(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_37), .B(n_212), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_38), .A2(n_48), .B1(n_152), .B2(n_154), .Y(n_151) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_39), .A2(n_60), .B1(n_90), .B2(n_94), .Y(n_93) );
OAI22xp5_ASAP7_75t_SL g157 ( .A1(n_40), .A2(n_158), .B1(n_159), .B2(n_165), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_40), .Y(n_165) );
AND2x2_ASAP7_75t_L g298 ( .A(n_41), .B(n_226), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_42), .B(n_226), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_43), .A2(n_53), .B1(n_146), .B2(n_149), .Y(n_145) );
INVx1_ASAP7_75t_L g200 ( .A(n_44), .Y(n_200) );
INVx1_ASAP7_75t_L g209 ( .A(n_44), .Y(n_209) );
OAI22xp5_ASAP7_75t_SL g161 ( .A1(n_45), .A2(n_55), .B1(n_162), .B2(n_163), .Y(n_161) );
INVx1_ASAP7_75t_L g163 ( .A(n_45), .Y(n_163) );
INVx1_ASAP7_75t_L g92 ( .A(n_46), .Y(n_92) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_47), .B(n_197), .Y(n_235) );
AND2x2_ASAP7_75t_L g227 ( .A(n_49), .B(n_226), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_50), .B(n_214), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_51), .B(n_212), .Y(n_223) );
AND2x2_ASAP7_75t_SL g266 ( .A(n_52), .B(n_192), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_54), .A2(n_205), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g162 ( .A(n_55), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_55), .B(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_SL g256 ( .A(n_56), .B(n_243), .Y(n_256) );
INVxp33_ASAP7_75t_L g174 ( .A(n_58), .Y(n_174) );
INVx1_ASAP7_75t_L g202 ( .A(n_59), .Y(n_202) );
INVx1_ASAP7_75t_L g207 ( .A(n_59), .Y(n_207) );
INVxp67_ASAP7_75t_L g173 ( .A(n_60), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_61), .B(n_197), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_62), .A2(n_64), .B1(n_197), .B2(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_66), .B(n_212), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_67), .B(n_212), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_68), .A2(n_205), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_70), .B(n_214), .Y(n_222) );
INVxp67_ASAP7_75t_L g276 ( .A(n_71), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_72), .B(n_197), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_73), .B(n_214), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_73), .A2(n_80), .B1(n_81), .B2(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_73), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_74), .A2(n_205), .B(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_SL g171 ( .A(n_76), .Y(n_171) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_166), .B1(n_180), .B2(n_492), .C(n_493), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_157), .Y(n_78) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_81), .Y(n_80) );
OR2x2_ASAP7_75t_L g81 ( .A(n_82), .B(n_130), .Y(n_81) );
NAND3xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_111), .C(n_123), .Y(n_82) );
INVx3_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx6_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
AND2x4_ASAP7_75t_L g104 ( .A(n_87), .B(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g113 ( .A(n_87), .B(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
INVx2_ASAP7_75t_L g110 ( .A(n_88), .Y(n_110) );
AND2x2_ASAP7_75t_L g121 ( .A(n_88), .B(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_88), .Y(n_127) );
OAI22x1_ASAP7_75t_L g88 ( .A1(n_89), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g94 ( .A(n_90), .Y(n_94) );
INVx2_ASAP7_75t_L g98 ( .A(n_90), .Y(n_98) );
INVx1_ASAP7_75t_L g101 ( .A(n_90), .Y(n_101) );
AND2x2_ASAP7_75t_L g109 ( .A(n_93), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g122 ( .A(n_93), .Y(n_122) );
BUFx2_ASAP7_75t_L g150 ( .A(n_93), .Y(n_150) );
AND2x4_ASAP7_75t_L g134 ( .A(n_95), .B(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g141 ( .A(n_95), .B(n_109), .Y(n_141) );
AND2x4_ASAP7_75t_L g153 ( .A(n_95), .B(n_121), .Y(n_153) );
AND2x4_ASAP7_75t_L g95 ( .A(n_96), .B(n_99), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x4_ASAP7_75t_L g108 ( .A(n_97), .B(n_99), .Y(n_108) );
INVx1_ASAP7_75t_L g116 ( .A(n_97), .Y(n_116) );
AND2x2_ASAP7_75t_L g126 ( .A(n_97), .B(n_100), .Y(n_126) );
INVxp67_ASAP7_75t_L g105 ( .A(n_99), .Y(n_105) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g120 ( .A(n_100), .B(n_116), .Y(n_120) );
INVx2_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx6_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g129 ( .A(n_108), .B(n_121), .Y(n_129) );
AND2x4_ASAP7_75t_L g138 ( .A(n_108), .B(n_135), .Y(n_138) );
AND2x2_ASAP7_75t_L g148 ( .A(n_109), .B(n_120), .Y(n_148) );
AND2x4_ASAP7_75t_L g135 ( .A(n_110), .B(n_122), .Y(n_135) );
BUFx6f_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x4_ASAP7_75t_L g144 ( .A(n_120), .B(n_135), .Y(n_144) );
BUFx12f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x4_ASAP7_75t_L g149 ( .A(n_126), .B(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g155 ( .A(n_126), .B(n_135), .Y(n_155) );
BUFx5_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NAND4xp25_ASAP7_75t_L g130 ( .A(n_131), .B(n_139), .C(n_145), .D(n_151), .Y(n_130) );
INVx2_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
INVx8_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx8_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_159), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
AND3x1_ASAP7_75t_SL g168 ( .A(n_169), .B(n_175), .C(n_178), .Y(n_168) );
INVxp67_ASAP7_75t_L g501 ( .A(n_169), .Y(n_501) );
CKINVDCx8_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_175), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_175), .A2(n_509), .B(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g248 ( .A(n_176), .B(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_SL g506 ( .A(n_176), .B(n_178), .Y(n_506) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g208 ( .A(n_177), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_178), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2x1p5_ASAP7_75t_L g253 ( .A(n_179), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_414), .Y(n_183) );
NOR3xp33_ASAP7_75t_SL g184 ( .A(n_185), .B(n_338), .C(n_388), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_318), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_257), .B(n_299), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_237), .Y(n_188) );
INVx1_ASAP7_75t_SL g424 ( .A(n_189), .Y(n_424) );
AOI32xp33_ASAP7_75t_L g455 ( .A1(n_189), .A2(n_437), .A3(n_456), .B1(n_457), .B2(n_458), .Y(n_455) );
AND2x2_ASAP7_75t_L g457 ( .A(n_189), .B(n_314), .Y(n_457) );
AND2x4_ASAP7_75t_SL g189 ( .A(n_190), .B(n_217), .Y(n_189) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_190), .Y(n_238) );
INVx5_ASAP7_75t_L g317 ( .A(n_190), .Y(n_317) );
OR2x2_ASAP7_75t_L g324 ( .A(n_190), .B(n_316), .Y(n_324) );
INVx2_ASAP7_75t_L g329 ( .A(n_190), .Y(n_329) );
AND2x2_ASAP7_75t_L g341 ( .A(n_190), .B(n_218), .Y(n_341) );
AND2x2_ASAP7_75t_L g346 ( .A(n_190), .B(n_228), .Y(n_346) );
OR2x2_ASAP7_75t_L g353 ( .A(n_190), .B(n_240), .Y(n_353) );
AND2x4_ASAP7_75t_L g362 ( .A(n_190), .B(n_229), .Y(n_362) );
O2A1O1Ixp33_ASAP7_75t_SL g404 ( .A1(n_190), .A2(n_320), .B(n_355), .C(n_393), .Y(n_404) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_195), .Y(n_190) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_192), .Y(n_226) );
AND2x2_ASAP7_75t_SL g192 ( .A(n_193), .B(n_194), .Y(n_192) );
AND2x4_ASAP7_75t_L g216 ( .A(n_193), .B(n_194), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_204), .B(n_216), .Y(n_195) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_203), .Y(n_197) );
INVx1_ASAP7_75t_L g281 ( .A(n_198), .Y(n_281) );
AND2x4_ASAP7_75t_L g198 ( .A(n_199), .B(n_201), .Y(n_198) );
AND2x6_ASAP7_75t_L g212 ( .A(n_199), .B(n_207), .Y(n_212) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_L g214 ( .A(n_201), .B(n_209), .Y(n_214) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx5_ASAP7_75t_L g215 ( .A(n_203), .Y(n_215) );
AND2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_208), .Y(n_205) );
BUFx3_ASAP7_75t_L g250 ( .A(n_206), .Y(n_250) );
INVx2_ASAP7_75t_L g255 ( .A(n_207), .Y(n_255) );
AND2x4_ASAP7_75t_L g252 ( .A(n_208), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g249 ( .A(n_209), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_213), .B(n_215), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_215), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_215), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_215), .A2(n_264), .B(n_265), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_215), .A2(n_287), .B(n_288), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_215), .A2(n_295), .B(n_296), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_216), .B(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_216), .B(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_216), .B(n_276), .Y(n_275) );
NOR3xp33_ASAP7_75t_L g279 ( .A(n_216), .B(n_280), .C(n_281), .Y(n_279) );
INVx3_ASAP7_75t_SL g354 ( .A(n_217), .Y(n_354) );
AND2x2_ASAP7_75t_L g400 ( .A(n_217), .B(n_317), .Y(n_400) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_228), .Y(n_217) );
AND2x2_ASAP7_75t_L g239 ( .A(n_218), .B(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g331 ( .A(n_218), .B(n_229), .Y(n_331) );
AND2x2_ASAP7_75t_L g335 ( .A(n_218), .B(n_314), .Y(n_335) );
INVx1_ASAP7_75t_L g361 ( .A(n_218), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_218), .B(n_229), .Y(n_383) );
INVx2_ASAP7_75t_L g387 ( .A(n_218), .Y(n_387) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_218), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_218), .B(n_317), .Y(n_464) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_225), .B(n_227), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_225), .A2(n_230), .B(n_236), .Y(n_229) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_225), .A2(n_230), .B(n_236), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_226), .Y(n_225) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_226), .A2(n_285), .B(n_289), .Y(n_284) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g398 ( .A(n_229), .B(n_240), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_235), .Y(n_230) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx1_ASAP7_75t_L g408 ( .A(n_238), .Y(n_408) );
NAND2xp33_ASAP7_75t_SL g433 ( .A(n_238), .B(n_325), .Y(n_433) );
AND2x2_ASAP7_75t_L g475 ( .A(n_239), .B(n_317), .Y(n_475) );
AND2x2_ASAP7_75t_L g386 ( .A(n_240), .B(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g449 ( .A(n_240), .Y(n_449) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_241), .Y(n_314) );
AOI21x1_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_245), .B(n_256), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_243), .A2(n_261), .B(n_262), .Y(n_260) );
BUFx4f_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx3_ASAP7_75t_L g278 ( .A(n_244), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_251), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_247), .A2(n_252), .B1(n_270), .B2(n_272), .Y(n_269) );
AND2x4_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
INVx1_ASAP7_75t_L g510 ( .A(n_248), .Y(n_510) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_252), .Y(n_492) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_253), .Y(n_509) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_257), .A2(n_340), .B1(n_442), .B2(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_282), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_258), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_258), .B(n_365), .Y(n_364) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_267), .Y(n_258) );
INVx2_ASAP7_75t_L g305 ( .A(n_259), .Y(n_305) );
OR2x2_ASAP7_75t_L g309 ( .A(n_259), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_259), .B(n_322), .Y(n_327) );
AND2x4_ASAP7_75t_SL g337 ( .A(n_259), .B(n_268), .Y(n_337) );
OR2x2_ASAP7_75t_L g344 ( .A(n_259), .B(n_284), .Y(n_344) );
OR2x2_ASAP7_75t_L g356 ( .A(n_259), .B(n_268), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_259), .B(n_284), .Y(n_370) );
INVx1_ASAP7_75t_L g375 ( .A(n_259), .Y(n_375) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_259), .Y(n_393) );
AND2x2_ASAP7_75t_L g456 ( .A(n_259), .B(n_376), .Y(n_456) );
INVx2_ASAP7_75t_L g460 ( .A(n_259), .Y(n_460) );
OR2x2_ASAP7_75t_L g467 ( .A(n_259), .B(n_357), .Y(n_467) );
OR2x2_ASAP7_75t_L g489 ( .A(n_259), .B(n_490), .Y(n_489) );
OR2x6_ASAP7_75t_L g259 ( .A(n_260), .B(n_266), .Y(n_259) );
AND2x2_ASAP7_75t_L g306 ( .A(n_267), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_267), .B(n_290), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_267), .B(n_366), .Y(n_428) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g325 ( .A(n_268), .Y(n_325) );
AND2x4_ASAP7_75t_L g376 ( .A(n_268), .B(n_377), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_268), .B(n_321), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_268), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_268), .B(n_310), .Y(n_469) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_274), .Y(n_268) );
INVx4_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI21x1_ASAP7_75t_L g291 ( .A1(n_278), .A2(n_292), .B(n_298), .Y(n_291) );
AND2x2_ASAP7_75t_L g336 ( .A(n_282), .B(n_337), .Y(n_336) );
AO221x1_ASAP7_75t_L g410 ( .A1(n_282), .A2(n_325), .B1(n_356), .B2(n_411), .C(n_412), .Y(n_410) );
OAI322xp33_ASAP7_75t_L g462 ( .A1(n_282), .A2(n_382), .A3(n_463), .B1(n_465), .B2(n_466), .C1(n_467), .C2(n_468), .Y(n_462) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_290), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx3_ASAP7_75t_L g304 ( .A(n_284), .Y(n_304) );
INVx2_ASAP7_75t_L g310 ( .A(n_284), .Y(n_310) );
AND2x2_ASAP7_75t_L g322 ( .A(n_284), .B(n_290), .Y(n_322) );
INVx1_ASAP7_75t_L g367 ( .A(n_284), .Y(n_367) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_284), .Y(n_423) );
INVx1_ASAP7_75t_L g307 ( .A(n_290), .Y(n_307) );
OR2x2_ASAP7_75t_L g357 ( .A(n_290), .B(n_310), .Y(n_357) );
INVx2_ASAP7_75t_L g377 ( .A(n_290), .Y(n_377) );
INVx1_ASAP7_75t_L g430 ( .A(n_290), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_290), .B(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI21xp33_ASAP7_75t_SL g300 ( .A1(n_301), .A2(n_308), .B(n_311), .Y(n_300) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_301), .A2(n_340), .B1(n_342), .B2(n_346), .C(n_347), .Y(n_339) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
NOR2x1p5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g426 ( .A(n_305), .Y(n_426) );
INVx1_ASAP7_75t_SL g345 ( .A(n_306), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_306), .A2(n_451), .B(n_453), .Y(n_450) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_307), .Y(n_350) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_310), .Y(n_413) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
OAI211xp5_ASAP7_75t_L g388 ( .A1(n_313), .A2(n_389), .B(n_394), .C(n_405), .Y(n_388) );
OR2x2_ASAP7_75t_L g478 ( .A(n_313), .B(n_383), .Y(n_478) );
AND2x2_ASAP7_75t_L g480 ( .A(n_313), .B(n_346), .Y(n_480) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g320 ( .A(n_314), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g382 ( .A(n_314), .B(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g420 ( .A(n_314), .B(n_387), .Y(n_420) );
OA33x2_ASAP7_75t_L g427 ( .A1(n_314), .A2(n_344), .A3(n_428), .B1(n_429), .B2(n_431), .B3(n_433), .Y(n_427) );
OR2x2_ASAP7_75t_L g438 ( .A(n_314), .B(n_423), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_314), .B(n_362), .Y(n_452) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g340 ( .A(n_316), .B(n_341), .Y(n_340) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_316), .A2(n_346), .B1(n_390), .B2(n_391), .Y(n_389) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_317), .B(n_397), .C(n_430), .Y(n_429) );
AOI322xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_323), .A3(n_325), .B1(n_326), .B2(n_328), .C1(n_332), .C2(n_336), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g425 ( .A(n_321), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
A2O1A1Ixp33_ASAP7_75t_L g380 ( .A1(n_322), .A2(n_337), .B(n_381), .C(n_384), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_323), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
NAND4xp25_ASAP7_75t_SL g444 ( .A(n_324), .B(n_353), .C(n_445), .D(n_447), .Y(n_444) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx2_ASAP7_75t_L g334 ( .A(n_329), .Y(n_334) );
OR2x2_ASAP7_75t_L g379 ( .A(n_329), .B(n_331), .Y(n_379) );
AND2x2_ASAP7_75t_L g448 ( .A(n_330), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g453 ( .A(n_334), .B(n_448), .Y(n_453) );
BUFx2_ASAP7_75t_L g446 ( .A(n_335), .Y(n_446) );
INVx1_ASAP7_75t_SL g476 ( .A(n_336), .Y(n_476) );
AND2x4_ASAP7_75t_L g412 ( .A(n_337), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g465 ( .A(n_337), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_358), .C(n_380), .Y(n_338) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_SL g402 ( .A(n_344), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g470 ( .A1(n_344), .A2(n_471), .B(n_472), .C(n_481), .Y(n_470) );
OR2x2_ASAP7_75t_L g392 ( .A(n_345), .B(n_393), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_351), .B1(n_354), .B2(n_355), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_349), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_352), .B(n_409), .Y(n_491) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g466 ( .A(n_353), .B(n_354), .Y(n_466) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g411 ( .A(n_357), .Y(n_411) );
AOI222xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_363), .B1(n_368), .B2(n_372), .C1(n_373), .C2(n_378), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_361), .Y(n_372) );
AND2x2_ASAP7_75t_L g419 ( .A(n_362), .B(n_420), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_362), .A2(n_435), .B1(n_440), .B2(n_444), .Y(n_434) );
INVx2_ASAP7_75t_SL g487 ( .A(n_362), .Y(n_487) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g443 ( .A(n_367), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_367), .B(n_430), .Y(n_490) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_373), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g441 ( .A(n_375), .Y(n_441) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_376), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g484 ( .A(n_376), .B(n_413), .Y(n_484) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g409 ( .A(n_383), .Y(n_409) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g488 ( .A(n_386), .Y(n_488) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_387), .Y(n_432) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_399), .B(n_401), .C(n_404), .Y(n_394) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_396), .B(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g439 ( .A(n_401), .Y(n_439) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_410), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_408), .B(n_409), .Y(n_407) );
NOR3xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_454), .C(n_470), .Y(n_414) );
NAND3xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_434), .C(n_450), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .B1(n_424), .B2(n_425), .C(n_427), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_436), .B(n_439), .Y(n_435) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g463 ( .A(n_449), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g471 ( .A(n_453), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_461), .Y(n_454) );
INVx2_ASAP7_75t_L g477 ( .A(n_456), .Y(n_477) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g468 ( .A(n_459), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_476), .B1(n_477), .B2(n_478), .C(n_479), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_485), .B1(n_489), .B2(n_491), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
OAI222xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_496), .B2(n_502), .C1(n_504), .C2(n_507), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
endmodule