module fake_netlist_5_1595_n_1271 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1271);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1271;

wire n_924;
wire n_1263;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_292;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_307;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_600;
wire n_223;
wire n_264;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_254;
wire n_1233;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1121;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_582;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_261;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_222;
wire n_1123;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_302;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_212;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_205;
wire n_1136;
wire n_754;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_202;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_605;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_522;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1012;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_277;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_312;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_246;
wire n_1042;
wire n_269;
wire n_285;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_533;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_92),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_143),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_108),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_87),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_49),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_5),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_5),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_3),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_88),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_6),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_29),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_86),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_17),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_27),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_131),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_141),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_17),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_76),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_45),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_9),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_49),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_0),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_28),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_0),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_61),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_38),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_38),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_45),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_165),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_21),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_44),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_122),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_148),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_53),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_58),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_115),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_12),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_35),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_170),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_28),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_149),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_25),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_26),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_145),
.Y(n_237)
);

BUFx8_ASAP7_75t_SL g238 ( 
.A(n_93),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_114),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_117),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_31),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_79),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_50),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_24),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_54),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_164),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_22),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_21),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_171),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_101),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_57),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_124),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_140),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_7),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_97),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_129),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_14),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_74),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_89),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_90),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_146),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_173),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_135),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_50),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_144),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_91),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_40),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_8),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_159),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_160),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_24),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_70),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_1),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_147),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_152),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_161),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_51),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_163),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_100),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_44),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_6),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_156),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_119),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_172),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_151),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_52),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_176),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_3),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_111),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_162),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_37),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_104),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_12),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_11),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_42),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_138),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_121),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_82),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_236),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_238),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_216),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_178),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_236),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_197),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_216),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_236),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_179),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_204),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_252),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_244),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_236),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_236),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_205),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_217),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_206),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_210),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_236),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_242),
.B(n_1),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_235),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_235),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_241),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_2),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_241),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_252),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_197),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_270),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_241),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_188),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_218),
.B(n_2),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_221),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_188),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_193),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_225),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_218),
.B(n_4),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_241),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_241),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_226),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_193),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_189),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_203),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_209),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_270),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_213),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_227),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_219),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_220),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_233),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_231),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_232),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_237),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_194),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_254),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_267),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_277),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_239),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_291),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_250),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_234),
.B(n_4),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_251),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_194),
.Y(n_362)
);

INVxp33_ASAP7_75t_SL g363 ( 
.A(n_198),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_200),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_197),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_200),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_243),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_212),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_243),
.B(n_7),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_214),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_198),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_201),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_294),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_295),
.Y(n_375)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_201),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_278),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_234),
.B(n_8),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_273),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_278),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_273),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_280),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_180),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_181),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_280),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_281),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_184),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_256),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_186),
.Y(n_389)
);

CKINVDCx8_ASAP7_75t_R g390 ( 
.A(n_300),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_337),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_313),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_364),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_330),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_330),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_182),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_283),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

AND3x1_ASAP7_75t_L g401 ( 
.A(n_320),
.B(n_271),
.C(n_268),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_310),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_364),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_325),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_364),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_224),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_338),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_182),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_389),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_364),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_367),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_299),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_283),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_303),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_326),
.B(n_268),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_307),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_328),
.B(n_271),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_366),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_324),
.B(n_253),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_344),
.B(n_183),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_366),
.Y(n_425)
);

BUFx8_ASAP7_75t_L g426 ( 
.A(n_334),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_366),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_312),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_316),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_319),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_366),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_342),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_343),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_360),
.B(n_183),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_345),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_333),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_348),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_349),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_333),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_355),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_356),
.Y(n_444)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_336),
.A2(n_190),
.B(n_187),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_358),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_310),
.B(n_199),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_372),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_375),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_321),
.Y(n_450)
);

OA21x2_ASAP7_75t_L g451 ( 
.A1(n_369),
.A2(n_192),
.B(n_191),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_322),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_374),
.B(n_199),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_302),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_331),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_379),
.B(n_195),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_308),
.B(n_196),
.Y(n_457)
);

AND2x6_ASAP7_75t_L g458 ( 
.A(n_309),
.B(n_200),
.Y(n_458)
);

BUFx12f_ASAP7_75t_L g459 ( 
.A(n_388),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_393),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_415),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_402),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_393),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_393),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_415),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_408),
.B(n_314),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_408),
.B(n_315),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_418),
.B(n_304),
.Y(n_468)
);

BUFx10_ASAP7_75t_L g469 ( 
.A(n_458),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_447),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_392),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_403),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_403),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_403),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_L g475 ( 
.A(n_401),
.B(n_207),
.C(n_202),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_454),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_417),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_391),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_419),
.Y(n_480)
);

CKINVDCx6p67_ASAP7_75t_R g481 ( 
.A(n_459),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_395),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_419),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_402),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_402),
.B(n_332),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_422),
.B(n_335),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_401),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_422),
.A2(n_386),
.B1(n_385),
.B2(n_382),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_392),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_200),
.Y(n_491)
);

OAI22xp33_ASAP7_75t_L g492 ( 
.A1(n_435),
.A2(n_248),
.B1(n_264),
.B2(n_222),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_435),
.B(n_339),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_428),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_458),
.B(n_346),
.Y(n_495)
);

OR2x6_ASAP7_75t_L g496 ( 
.A(n_459),
.B(n_208),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_399),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_428),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_458),
.B(n_350),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_457),
.B(n_200),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_429),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_424),
.B(n_351),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_458),
.B(n_352),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_429),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_L g505 ( 
.A(n_418),
.B(n_215),
.C(n_211),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_424),
.B(n_357),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_430),
.Y(n_507)
);

NAND2xp33_ASAP7_75t_L g508 ( 
.A(n_458),
.B(n_359),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_418),
.B(n_317),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_399),
.Y(n_510)
);

AOI22x1_ASAP7_75t_L g511 ( 
.A1(n_456),
.A2(n_318),
.B1(n_368),
.B2(n_370),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_420),
.B(n_317),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_420),
.B(n_318),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_430),
.Y(n_514)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_392),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_453),
.B(n_361),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

INVxp33_ASAP7_75t_SL g518 ( 
.A(n_395),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_458),
.B(n_368),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_392),
.Y(n_520)
);

CKINVDCx6p67_ASAP7_75t_R g521 ( 
.A(n_454),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_400),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_392),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_458),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_447),
.B(n_353),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_437),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_458),
.B(n_370),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_457),
.B(n_353),
.Y(n_528)
);

NOR3xp33_ASAP7_75t_L g529 ( 
.A(n_437),
.B(n_327),
.C(n_305),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_453),
.B(n_365),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_461),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_466),
.B(n_493),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_478),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_468),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_478),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_461),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_470),
.B(n_454),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_470),
.B(n_458),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_502),
.B(n_458),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_520),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_478),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_462),
.B(n_456),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_484),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_465),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_484),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_525),
.A2(n_456),
.B1(n_454),
.B2(n_420),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_487),
.A2(n_411),
.B1(n_410),
.B2(n_397),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_484),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_462),
.B(n_455),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_469),
.B(n_445),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_469),
.B(n_445),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_510),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_518),
.A2(n_306),
.B1(n_301),
.B2(n_340),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_462),
.B(n_455),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_481),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_485),
.B(n_450),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_485),
.B(n_450),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_485),
.B(n_450),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_481),
.B(n_390),
.Y(n_560)
);

NOR2xp67_ASAP7_75t_L g561 ( 
.A(n_530),
.B(n_528),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_467),
.B(n_530),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_468),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_477),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_469),
.B(n_445),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_506),
.B(n_363),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_477),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_501),
.B(n_450),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_479),
.B(n_480),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_469),
.B(n_240),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_479),
.B(n_450),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_480),
.Y(n_572)
);

AO221x1_ASAP7_75t_L g573 ( 
.A1(n_492),
.A2(n_488),
.B1(n_240),
.B2(n_475),
.C(n_498),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_520),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_L g575 ( 
.A1(n_475),
.A2(n_410),
.B1(n_397),
.B2(n_373),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_483),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_483),
.B(n_442),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_510),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_488),
.A2(n_451),
.B1(n_376),
.B2(n_363),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_494),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_L g581 ( 
.A(n_491),
.B(n_240),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_494),
.B(n_442),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_509),
.A2(n_411),
.B1(n_416),
.B2(n_398),
.Y(n_583)
);

INVx8_ASAP7_75t_L g584 ( 
.A(n_491),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_524),
.B(n_240),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_524),
.B(n_240),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_498),
.B(n_442),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_504),
.B(n_442),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_510),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_504),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_507),
.A2(n_451),
.B1(n_376),
.B2(n_442),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_507),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_516),
.B(n_340),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_514),
.B(n_491),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_514),
.B(n_411),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_522),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_491),
.B(n_411),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_522),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_486),
.B(n_362),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_497),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_497),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_491),
.B(n_411),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_509),
.A2(n_416),
.B1(n_398),
.B2(n_373),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_524),
.B(n_436),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_512),
.B(n_436),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_491),
.B(n_398),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_512),
.B(n_436),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_513),
.B(n_436),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_513),
.B(n_436),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_491),
.B(n_416),
.Y(n_610)
);

HB1xp67_ASAP7_75t_SL g611 ( 
.A(n_529),
.Y(n_611)
);

NOR2xp67_ASAP7_75t_SL g612 ( 
.A(n_505),
.B(n_390),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_500),
.B(n_436),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_472),
.Y(n_614)
);

NOR3xp33_ASAP7_75t_L g615 ( 
.A(n_482),
.B(n_441),
.C(n_396),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_500),
.B(n_436),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_519),
.B(n_436),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_460),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_500),
.B(n_444),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_527),
.B(n_495),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_500),
.B(n_444),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_521),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_520),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_499),
.B(n_444),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_500),
.A2(n_362),
.B1(n_371),
.B2(n_381),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_526),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_472),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_500),
.B(n_444),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_473),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_551),
.A2(n_508),
.B(n_503),
.Y(n_630)
);

AO21x1_ASAP7_75t_L g631 ( 
.A1(n_532),
.A2(n_245),
.B(n_228),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_626),
.B(n_396),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_561),
.B(n_489),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_551),
.A2(n_520),
.B(n_523),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_542),
.B(n_500),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_562),
.B(n_489),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_546),
.B(n_511),
.Y(n_637)
);

A2O1A1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_547),
.A2(n_505),
.B(n_266),
.C(n_269),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_534),
.B(n_521),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_552),
.A2(n_520),
.B(n_523),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_552),
.A2(n_520),
.B(n_523),
.Y(n_641)
);

OAI21xp33_ASAP7_75t_L g642 ( 
.A1(n_566),
.A2(n_511),
.B(n_288),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_579),
.A2(n_569),
.B1(n_591),
.B2(n_583),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_565),
.A2(n_523),
.B(n_515),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_563),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_531),
.B(n_471),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_536),
.B(n_544),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_599),
.B(n_371),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_556),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_600),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_565),
.A2(n_523),
.B(n_515),
.Y(n_651)
);

INVx11_ASAP7_75t_L g652 ( 
.A(n_560),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_623),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_600),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_622),
.Y(n_655)
);

O2A1O1Ixp5_ASAP7_75t_L g656 ( 
.A1(n_620),
.A2(n_471),
.B(n_517),
.C(n_490),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_537),
.Y(n_657)
);

OAI21xp33_ASAP7_75t_L g658 ( 
.A1(n_593),
.A2(n_603),
.B(n_625),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_620),
.A2(n_523),
.B(n_515),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_574),
.A2(n_515),
.B(n_490),
.Y(n_660)
);

AOI21x1_ASAP7_75t_L g661 ( 
.A1(n_538),
.A2(n_474),
.B(n_473),
.Y(n_661)
);

A2O1A1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_595),
.A2(n_260),
.B(n_246),
.C(n_249),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_533),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_549),
.B(n_471),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_574),
.A2(n_515),
.B(n_490),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_540),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_573),
.A2(n_607),
.B1(n_608),
.B2(n_605),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_623),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_622),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_601),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_564),
.A2(n_476),
.B1(n_496),
.B2(n_311),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_537),
.B(n_381),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_567),
.B(n_572),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_574),
.A2(n_515),
.B(n_490),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_574),
.A2(n_517),
.B(n_471),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_596),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_576),
.B(n_580),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_540),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_539),
.A2(n_463),
.B(n_460),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_575),
.B(n_426),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_612),
.B(n_382),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_550),
.A2(n_476),
.B1(n_496),
.B2(n_185),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_624),
.A2(n_517),
.B(n_474),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_590),
.A2(n_592),
.B1(n_555),
.B2(n_605),
.Y(n_684)
);

A2O1A1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_607),
.A2(n_276),
.B(n_255),
.C(n_279),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_623),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_608),
.A2(n_476),
.B1(n_496),
.B2(n_386),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_609),
.B(n_517),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_617),
.A2(n_463),
.B(n_460),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_617),
.A2(n_464),
.B(n_463),
.Y(n_690)
);

OAI21xp33_ASAP7_75t_L g691 ( 
.A1(n_609),
.A2(n_288),
.B(n_281),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_598),
.A2(n_582),
.B(n_587),
.C(n_577),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_623),
.Y(n_693)
);

NOR2xp67_ASAP7_75t_L g694 ( 
.A(n_614),
.B(n_627),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_624),
.A2(n_464),
.B(n_394),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_557),
.A2(n_464),
.B(n_394),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_568),
.B(n_444),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_554),
.B(n_385),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_533),
.Y(n_699)
);

O2A1O1Ixp5_ASAP7_75t_L g700 ( 
.A1(n_570),
.A2(n_289),
.B(n_452),
.C(n_440),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_535),
.B(n_444),
.Y(n_701)
);

OAI21xp33_ASAP7_75t_SL g702 ( 
.A1(n_570),
.A2(n_476),
.B(n_496),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_615),
.B(n_396),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_SL g704 ( 
.A(n_584),
.B(n_476),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_558),
.A2(n_394),
.B(n_392),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_559),
.A2(n_394),
.B(n_392),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_588),
.A2(n_292),
.B(n_261),
.C(n_432),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_540),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_604),
.A2(n_425),
.B(n_394),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_535),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_541),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_604),
.A2(n_425),
.B(n_394),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_611),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_571),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_585),
.B(n_441),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_584),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_584),
.A2(n_425),
.B(n_394),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_585),
.B(n_441),
.Y(n_718)
);

BUFx12f_ASAP7_75t_L g719 ( 
.A(n_584),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_606),
.A2(n_610),
.B1(n_597),
.B2(n_602),
.Y(n_720)
);

NAND3xp33_ASAP7_75t_L g721 ( 
.A(n_594),
.B(n_426),
.C(n_390),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_613),
.A2(n_425),
.B(n_394),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_616),
.A2(n_431),
.B(n_425),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_541),
.A2(n_443),
.B(n_438),
.C(n_432),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_619),
.A2(n_431),
.B(n_425),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_621),
.A2(n_431),
.B(n_425),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_586),
.B(n_301),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_543),
.B(n_545),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_543),
.B(n_496),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_714),
.B(n_426),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_636),
.B(n_306),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_630),
.A2(n_581),
.B(n_628),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_697),
.A2(n_581),
.B(n_586),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_649),
.Y(n_734)
);

O2A1O1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_637),
.A2(n_545),
.B(n_589),
.C(n_578),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_648),
.B(n_311),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_657),
.B(n_548),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_632),
.B(n_548),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_669),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_672),
.B(n_426),
.Y(n_740)
);

NOR2x1_ASAP7_75t_SL g741 ( 
.A(n_716),
.B(n_553),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_663),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_634),
.A2(n_578),
.B(n_553),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_650),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_647),
.B(n_589),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_716),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_640),
.A2(n_618),
.B(n_629),
.Y(n_747)
);

O2A1O1Ixp5_ASAP7_75t_L g748 ( 
.A1(n_631),
.A2(n_618),
.B(n_407),
.C(n_405),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_654),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_641),
.A2(n_431),
.B(n_425),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_699),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_658),
.B(n_426),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_668),
.Y(n_753)
);

BUFx2_ASAP7_75t_L g754 ( 
.A(n_645),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_673),
.B(n_452),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_667),
.A2(n_451),
.B1(n_265),
.B2(n_297),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_633),
.B(n_223),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_727),
.B(n_715),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_720),
.A2(n_451),
.B1(n_272),
.B2(n_297),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_635),
.A2(n_431),
.B(n_451),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_716),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_SL g762 ( 
.A1(n_638),
.A2(n_407),
.B(n_409),
.C(n_405),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_642),
.A2(n_718),
.B(n_643),
.C(n_702),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_644),
.A2(n_431),
.B(n_406),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_643),
.A2(n_434),
.B(n_433),
.C(n_448),
.Y(n_765)
);

NOR2x1_ASAP7_75t_L g766 ( 
.A(n_721),
.B(n_433),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_668),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_651),
.A2(n_431),
.B(n_406),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_713),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_681),
.B(n_229),
.Y(n_770)
);

INVx4_ASAP7_75t_L g771 ( 
.A(n_668),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_688),
.A2(n_431),
.B(n_406),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_680),
.A2(n_434),
.B(n_448),
.C(n_446),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_710),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_686),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_684),
.A2(n_406),
.B(n_404),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_686),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_655),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_711),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_707),
.A2(n_409),
.B(n_400),
.C(n_452),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_684),
.A2(n_679),
.B(n_659),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_724),
.A2(n_438),
.B(n_446),
.C(n_439),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_679),
.A2(n_413),
.B(n_404),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_677),
.B(n_230),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_687),
.A2(n_439),
.B(n_443),
.C(n_265),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_670),
.B(n_449),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_639),
.B(n_272),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_671),
.B(n_274),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_703),
.B(n_440),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_729),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_686),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_692),
.A2(n_421),
.B(n_413),
.Y(n_792)
);

CKINVDCx6p67_ASAP7_75t_R g793 ( 
.A(n_719),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_676),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_694),
.A2(n_290),
.B1(n_296),
.B2(n_285),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_646),
.A2(n_290),
.B1(n_296),
.B2(n_285),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_671),
.B(n_274),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_664),
.A2(n_284),
.B1(n_282),
.B2(n_275),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_693),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_728),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_751),
.Y(n_801)
);

OA21x2_ASAP7_75t_L g802 ( 
.A1(n_781),
.A2(n_656),
.B(n_689),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_778),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_758),
.A2(n_691),
.B(n_698),
.C(n_682),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_752),
.A2(n_662),
.B(n_685),
.C(n_704),
.Y(n_805)
);

AO32x2_ASAP7_75t_L g806 ( 
.A1(n_756),
.A2(n_759),
.A3(n_798),
.B1(n_796),
.B2(n_763),
.Y(n_806)
);

OA21x2_ASAP7_75t_L g807 ( 
.A1(n_748),
.A2(n_690),
.B(n_689),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_784),
.B(n_666),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_733),
.A2(n_683),
.B(n_700),
.Y(n_809)
);

OAI21x1_ASAP7_75t_L g810 ( 
.A1(n_792),
.A2(n_661),
.B(n_695),
.Y(n_810)
);

NOR2xp67_ASAP7_75t_L g811 ( 
.A(n_746),
.B(n_666),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_732),
.A2(n_704),
.B(n_653),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_767),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_752),
.A2(n_696),
.B(n_705),
.C(n_706),
.Y(n_814)
);

AO31x2_ASAP7_75t_L g815 ( 
.A1(n_765),
.A2(n_701),
.A3(n_712),
.B(n_709),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_745),
.A2(n_653),
.B(n_717),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_757),
.A2(n_726),
.B(n_725),
.C(n_723),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_774),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_794),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_738),
.B(n_678),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_744),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_743),
.A2(n_693),
.B(n_690),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_739),
.B(n_708),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_734),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_789),
.B(n_731),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_736),
.A2(n_440),
.B(n_449),
.C(n_412),
.Y(n_826)
);

O2A1O1Ixp5_ASAP7_75t_SL g827 ( 
.A1(n_740),
.A2(n_678),
.B(n_414),
.C(n_412),
.Y(n_827)
);

AO21x1_ASAP7_75t_L g828 ( 
.A1(n_770),
.A2(n_722),
.B(n_675),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_785),
.A2(n_784),
.B(n_780),
.C(n_773),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_SL g830 ( 
.A1(n_800),
.A2(n_674),
.B(n_665),
.C(n_660),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_754),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_749),
.Y(n_832)
);

AO22x2_ASAP7_75t_L g833 ( 
.A1(n_788),
.A2(n_797),
.B1(n_730),
.B2(n_790),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_779),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_769),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_737),
.B(n_755),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_787),
.B(n_708),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_742),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_748),
.A2(n_421),
.B(n_404),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_780),
.A2(n_708),
.B(n_652),
.C(n_693),
.Y(n_840)
);

OAI21x1_ASAP7_75t_L g841 ( 
.A1(n_747),
.A2(n_427),
.B(n_423),
.Y(n_841)
);

AO31x2_ASAP7_75t_L g842 ( 
.A1(n_776),
.A2(n_449),
.A3(n_421),
.B(n_427),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_SL g843 ( 
.A1(n_786),
.A2(n_414),
.B(n_427),
.C(n_423),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_782),
.A2(n_284),
.B(n_275),
.C(n_282),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_753),
.B(n_258),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_753),
.B(n_259),
.Y(n_846)
);

NOR4xp25_ASAP7_75t_L g847 ( 
.A(n_782),
.B(n_253),
.C(n_10),
.D(n_11),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_746),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_793),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_760),
.A2(n_423),
.B(n_413),
.Y(n_850)
);

AOI221x1_ASAP7_75t_L g851 ( 
.A1(n_783),
.A2(n_444),
.B1(n_253),
.B2(n_257),
.C(n_247),
.Y(n_851)
);

NAND2x1_ASAP7_75t_L g852 ( 
.A(n_761),
.B(n_444),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_791),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_795),
.B(n_262),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_766),
.A2(n_298),
.B1(n_263),
.B2(n_13),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_735),
.A2(n_741),
.B(n_750),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_791),
.Y(n_857)
);

AO31x2_ASAP7_75t_L g858 ( 
.A1(n_764),
.A2(n_9),
.A3(n_10),
.B(n_13),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_735),
.A2(n_78),
.B(n_169),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_768),
.A2(n_77),
.B(n_168),
.Y(n_860)
);

AO31x2_ASAP7_75t_L g861 ( 
.A1(n_772),
.A2(n_762),
.A3(n_777),
.B(n_775),
.Y(n_861)
);

AO31x2_ASAP7_75t_L g862 ( 
.A1(n_771),
.A2(n_14),
.A3(n_15),
.B(n_16),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_761),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_801),
.Y(n_864)
);

BUFx4f_ASAP7_75t_SL g865 ( 
.A(n_831),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_804),
.A2(n_777),
.B1(n_775),
.B2(n_771),
.Y(n_866)
);

OAI22xp33_ASAP7_75t_SL g867 ( 
.A1(n_855),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_813),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_818),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_SL g870 ( 
.A1(n_833),
.A2(n_799),
.B1(n_767),
.B2(n_22),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_825),
.B(n_808),
.Y(n_871)
);

BUFx8_ASAP7_75t_L g872 ( 
.A(n_849),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_823),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_821),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_832),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_813),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_833),
.A2(n_799),
.B1(n_767),
.B2(n_23),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_824),
.Y(n_878)
);

AOI21xp33_ASAP7_75t_L g879 ( 
.A1(n_829),
.A2(n_799),
.B(n_767),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_803),
.A2(n_799),
.B1(n_20),
.B2(n_23),
.Y(n_880)
);

CKINVDCx8_ASAP7_75t_R g881 ( 
.A(n_823),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_834),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_819),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_842),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_820),
.B(n_19),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_813),
.Y(n_886)
);

CKINVDCx11_ASAP7_75t_R g887 ( 
.A(n_838),
.Y(n_887)
);

CKINVDCx12_ASAP7_75t_R g888 ( 
.A(n_835),
.Y(n_888)
);

NAND2x1p5_ASAP7_75t_L g889 ( 
.A(n_848),
.B(n_55),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_SL g890 ( 
.A1(n_854),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_890)
);

CKINVDCx11_ASAP7_75t_R g891 ( 
.A(n_853),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_857),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_848),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_836),
.B(n_29),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_842),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_837),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_SL g897 ( 
.A1(n_855),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_863),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_845),
.Y(n_899)
);

BUFx10_ASAP7_75t_L g900 ( 
.A(n_847),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_863),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_SL g902 ( 
.A1(n_846),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_902)
);

INVx6_ASAP7_75t_L g903 ( 
.A(n_811),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_842),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_802),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_847),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_852),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_858),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_828),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_858),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_858),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_860),
.A2(n_802),
.B1(n_807),
.B2(n_806),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_840),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_805),
.A2(n_844),
.B1(n_811),
.B2(n_812),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_817),
.A2(n_856),
.B1(n_816),
.B2(n_814),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_839),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_809),
.Y(n_917)
);

NAND2x1p5_ASAP7_75t_L g918 ( 
.A(n_859),
.B(n_56),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_SL g919 ( 
.A1(n_851),
.A2(n_39),
.B(n_41),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_815),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_822),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_807),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_861),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_862),
.Y(n_924)
);

INVx6_ASAP7_75t_L g925 ( 
.A(n_861),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_862),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_925),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_908),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_920),
.B(n_862),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_920),
.B(n_806),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_884),
.B(n_810),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_910),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_898),
.B(n_826),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_911),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_925),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_884),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_905),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_925),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_904),
.B(n_815),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_923),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_923),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_924),
.B(n_815),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_904),
.Y(n_943)
);

AO21x1_ASAP7_75t_SL g944 ( 
.A1(n_909),
.A2(n_806),
.B(n_827),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_926),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_895),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_895),
.B(n_861),
.Y(n_947)
);

CKINVDCx16_ASAP7_75t_R g948 ( 
.A(n_917),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_869),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_869),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_912),
.B(n_850),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_912),
.B(n_864),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_918),
.Y(n_953)
);

OA21x2_ASAP7_75t_L g954 ( 
.A1(n_915),
.A2(n_906),
.B(n_909),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_874),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_898),
.A2(n_841),
.B1(n_47),
.B2(n_48),
.Y(n_956)
);

OA21x2_ASAP7_75t_L g957 ( 
.A1(n_906),
.A2(n_843),
.B(n_830),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_875),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_882),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_900),
.Y(n_960)
);

CKINVDCx6p67_ASAP7_75t_R g961 ( 
.A(n_913),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_900),
.B(n_46),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_892),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_918),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_914),
.A2(n_110),
.B(n_166),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_927),
.B(n_896),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_949),
.Y(n_967)
);

AO32x2_ASAP7_75t_L g968 ( 
.A1(n_964),
.A2(n_921),
.A3(n_880),
.B1(n_866),
.B2(n_877),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_952),
.B(n_929),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_952),
.B(n_871),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_959),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_964),
.B(n_919),
.Y(n_972)
);

CKINVDCx11_ASAP7_75t_R g973 ( 
.A(n_948),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_942),
.B(n_960),
.Y(n_974)
);

AOI221xp5_ASAP7_75t_L g975 ( 
.A1(n_933),
.A2(n_867),
.B1(n_901),
.B2(n_897),
.C(n_890),
.Y(n_975)
);

AO32x2_ASAP7_75t_L g976 ( 
.A1(n_964),
.A2(n_952),
.A3(n_959),
.B1(n_929),
.B2(n_945),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_955),
.Y(n_977)
);

BUFx10_ASAP7_75t_L g978 ( 
.A(n_933),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_948),
.B(n_899),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_948),
.B(n_894),
.Y(n_980)
);

NAND2xp33_ASAP7_75t_R g981 ( 
.A(n_954),
.B(n_885),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_952),
.B(n_870),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_955),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_955),
.Y(n_984)
);

OA21x2_ASAP7_75t_L g985 ( 
.A1(n_965),
.A2(n_922),
.B(n_879),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_927),
.B(n_873),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_952),
.B(n_883),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_942),
.B(n_893),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_965),
.A2(n_901),
.B(n_902),
.Y(n_989)
);

NOR2x1_ASAP7_75t_SL g990 ( 
.A(n_964),
.B(n_960),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_961),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_961),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_942),
.B(n_873),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_964),
.B(n_889),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_927),
.B(n_868),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_952),
.B(n_929),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_927),
.B(n_868),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_952),
.B(n_916),
.Y(n_998)
);

BUFx12f_ASAP7_75t_L g999 ( 
.A(n_962),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_958),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_961),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_929),
.B(n_930),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_958),
.Y(n_1003)
);

AO21x1_ASAP7_75t_L g1004 ( 
.A1(n_960),
.A2(n_889),
.B(n_878),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_962),
.B(n_878),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_930),
.B(n_876),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_928),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_971),
.B(n_958),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_974),
.B(n_942),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_969),
.B(n_939),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_969),
.B(n_939),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1007),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1007),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_974),
.B(n_937),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_996),
.B(n_939),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_996),
.B(n_939),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_967),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_994),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_976),
.B(n_939),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_967),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_977),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_976),
.B(n_939),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_976),
.B(n_939),
.Y(n_1023)
);

AND2x2_ASAP7_75t_SL g1024 ( 
.A(n_982),
.B(n_954),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_976),
.B(n_937),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_970),
.B(n_928),
.Y(n_1026)
);

CKINVDCx14_ASAP7_75t_R g1027 ( 
.A(n_973),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_970),
.B(n_928),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_976),
.B(n_937),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1003),
.B(n_932),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_983),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1002),
.B(n_937),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_984),
.B(n_932),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_991),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1012),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1012),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_1017),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1019),
.B(n_1002),
.Y(n_1038)
);

INVxp67_ASAP7_75t_SL g1039 ( 
.A(n_1017),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_1034),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_1021),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_1024),
.A2(n_975),
.B1(n_954),
.B2(n_989),
.Y(n_1042)
);

OAI31xp33_ASAP7_75t_L g1043 ( 
.A1(n_1027),
.A2(n_962),
.A3(n_982),
.B(n_979),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_1018),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1013),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1019),
.B(n_987),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_1018),
.B(n_972),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_1026),
.B(n_988),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1025),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1013),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_1024),
.A2(n_954),
.B1(n_978),
.B2(n_972),
.Y(n_1051)
);

NOR2xp67_ASAP7_75t_L g1052 ( 
.A(n_1019),
.B(n_1000),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1021),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1022),
.B(n_1023),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1025),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_1043),
.B(n_1024),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1048),
.B(n_1026),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_1048),
.B(n_1028),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1054),
.B(n_1022),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1042),
.B(n_1028),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1042),
.B(n_1024),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1054),
.B(n_1022),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1035),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1044),
.B(n_1023),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1038),
.B(n_1023),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_1044),
.B(n_1018),
.Y(n_1066)
);

NOR2x1_ASAP7_75t_L g1067 ( 
.A(n_1040),
.B(n_1005),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1040),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1063),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1060),
.B(n_1043),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_1068),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1058),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1064),
.B(n_1038),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_1064),
.Y(n_1074)
);

INVxp67_ASAP7_75t_SL g1075 ( 
.A(n_1067),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1059),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1069),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1070),
.A2(n_1056),
.B(n_1061),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1069),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1071),
.B(n_1058),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1071),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_1081),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1078),
.A2(n_1056),
.B1(n_1075),
.B2(n_1027),
.Y(n_1083)
);

NAND4xp25_ASAP7_75t_L g1084 ( 
.A(n_1080),
.B(n_1051),
.C(n_980),
.D(n_1072),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1079),
.A2(n_1072),
.B(n_1074),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1077),
.A2(n_1074),
.B1(n_1047),
.B2(n_1076),
.Y(n_1086)
);

OAI221xp5_ASAP7_75t_SL g1087 ( 
.A1(n_1077),
.A2(n_962),
.B1(n_1076),
.B2(n_972),
.C(n_1047),
.Y(n_1087)
);

OAI221xp5_ASAP7_75t_L g1088 ( 
.A1(n_1078),
.A2(n_1047),
.B1(n_981),
.B2(n_1044),
.C(n_1073),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1081),
.B(n_1073),
.Y(n_1089)
);

AOI211xp5_ASAP7_75t_L g1090 ( 
.A1(n_1078),
.A2(n_1004),
.B(n_1066),
.C(n_998),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_SL g1091 ( 
.A1(n_1078),
.A2(n_1066),
.B(n_1064),
.Y(n_1091)
);

NAND2xp33_ASAP7_75t_L g1092 ( 
.A(n_1078),
.B(n_1001),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1078),
.A2(n_1066),
.B(n_965),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1089),
.B(n_1082),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1085),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1092),
.A2(n_1004),
.B(n_954),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_1083),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1086),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1084),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1091),
.B(n_1065),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_1092),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1088),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_1093),
.B(n_1059),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1090),
.A2(n_954),
.B(n_1047),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1087),
.A2(n_978),
.B1(n_973),
.B2(n_999),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_1082),
.B(n_1057),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1082),
.B(n_1065),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1082),
.Y(n_1108)
);

AOI211xp5_ASAP7_75t_L g1109 ( 
.A1(n_1083),
.A2(n_965),
.B(n_998),
.C(n_978),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1108),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1104),
.A2(n_1052),
.B(n_992),
.C(n_991),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1094),
.B(n_1062),
.Y(n_1112)
);

AOI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_1097),
.A2(n_872),
.B(n_1047),
.Y(n_1113)
);

INVx3_ASAP7_75t_SL g1114 ( 
.A(n_1094),
.Y(n_1114)
);

OAI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1101),
.A2(n_1047),
.B1(n_1044),
.B2(n_999),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_1106),
.B(n_1062),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1097),
.A2(n_972),
.B(n_956),
.C(n_954),
.Y(n_1117)
);

AOI222xp33_ASAP7_75t_L g1118 ( 
.A1(n_1099),
.A2(n_1095),
.B1(n_1102),
.B2(n_1098),
.C1(n_1105),
.C2(n_1100),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_1107),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1096),
.B(n_1046),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1105),
.B(n_1046),
.Y(n_1121)
);

HAxp5_ASAP7_75t_SL g1122 ( 
.A(n_1109),
.B(n_872),
.CON(n_1122),
.SN(n_1122)
);

NAND2x1_ASAP7_75t_L g1123 ( 
.A(n_1103),
.B(n_1049),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1103),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1103),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1094),
.B(n_1052),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1094),
.B(n_1049),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1094),
.B(n_1049),
.Y(n_1128)
);

AO221x1_ASAP7_75t_L g1129 ( 
.A1(n_1115),
.A2(n_1034),
.B1(n_1055),
.B2(n_1050),
.C(n_1045),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_L g1130 ( 
.A(n_1118),
.B(n_891),
.C(n_887),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1114),
.B(n_1055),
.Y(n_1131)
);

AOI321xp33_ASAP7_75t_L g1132 ( 
.A1(n_1125),
.A2(n_956),
.A3(n_992),
.B1(n_1039),
.B2(n_966),
.C(n_968),
.Y(n_1132)
);

INVxp67_ASAP7_75t_SL g1133 ( 
.A(n_1124),
.Y(n_1133)
);

NAND2xp33_ASAP7_75t_L g1134 ( 
.A(n_1110),
.B(n_1112),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1119),
.B(n_1113),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1118),
.B(n_1055),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_SL g1137 ( 
.A(n_1117),
.B(n_881),
.C(n_888),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1111),
.B(n_865),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_1122),
.B(n_891),
.C(n_887),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1121),
.B(n_865),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1116),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_SL g1142 ( 
.A(n_1126),
.B(n_1123),
.C(n_1120),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1128),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1127),
.B(n_1041),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1118),
.A2(n_961),
.B1(n_1018),
.B2(n_995),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1133),
.B(n_1037),
.Y(n_1146)
);

OAI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_1130),
.A2(n_1039),
.B1(n_1018),
.B2(n_994),
.C(n_985),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1145),
.B(n_1139),
.Y(n_1148)
);

NAND5xp2_ASAP7_75t_L g1149 ( 
.A(n_1135),
.B(n_987),
.C(n_1010),
.D(n_1011),
.E(n_1015),
.Y(n_1149)
);

AOI222xp33_ASAP7_75t_L g1150 ( 
.A1(n_1136),
.A2(n_1025),
.B1(n_1029),
.B2(n_1037),
.C1(n_968),
.C2(n_1041),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_SL g1151 ( 
.A1(n_1141),
.A2(n_1137),
.B(n_1140),
.Y(n_1151)
);

AOI221xp5_ASAP7_75t_L g1152 ( 
.A1(n_1134),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.C(n_1041),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1142),
.A2(n_995),
.B1(n_997),
.B2(n_966),
.Y(n_1153)
);

O2A1O1Ixp5_ASAP7_75t_L g1154 ( 
.A1(n_1138),
.A2(n_1035),
.B(n_1050),
.C(n_1045),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1143),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1131),
.A2(n_997),
.B1(n_995),
.B2(n_966),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1144),
.Y(n_1157)
);

NAND4xp25_ASAP7_75t_SL g1158 ( 
.A(n_1144),
.B(n_1029),
.C(n_1036),
.D(n_1009),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1129),
.A2(n_997),
.B1(n_986),
.B2(n_1036),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1132),
.B(n_1053),
.Y(n_1160)
);

OAI221xp5_ASAP7_75t_L g1161 ( 
.A1(n_1130),
.A2(n_994),
.B1(n_985),
.B2(n_964),
.C(n_953),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_L g1162 ( 
.A(n_1130),
.B(n_886),
.C(n_876),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1130),
.B(n_1053),
.Y(n_1163)
);

OAI221xp5_ASAP7_75t_SL g1164 ( 
.A1(n_1145),
.A2(n_994),
.B1(n_968),
.B2(n_1009),
.C(n_953),
.Y(n_1164)
);

OAI221xp5_ASAP7_75t_L g1165 ( 
.A1(n_1130),
.A2(n_985),
.B1(n_964),
.B2(n_953),
.C(n_1008),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1133),
.B(n_1010),
.Y(n_1166)
);

AOI211xp5_ASAP7_75t_L g1167 ( 
.A1(n_1130),
.A2(n_1008),
.B(n_1029),
.C(n_886),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1133),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1133),
.B(n_1010),
.Y(n_1169)
);

AOI221x1_ASAP7_75t_L g1170 ( 
.A1(n_1157),
.A2(n_1030),
.B1(n_1033),
.B2(n_1031),
.C(n_1021),
.Y(n_1170)
);

NOR4xp25_ASAP7_75t_L g1171 ( 
.A(n_1151),
.B(n_1148),
.C(n_1152),
.D(n_1163),
.Y(n_1171)
);

AOI32xp33_ASAP7_75t_L g1172 ( 
.A1(n_1152),
.A2(n_1011),
.A3(n_1015),
.B1(n_1016),
.B2(n_968),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1168),
.B(n_1011),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1162),
.A2(n_1009),
.B1(n_988),
.B2(n_1030),
.Y(n_1174)
);

OAI221xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1153),
.A2(n_968),
.B1(n_953),
.B2(n_1014),
.C(n_993),
.Y(n_1175)
);

NAND3xp33_ASAP7_75t_L g1176 ( 
.A(n_1155),
.B(n_1146),
.C(n_1167),
.Y(n_1176)
);

OAI211xp5_ASAP7_75t_SL g1177 ( 
.A1(n_1147),
.A2(n_953),
.B(n_993),
.C(n_1033),
.Y(n_1177)
);

OAI211xp5_ASAP7_75t_SL g1178 ( 
.A1(n_1161),
.A2(n_953),
.B(n_963),
.C(n_951),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_1160),
.A2(n_1031),
.B1(n_963),
.B2(n_1015),
.C(n_1016),
.Y(n_1179)
);

AOI221xp5_ASAP7_75t_L g1180 ( 
.A1(n_1165),
.A2(n_1031),
.B1(n_963),
.B2(n_1016),
.C(n_986),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1154),
.A2(n_1169),
.B(n_1166),
.C(n_1164),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_L g1182 ( 
.A1(n_1149),
.A2(n_963),
.B1(n_986),
.B2(n_1020),
.C(n_932),
.Y(n_1182)
);

AOI211xp5_ASAP7_75t_L g1183 ( 
.A1(n_1158),
.A2(n_1014),
.B(n_938),
.C(n_951),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1150),
.A2(n_990),
.B(n_957),
.Y(n_1184)
);

XNOR2x1_ASAP7_75t_L g1185 ( 
.A(n_1156),
.B(n_59),
.Y(n_1185)
);

AOI211xp5_ASAP7_75t_L g1186 ( 
.A1(n_1159),
.A2(n_1014),
.B(n_938),
.C(n_951),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1168),
.A2(n_957),
.B(n_951),
.C(n_1020),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1168),
.A2(n_1020),
.B1(n_934),
.B2(n_938),
.C(n_946),
.Y(n_1188)
);

NAND3xp33_ASAP7_75t_L g1189 ( 
.A(n_1168),
.B(n_907),
.C(n_957),
.Y(n_1189)
);

OAI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1151),
.A2(n_903),
.B1(n_957),
.B2(n_934),
.C(n_950),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1148),
.A2(n_903),
.B1(n_1006),
.B2(n_1032),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1168),
.B(n_1032),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1168),
.A2(n_957),
.B(n_945),
.C(n_950),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_1176),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_1192),
.Y(n_1195)
);

NOR2xp67_ASAP7_75t_L g1196 ( 
.A(n_1173),
.B(n_60),
.Y(n_1196)
);

NAND4xp75_ASAP7_75t_L g1197 ( 
.A(n_1179),
.B(n_1180),
.C(n_1170),
.D(n_1191),
.Y(n_1197)
);

NAND4xp75_ASAP7_75t_L g1198 ( 
.A(n_1188),
.B(n_957),
.C(n_1032),
.D(n_1006),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1181),
.Y(n_1199)
);

NAND4xp75_ASAP7_75t_L g1200 ( 
.A(n_1171),
.B(n_957),
.C(n_934),
.D(n_946),
.Y(n_1200)
);

NOR2x1_ASAP7_75t_L g1201 ( 
.A(n_1185),
.B(n_62),
.Y(n_1201)
);

XNOR2xp5_ASAP7_75t_L g1202 ( 
.A(n_1186),
.B(n_63),
.Y(n_1202)
);

NOR2x1_ASAP7_75t_L g1203 ( 
.A(n_1189),
.B(n_64),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1177),
.B(n_1190),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1183),
.B(n_990),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1175),
.A2(n_903),
.B1(n_946),
.B2(n_935),
.Y(n_1206)
);

XNOR2x1_ASAP7_75t_L g1207 ( 
.A(n_1174),
.B(n_65),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1193),
.Y(n_1208)
);

NOR3xp33_ASAP7_75t_L g1209 ( 
.A(n_1178),
.B(n_1172),
.C(n_1187),
.Y(n_1209)
);

AND3x1_ASAP7_75t_L g1210 ( 
.A(n_1182),
.B(n_935),
.C(n_927),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1184),
.B(n_949),
.Y(n_1211)
);

NOR2x1_ASAP7_75t_L g1212 ( 
.A(n_1176),
.B(n_66),
.Y(n_1212)
);

NOR2x1_ASAP7_75t_L g1213 ( 
.A(n_1176),
.B(n_67),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1173),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1173),
.Y(n_1215)
);

AND4x1_ASAP7_75t_L g1216 ( 
.A(n_1212),
.B(n_68),
.C(n_69),
.D(n_71),
.Y(n_1216)
);

NAND4xp75_ASAP7_75t_L g1217 ( 
.A(n_1213),
.B(n_72),
.C(n_73),
.D(n_75),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_SL g1218 ( 
.A1(n_1194),
.A2(n_907),
.B(n_81),
.Y(n_1218)
);

AND2x4_ASAP7_75t_SL g1219 ( 
.A(n_1214),
.B(n_907),
.Y(n_1219)
);

NAND3x1_ASAP7_75t_L g1220 ( 
.A(n_1199),
.B(n_935),
.C(n_927),
.Y(n_1220)
);

NOR3xp33_ASAP7_75t_L g1221 ( 
.A(n_1201),
.B(n_1195),
.C(n_1215),
.Y(n_1221)
);

OAI221xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1209),
.A2(n_950),
.B1(n_949),
.B2(n_935),
.C(n_947),
.Y(n_1222)
);

AND4x1_ASAP7_75t_L g1223 ( 
.A(n_1203),
.B(n_80),
.C(n_83),
.D(n_84),
.Y(n_1223)
);

AOI222xp33_ASAP7_75t_L g1224 ( 
.A1(n_1208),
.A2(n_950),
.B1(n_949),
.B2(n_907),
.C1(n_930),
.C2(n_931),
.Y(n_1224)
);

NAND4xp75_ASAP7_75t_L g1225 ( 
.A(n_1196),
.B(n_85),
.C(n_94),
.D(n_95),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1207),
.B(n_96),
.Y(n_1226)
);

NAND4xp75_ASAP7_75t_L g1227 ( 
.A(n_1210),
.B(n_98),
.C(n_99),
.D(n_103),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1204),
.B(n_1202),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1200),
.B(n_950),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1197),
.B(n_105),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1220),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1216),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1221),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1230),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1226),
.B(n_1205),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1228),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1219),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1217),
.A2(n_1206),
.B1(n_1198),
.B2(n_1211),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_1218),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1222),
.A2(n_1211),
.B(n_109),
.C(n_112),
.Y(n_1240)
);

NOR2x1p5_ASAP7_75t_L g1241 ( 
.A(n_1225),
.B(n_935),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1227),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1223),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1224),
.A2(n_106),
.B(n_113),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1229),
.B(n_949),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1236),
.A2(n_935),
.B1(n_947),
.B2(n_930),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1233),
.A2(n_940),
.B1(n_947),
.B2(n_931),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1231),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1232),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1234),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1239),
.A2(n_941),
.B1(n_936),
.B2(n_943),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1243),
.A2(n_947),
.B1(n_941),
.B2(n_931),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1237),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1242),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1241),
.A2(n_944),
.B1(n_941),
.B2(n_931),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1253),
.A2(n_1238),
.B1(n_1235),
.B2(n_1244),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1248),
.A2(n_1245),
.B1(n_1240),
.B2(n_1244),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1249),
.B(n_118),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1254),
.B(n_120),
.Y(n_1259)
);

AOI22x1_ASAP7_75t_L g1260 ( 
.A1(n_1250),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1252),
.A2(n_941),
.B1(n_943),
.B2(n_936),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1258),
.A2(n_1251),
.B(n_1247),
.Y(n_1262)
);

OAI22x1_ASAP7_75t_L g1263 ( 
.A1(n_1256),
.A2(n_1246),
.B1(n_1255),
.B2(n_130),
.Y(n_1263)
);

BUFx4f_ASAP7_75t_SL g1264 ( 
.A(n_1259),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1257),
.A2(n_941),
.B1(n_943),
.B2(n_936),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1264),
.A2(n_1260),
.B1(n_1261),
.B2(n_941),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1266),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1267),
.A2(n_1263),
.B1(n_1262),
.B2(n_1265),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1268),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1269),
.A2(n_127),
.B1(n_128),
.B2(n_133),
.Y(n_1270)
);

AOI211xp5_ASAP7_75t_L g1271 ( 
.A1(n_1270),
.A2(n_136),
.B(n_137),
.C(n_142),
.Y(n_1271)
);


endmodule