module fake_jpeg_2470_n_201 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_201);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_26),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_30),
.B(n_18),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_61),
.Y(n_71)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_77),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_82),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_59),
.B1(n_70),
.B2(n_55),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_77),
.B(n_53),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_59),
.B1(n_70),
.B2(n_55),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_85),
.B(n_77),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_70),
.B1(n_55),
.B2(n_49),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_49),
.B1(n_57),
.B2(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_93),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_64),
.B1(n_65),
.B2(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_69),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_77),
.B1(n_73),
.B2(n_72),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_47),
.B1(n_41),
.B2(n_39),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_67),
.B(n_50),
.C(n_61),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_110),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_111),
.Y(n_120)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_62),
.C(n_76),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_98),
.C(n_110),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_79),
.A2(n_77),
.B(n_73),
.C(n_72),
.Y(n_107)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_1),
.B(n_2),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_84),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_109),
.A2(n_84),
.B(n_86),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_67),
.B(n_66),
.C(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_68),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_29),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_28),
.B(n_27),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_0),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_122),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_90),
.B(n_65),
.C(n_86),
.Y(n_118)
);

AO22x1_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_139)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_65),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_1),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_48),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_131),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_102),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_109),
.B(n_95),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_149),
.B(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_130),
.A2(n_95),
.B1(n_104),
.B2(n_105),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_153),
.B(n_118),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_124),
.B1(n_128),
.B2(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_2),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_140),
.B(n_123),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_32),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_144),
.C(n_148),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_31),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_120),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_3),
.B(n_4),
.Y(n_149)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_154),
.B(n_161),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_164),
.B(n_165),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_124),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_167),
.C(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_138),
.B(n_129),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_3),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_163),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_118),
.B(n_25),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_23),
.C(n_6),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_132),
.B(n_21),
.Y(n_168)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_141),
.C(n_149),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_180),
.C(n_182),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_151),
.C(n_150),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_159),
.A2(n_150),
.B1(n_151),
.B2(n_139),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_181),
.A2(n_169),
.B1(n_176),
.B2(n_162),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_134),
.C(n_8),
.Y(n_182)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_185),
.B(n_187),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_155),
.B(n_164),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_158),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_189),
.A3(n_175),
.B1(n_9),
.B2(n_10),
.C1(n_12),
.C2(n_13),
.Y(n_191)
);

OAI221xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_157),
.B1(n_134),
.B2(n_170),
.C(n_12),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_193),
.B(n_194),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_177),
.A3(n_182),
.B1(n_10),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_7),
.A3(n_9),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_17),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_192),
.B(n_183),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_197),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_16),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_17),
.B(n_19),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_20),
.B(n_199),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_20),
.Y(n_201)
);


endmodule