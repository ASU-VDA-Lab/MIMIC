module fake_jpeg_29573_n_438 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_438);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_438;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_SL g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_15),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_47),
.B(n_50),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_49),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_60),
.Y(n_95)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_64),
.Y(n_110)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_66),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_34),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_13),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_75),
.Y(n_116)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_13),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_34),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_84),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_92),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_1),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_23),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_93),
.B(n_121),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_37),
.B1(n_23),
.B2(n_31),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_98),
.B(n_57),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_105),
.A2(n_111),
.B1(n_117),
.B2(n_79),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_50),
.B(n_17),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_106),
.B(n_25),
.C(n_40),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_46),
.C(n_43),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_89),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_53),
.A2(n_37),
.B1(n_36),
.B2(n_22),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_36),
.B1(n_22),
.B2(n_41),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_48),
.B(n_17),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_56),
.B(n_31),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_142),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_51),
.B(n_24),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_137),
.B(n_141),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_55),
.A2(n_41),
.B1(n_24),
.B2(n_42),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_69),
.B1(n_3),
.B2(n_4),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_61),
.B(n_46),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_49),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_86),
.B1(n_82),
.B2(n_72),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_145),
.A2(n_157),
.B1(n_130),
.B2(n_127),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_151),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_43),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_40),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_167),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_76),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_34),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_161),
.Y(n_201)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_77),
.B1(n_41),
.B2(n_90),
.Y(n_157)
);

AO22x2_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_59),
.B1(n_25),
.B2(n_67),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_187),
.B1(n_191),
.B2(n_132),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_40),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_171),
.Y(n_204)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_94),
.B(n_34),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_95),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_163),
.B(n_164),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_110),
.B(n_99),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_96),
.B(n_34),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_181),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_166),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_105),
.A2(n_25),
.B1(n_68),
.B2(n_40),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_168),
.A2(n_174),
.B1(n_185),
.B2(n_186),
.Y(n_214)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_100),
.Y(n_172)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_144),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_173),
.Y(n_233)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_101),
.B(n_22),
.Y(n_179)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_80),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_108),
.B(n_22),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_112),
.A2(n_79),
.B1(n_80),
.B2(n_62),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_62),
.B1(n_4),
.B2(n_5),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_129),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_188)
);

AOI32xp33_ASAP7_75t_L g230 ( 
.A1(n_188),
.A2(n_97),
.A3(n_115),
.B1(n_109),
.B2(n_9),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_102),
.B(n_2),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_192),
.Y(n_215)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_118),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_120),
.B(n_2),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_102),
.B(n_6),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_189),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_194),
.A2(n_206),
.B1(n_220),
.B2(n_189),
.Y(n_246)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_197),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_200),
.A2(n_187),
.B1(n_181),
.B2(n_172),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_168),
.A2(n_174),
.B1(n_154),
.B2(n_167),
.Y(n_206)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

BUFx8_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_216),
.B(n_224),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_157),
.A2(n_120),
.B1(n_127),
.B2(n_126),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_217),
.A2(n_227),
.B1(n_177),
.B2(n_178),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_148),
.A2(n_126),
.B1(n_119),
.B2(n_133),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_155),
.B(n_133),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_192),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_152),
.A2(n_124),
.B(n_113),
.C(n_8),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_149),
.A2(n_97),
.B1(n_115),
.B2(n_113),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_188),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_152),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_238),
.B(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_239),
.Y(n_301)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_146),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_254),
.C(n_263),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_244),
.B(n_252),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_247),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_246),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_201),
.B(n_165),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_248),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_205),
.A2(n_214),
.B(n_194),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_249),
.A2(n_271),
.B(n_124),
.Y(n_296)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_251),
.Y(n_295)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_213),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_253),
.B(n_256),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_161),
.C(n_164),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_262),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_198),
.B(n_163),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_145),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

AND2x2_ASAP7_75t_SL g258 ( 
.A(n_211),
.B(n_153),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_259),
.A2(n_224),
.B(n_216),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_260),
.A2(n_264),
.B1(n_272),
.B2(n_257),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_202),
.B(n_233),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_261),
.B(n_265),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_195),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_205),
.B(n_176),
.C(n_158),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_210),
.B(n_150),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_221),
.B(n_158),
.C(n_156),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_228),
.C(n_199),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_222),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_269),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_226),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_215),
.B(n_193),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_219),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_206),
.B(n_158),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_200),
.A2(n_158),
.B1(n_162),
.B2(n_190),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_246),
.A2(n_217),
.B1(n_231),
.B2(n_215),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_274),
.A2(n_297),
.B1(n_306),
.B2(n_264),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_276),
.B(n_298),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_238),
.B(n_223),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_279),
.B(n_284),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_244),
.B(n_196),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_290),
.Y(n_312)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_160),
.C(n_235),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_288),
.C(n_294),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_287),
.A2(n_304),
.B1(n_237),
.B2(n_269),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_243),
.B(n_228),
.C(n_219),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_271),
.A2(n_209),
.B1(n_197),
.B2(n_170),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_272),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_247),
.B(n_225),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_296),
.A2(n_257),
.B(n_250),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_267),
.A2(n_209),
.B1(n_229),
.B2(n_225),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_245),
.B(n_218),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_258),
.B(n_199),
.C(n_208),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_263),
.C(n_249),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_271),
.A2(n_229),
.B1(n_180),
.B2(n_8),
.Y(n_304)
);

XOR2x2_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_281),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_279),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_310),
.Y(n_358)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_315),
.C(n_331),
.Y(n_337)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_314),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_270),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_285),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_316),
.B(n_326),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_297),
.B1(n_292),
.B2(n_299),
.Y(n_351)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_278),
.B(n_258),
.Y(n_319)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_319),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_320),
.A2(n_324),
.B1(n_287),
.B2(n_304),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_277),
.B(n_268),
.Y(n_321)
);

NOR4xp25_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_332),
.C(n_299),
.D(n_292),
.Y(n_352)
);

OAI32xp33_ASAP7_75t_L g323 ( 
.A1(n_275),
.A2(n_239),
.A3(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_327),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_274),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_324)
);

AO21x2_ASAP7_75t_SL g325 ( 
.A1(n_296),
.A2(n_237),
.B(n_273),
.Y(n_325)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_325),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_305),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_295),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_330),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_236),
.C(n_266),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_273),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_300),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_236),
.C(n_273),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_286),
.C(n_302),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_336),
.A2(n_325),
.B1(n_303),
.B2(n_11),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_312),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_340),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_322),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_342),
.B(n_345),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_344),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_284),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_308),
.B(n_288),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_348),
.C(n_350),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_308),
.B(n_275),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_354),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_313),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_351),
.A2(n_320),
.B1(n_324),
.B2(n_291),
.Y(n_363)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_329),
.B(n_276),
.Y(n_354)
);

BUFx24_ASAP7_75t_SL g360 ( 
.A(n_357),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_374),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_317),
.Y(n_361)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_338),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_362),
.B(n_370),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_363),
.A2(n_375),
.B1(n_345),
.B2(n_342),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_347),
.A2(n_314),
.B(n_310),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_365),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_309),
.Y(n_367)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_353),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_371),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_343),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_347),
.A2(n_310),
.B(n_325),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_372),
.A2(n_348),
.B(n_349),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_331),
.C(n_334),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_353),
.A2(n_323),
.B1(n_325),
.B2(n_293),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_329),
.C(n_301),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_346),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_378),
.A2(n_358),
.B1(n_355),
.B2(n_343),
.Y(n_387)
);

BUFx12f_ASAP7_75t_SL g380 ( 
.A(n_377),
.Y(n_380)
);

XNOR2x1_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_388),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_384),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_363),
.A2(n_358),
.B1(n_351),
.B2(n_354),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_387),
.A2(n_375),
.B1(n_359),
.B2(n_378),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_350),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_303),
.Y(n_389)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_389),
.Y(n_397)
);

INVx13_ASAP7_75t_L g390 ( 
.A(n_368),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_393),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_392),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_371),
.Y(n_392)
);

XNOR2x2_ASAP7_75t_SL g395 ( 
.A(n_380),
.B(n_372),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_395),
.B(n_402),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_398),
.B(n_403),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_367),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_379),
.A2(n_385),
.B1(n_394),
.B2(n_387),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_382),
.Y(n_404)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_404),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_389),
.B(n_386),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_406),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_373),
.C(n_374),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_399),
.A2(n_391),
.B(n_379),
.Y(n_407)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_407),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_403),
.B(n_384),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_410),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_401),
.B(n_393),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_397),
.A2(n_394),
.B1(n_385),
.B2(n_392),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_411),
.B(n_413),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_406),
.B(n_361),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_366),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_400),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_416),
.A2(n_395),
.B(n_373),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_417),
.B(n_423),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_415),
.B(n_396),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_424),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_388),
.C(n_400),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_414),
.C(n_410),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_409),
.B(n_382),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_420),
.A2(n_412),
.B1(n_408),
.B2(n_376),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_425),
.B(n_428),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_421),
.B(n_364),
.Y(n_429)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_429),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_426),
.B(n_419),
.C(n_421),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_431),
.A2(n_427),
.B(n_422),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_433),
.A2(n_434),
.B1(n_432),
.B2(n_390),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_430),
.A2(n_427),
.B(n_423),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_435),
.B(n_365),
.C(n_364),
.Y(n_436)
);

OAI31xp33_ASAP7_75t_L g437 ( 
.A1(n_436),
.A2(n_9),
.A3(n_10),
.B(n_11),
.Y(n_437)
);

NAND3xp33_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_9),
.C(n_11),
.Y(n_438)
);


endmodule