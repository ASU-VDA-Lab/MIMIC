module fake_jpeg_29307_n_515 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_515);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_515;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_56),
.B(n_82),
.Y(n_123)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_63),
.B(n_68),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_25),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_34),
.A2(n_7),
.B(n_11),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_69),
.A2(n_30),
.B(n_47),
.C(n_33),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_74),
.B(n_88),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_77),
.Y(n_146)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g167 ( 
.A(n_79),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_6),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_35),
.B(n_12),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g149 ( 
.A(n_89),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_16),
.B(n_6),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_90),
.B(n_28),
.Y(n_145)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_63),
.A2(n_44),
.B1(n_37),
.B2(n_42),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_110),
.A2(n_117),
.B1(n_129),
.B2(n_135),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_60),
.A2(n_44),
.B1(n_37),
.B2(n_42),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_50),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_118),
.B(n_119),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_88),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_83),
.A2(n_44),
.B1(n_39),
.B2(n_43),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_33),
.B(n_47),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_58),
.A2(n_44),
.B1(n_39),
.B2(n_43),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_50),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_140),
.B(n_0),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_24),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_61),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_154),
.A2(n_163),
.B1(n_166),
.B2(n_3),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_62),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_64),
.A2(n_28),
.B1(n_46),
.B2(n_45),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_27),
.B1(n_17),
.B2(n_32),
.Y(n_191)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_70),
.A2(n_39),
.B1(n_18),
.B2(n_30),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_103),
.C(n_101),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_177),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_146),
.A2(n_41),
.B1(n_47),
.B2(n_30),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_174),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_115),
.A2(n_99),
.B1(n_98),
.B2(n_97),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_175),
.A2(n_191),
.B1(n_163),
.B2(n_166),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_33),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_176),
.B(n_180),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_140),
.Y(n_177)
);

NOR2x1_ASAP7_75t_L g243 ( 
.A(n_178),
.B(n_149),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_48),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_107),
.A2(n_95),
.B1(n_93),
.B2(n_92),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_183),
.A2(n_186),
.B1(n_192),
.B2(n_204),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_120),
.A2(n_24),
.B1(n_46),
.B2(n_45),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_184),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_185),
.B(n_206),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_86),
.B1(n_81),
.B2(n_80),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_128),
.Y(n_187)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_146),
.A2(n_40),
.B1(n_27),
.B2(n_17),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_188),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_132),
.A2(n_79),
.B1(n_18),
.B2(n_32),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_138),
.A2(n_32),
.B1(n_38),
.B2(n_18),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_197),
.Y(n_261)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_38),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_210),
.Y(n_231)
);

BUFx2_ASAP7_75t_SL g200 ( 
.A(n_149),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_147),
.A2(n_18),
.B1(n_9),
.B2(n_12),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_201),
.A2(n_213),
.B1(n_154),
.B2(n_135),
.Y(n_254)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_202),
.Y(n_264)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_133),
.A2(n_38),
.B1(n_7),
.B2(n_10),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_159),
.A2(n_38),
.B1(n_10),
.B2(n_2),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_205),
.A2(n_212),
.B1(n_214),
.B2(n_221),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_160),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_207),
.Y(n_262)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_136),
.Y(n_208)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_118),
.B(n_160),
.Y(n_210)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_167),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_157),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_167),
.A2(n_139),
.B1(n_158),
.B2(n_171),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_220),
.Y(n_257)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_109),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_114),
.B(n_0),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_219),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_153),
.B(n_0),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_121),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_127),
.A2(n_152),
.B1(n_151),
.B2(n_148),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_110),
.B1(n_117),
.B2(n_129),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_122),
.B(n_3),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_1),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_116),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_162),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_184),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_246),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_159),
.B1(n_162),
.B2(n_137),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_233),
.A2(n_242),
.B1(n_201),
.B2(n_197),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_254),
.B1(n_204),
.B2(n_192),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_243),
.A2(n_213),
.B(n_217),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_191),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_251),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_176),
.B(n_137),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_194),
.B(n_141),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_209),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_237),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_266),
.B(n_278),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_231),
.B(n_199),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_273),
.Y(n_303)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_235),
.Y(n_268)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_290),
.B1(n_254),
.B2(n_240),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_241),
.A2(n_263),
.B1(n_226),
.B2(n_246),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_270),
.A2(n_274),
.B(n_280),
.Y(n_321)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_235),
.Y(n_271)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_272),
.A2(n_283),
.B1(n_232),
.B2(n_234),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_173),
.C(n_219),
.Y(n_273)
);

A2O1A1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_180),
.B(n_224),
.C(n_182),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_231),
.B(n_193),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_277),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_249),
.B(n_195),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_237),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_282),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_241),
.A2(n_187),
.B1(n_161),
.B2(n_216),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_281),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_186),
.B1(n_181),
.B2(n_190),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_263),
.A2(n_252),
.B1(n_242),
.B2(n_187),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_284),
.A2(n_256),
.B1(n_255),
.B2(n_253),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_285),
.A2(n_256),
.B(n_264),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_207),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_294),
.Y(n_307)
);

OAI32xp33_ASAP7_75t_L g287 ( 
.A1(n_250),
.A2(n_217),
.A3(n_202),
.B1(n_179),
.B2(n_108),
.Y(n_287)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_287),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_230),
.B(n_169),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_292),
.Y(n_310)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_261),
.A2(n_124),
.B1(n_126),
.B2(n_143),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_238),
.B(n_196),
.C(n_179),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_238),
.B(n_230),
.C(n_243),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_295),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_252),
.A2(n_211),
.B1(n_203),
.B2(n_208),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g295 ( 
.A(n_243),
.B(n_2),
.CI(n_3),
.CON(n_295),
.SN(n_295)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_306),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_298),
.A2(n_302),
.B1(n_308),
.B2(n_313),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_269),
.A2(n_232),
.B1(n_257),
.B2(n_236),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_256),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_265),
.A2(n_247),
.B1(n_240),
.B2(n_236),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_237),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_304),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_272),
.A2(n_143),
.B1(n_124),
.B2(n_126),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_245),
.B1(n_262),
.B2(n_189),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_286),
.A2(n_262),
.B1(n_225),
.B2(n_248),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_270),
.A2(n_248),
.B1(n_255),
.B2(n_227),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_323),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_316),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_317),
.A2(n_319),
.B(n_280),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_285),
.A2(n_229),
.B(n_264),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_267),
.B(n_256),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_271),
.Y(n_324)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_324),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_323),
.B(n_275),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_325),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_326),
.A2(n_328),
.B(n_347),
.Y(n_354)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_297),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_327),
.Y(n_368)
);

OAI21xp33_ASAP7_75t_SL g328 ( 
.A1(n_319),
.A2(n_304),
.B(n_321),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_311),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_329),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_273),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_330),
.B(n_293),
.C(n_291),
.Y(n_373)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_331),
.Y(n_352)
);

A2O1A1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_295),
.B(n_274),
.C(n_291),
.Y(n_333)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_333),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_316),
.B(n_307),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_334),
.A2(n_348),
.B(n_313),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_305),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_338),
.B(n_324),
.Y(n_353)
);

INVx3_ASAP7_75t_SL g339 ( 
.A(n_307),
.Y(n_339)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_339),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_311),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_343),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_307),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_345),
.Y(n_356)
);

OA21x2_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_287),
.B(n_294),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_298),
.A2(n_283),
.B1(n_292),
.B2(n_276),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_346),
.A2(n_315),
.B1(n_290),
.B2(n_288),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_319),
.A2(n_274),
.B(n_295),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_278),
.B(n_266),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_350),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_302),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_308),
.Y(n_363)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_353),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_351),
.A2(n_300),
.B1(n_322),
.B2(n_296),
.Y(n_355)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_310),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_372),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_309),
.Y(n_358)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_332),
.A2(n_309),
.B1(n_306),
.B2(n_303),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_376),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_318),
.Y(n_365)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_341),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_378),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_369),
.A2(n_335),
.B1(n_349),
.B2(n_346),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_371),
.A2(n_328),
.B(n_326),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_330),
.B(n_303),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_374),
.C(n_375),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_277),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_318),
.C(n_320),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_297),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_312),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_377),
.B(n_379),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_312),
.C(n_289),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_332),
.A2(n_279),
.B1(n_299),
.B2(n_295),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_387),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_360),
.B(n_366),
.Y(n_381)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_381),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_352),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_391),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_352),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_384),
.Y(n_411)
);

INVxp33_ASAP7_75t_L g387 ( 
.A(n_365),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_360),
.B(n_350),
.Y(n_390)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_390),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_358),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_338),
.Y(n_393)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_393),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_361),
.Y(n_394)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_394),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_359),
.B(n_336),
.Y(n_395)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_395),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_397),
.A2(n_337),
.B1(n_376),
.B2(n_339),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_368),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_398),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_368),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_400),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_355),
.A2(n_337),
.B1(n_340),
.B2(n_339),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_401),
.A2(n_356),
.B1(n_369),
.B2(n_339),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_370),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_402),
.A2(n_403),
.B1(n_341),
.B2(n_342),
.Y(n_410)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_377),
.B(n_349),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_374),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_407),
.B(n_421),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_395),
.B(n_364),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_409),
.Y(n_435)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_410),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_372),
.C(n_357),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_413),
.B(n_414),
.C(n_418),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_373),
.C(n_375),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_388),
.B(n_378),
.C(n_371),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_419),
.A2(n_397),
.B1(n_385),
.B2(n_399),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_396),
.A2(n_354),
.B1(n_334),
.B2(n_364),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_423),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_388),
.B(n_354),
.C(n_356),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_427),
.C(n_389),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_333),
.C(n_347),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_389),
.B(n_345),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_428),
.B(n_400),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_430),
.B(n_433),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_393),
.Y(n_431)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_431),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_380),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_434),
.A2(n_440),
.B1(n_423),
.B2(n_383),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_426),
.B(n_401),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_441),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_424),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_438),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_424),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_416),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_439),
.B(n_420),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_417),
.A2(n_385),
.B1(n_399),
.B2(n_391),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_382),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_425),
.B(n_414),
.Y(n_442)
);

CKINVDCx14_ASAP7_75t_R g453 ( 
.A(n_442),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_382),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_447),
.Y(n_456)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_415),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_446),
.B(n_381),
.Y(n_448)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_448),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_431),
.B(n_406),
.Y(n_449)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_449),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_445),
.B(n_407),
.C(n_386),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_451),
.B(n_452),
.C(n_459),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_419),
.C(n_412),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_433),
.A2(n_390),
.B(n_411),
.Y(n_454)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_454),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_455),
.B(n_432),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_406),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_457),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_402),
.C(n_403),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_443),
.A2(n_411),
.B(n_384),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_462),
.A2(n_443),
.B(n_422),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_463),
.B(n_392),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_441),
.B(n_427),
.C(n_421),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_444),
.C(n_434),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_436),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_327),
.C(n_299),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_466),
.B(n_470),
.Y(n_490)
);

INVx11_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_469),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_461),
.A2(n_429),
.B1(n_392),
.B2(n_460),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_473),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_432),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_474),
.B(n_478),
.C(n_452),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_476),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_450),
.A2(n_440),
.B1(n_398),
.B2(n_345),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_460),
.A2(n_345),
.B1(n_404),
.B2(n_342),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_486),
.Y(n_492)
);

NOR3xp33_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_458),
.C(n_459),
.Y(n_481)
);

NOR2x1_ASAP7_75t_L g499 ( 
.A(n_481),
.B(n_229),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_471),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_485),
.C(n_488),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_479),
.A2(n_451),
.B(n_464),
.C(n_331),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_484),
.B(n_472),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_468),
.A2(n_456),
.B1(n_398),
.B2(n_327),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_467),
.A2(n_299),
.B(n_281),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_487),
.A2(n_474),
.B(n_258),
.Y(n_498)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_469),
.Y(n_488)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_493),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_486),
.B(n_467),
.C(n_465),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_496),
.C(n_489),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_491),
.A2(n_476),
.B1(n_466),
.B2(n_478),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_495),
.A2(n_253),
.B(n_228),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_490),
.B(n_473),
.Y(n_496)
);

A2O1A1Ixp33_ASAP7_75t_SL g502 ( 
.A1(n_498),
.A2(n_499),
.B(n_481),
.C(n_484),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_229),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_500),
.B(n_482),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_502),
.B(n_503),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_504),
.B(n_494),
.C(n_492),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_505),
.A2(n_497),
.B(n_499),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_507),
.B(n_508),
.Y(n_510)
);

OAI311xp33_ASAP7_75t_L g509 ( 
.A1(n_506),
.A2(n_501),
.A3(n_495),
.B1(n_492),
.C1(n_496),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_509),
.A2(n_255),
.B(n_228),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_511),
.Y(n_512)
);

AO21x1_ASAP7_75t_L g513 ( 
.A1(n_512),
.A2(n_510),
.B(n_237),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_258),
.B(n_2),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_3),
.Y(n_515)
);


endmodule