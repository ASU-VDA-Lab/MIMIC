module fake_jpeg_15238_n_178 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_30),
.Y(n_43)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_34),
.B(n_26),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_35),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_21),
.B1(n_16),
.B2(n_26),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_27),
.B1(n_33),
.B2(n_35),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_16),
.B1(n_21),
.B2(n_23),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_35),
.B1(n_25),
.B2(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_30),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_31),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_46),
.B(n_42),
.C(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_64),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_34),
.B1(n_29),
.B2(n_16),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_27),
.B1(n_33),
.B2(n_32),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_65),
.B1(n_69),
.B2(n_38),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_15),
.B1(n_18),
.B2(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_57),
.Y(n_79)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_34),
.B(n_29),
.C(n_19),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_25),
.B1(n_26),
.B2(n_14),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_13),
.B1(n_24),
.B2(n_14),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_61),
.B(n_66),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_35),
.B1(n_28),
.B2(n_22),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_15),
.B1(n_18),
.B2(n_40),
.Y(n_76)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_25),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_36),
.A2(n_31),
.B1(n_22),
.B2(n_20),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_40),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_67),
.B(n_59),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_38),
.B1(n_20),
.B2(n_24),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_15),
.B1(n_18),
.B2(n_13),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_82),
.B1(n_63),
.B2(n_2),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_58),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_94),
.B(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_96),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_49),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_80),
.C(n_4),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_48),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_54),
.B1(n_66),
.B2(n_47),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_100),
.B1(n_71),
.B2(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_101),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_55),
.B1(n_53),
.B2(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_78),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_111),
.B1(n_2),
.B2(n_4),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_78),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_1),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_1),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_109),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_79),
.B(n_1),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_86),
.B(n_100),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_114),
.B1(n_123),
.B2(n_117),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_86),
.B(n_91),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_85),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_126),
.C(n_107),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_71),
.A3(n_82),
.B1(n_90),
.B2(n_84),
.C1(n_89),
.C2(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_121),
.Y(n_131)
);

XNOR2x2_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_71),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_96),
.B1(n_108),
.B2(n_5),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_139),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_110),
.B1(n_98),
.B2(n_103),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_122),
.B1(n_119),
.B2(n_123),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_136),
.C(n_137),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_138),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_140),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_109),
.C(n_105),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_105),
.C(n_102),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_125),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_115),
.C(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_137),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_122),
.B(n_119),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_114),
.B(n_126),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_131),
.B1(n_132),
.B2(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_159),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_149),
.B(n_147),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_157),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_133),
.Y(n_157)
);

OR2x2_ASAP7_75t_SL g165 ( 
.A(n_158),
.B(n_4),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_2),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_145),
.B1(n_146),
.B2(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_164),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_143),
.B1(n_145),
.B2(n_7),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_165),
.B(n_6),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_166),
.B(n_167),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_162),
.B(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_169),
.B(n_7),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_160),
.C(n_163),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_172),
.C(n_8),
.Y(n_174)
);

AOI31xp33_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_7),
.A3(n_8),
.B(n_9),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_174),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_9),
.B(n_10),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_11),
.Y(n_178)
);


endmodule