module real_aes_2102_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_763;
wire n_271;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_693;
wire n_496;
wire n_281;
wire n_468;
wire n_755;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_746;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_286;
wire n_416;
wire n_410;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_404;
wire n_713;
wire n_288;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_385;
wire n_275;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_668;
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_0), .A2(n_267), .B1(n_465), .B2(n_468), .Y(n_464) );
INVx1_ASAP7_75t_L g510 ( .A(n_1), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_2), .A2(n_230), .B1(n_559), .B2(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_3), .A2(n_227), .B1(n_652), .B2(n_653), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_4), .A2(n_145), .B1(n_392), .B2(n_415), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_5), .A2(n_100), .B1(n_578), .B2(n_648), .Y(n_647) );
OA22x2_ASAP7_75t_L g379 ( .A1(n_6), .A2(n_380), .B1(n_381), .B2(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_6), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_7), .A2(n_128), .B1(n_368), .B2(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_8), .A2(n_72), .B1(n_385), .B2(n_386), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_9), .A2(n_250), .B1(n_492), .B2(n_650), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_10), .A2(n_65), .B1(n_320), .B2(n_325), .Y(n_319) );
AO22x2_ASAP7_75t_L g307 ( .A1(n_11), .A2(n_201), .B1(n_297), .B2(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g708 ( .A(n_11), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_12), .A2(n_173), .B1(n_401), .B2(n_402), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_13), .A2(n_172), .B1(n_477), .B2(n_478), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_14), .A2(n_30), .B1(n_332), .B2(n_337), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_15), .A2(n_16), .B1(n_368), .B2(n_370), .Y(n_367) );
XOR2x2_ASAP7_75t_L g541 ( .A(n_17), .B(n_542), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_18), .A2(n_120), .B1(n_426), .B2(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_19), .A2(n_106), .B1(n_407), .B2(n_408), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_20), .A2(n_186), .B1(n_457), .B2(n_729), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_21), .A2(n_118), .B1(n_404), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_22), .A2(n_38), .B1(n_385), .B2(n_386), .Y(n_437) );
AO22x2_ASAP7_75t_L g304 ( .A1(n_23), .A2(n_70), .B1(n_297), .B2(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_23), .B(n_707), .Y(n_706) );
OA22x2_ASAP7_75t_L g660 ( .A1(n_24), .A2(n_661), .B1(n_674), .B2(n_675), .Y(n_660) );
INVx1_ASAP7_75t_L g674 ( .A(n_24), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_25), .A2(n_67), .B1(n_333), .B2(n_588), .Y(n_587) );
AOI22xp5_ASAP7_75t_SL g585 ( .A1(n_26), .A2(n_245), .B1(n_310), .B2(n_503), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_27), .A2(n_36), .B1(n_360), .B2(n_363), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_28), .A2(n_269), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_29), .A2(n_138), .B1(n_385), .B2(n_386), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_31), .A2(n_207), .B1(n_492), .B2(n_606), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_32), .A2(n_239), .B1(n_346), .B2(n_602), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_33), .A2(n_143), .B1(n_745), .B2(n_747), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_34), .A2(n_188), .B1(n_371), .B2(n_404), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_35), .A2(n_259), .B1(n_333), .B2(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_37), .A2(n_236), .B1(n_391), .B2(n_436), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_39), .A2(n_117), .B1(n_345), .B2(n_349), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_40), .B(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_41), .A2(n_237), .B1(n_388), .B2(n_417), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_42), .B(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_43), .A2(n_87), .B1(n_404), .B2(n_405), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_44), .A2(n_185), .B1(n_459), .B2(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_45), .A2(n_218), .B1(n_333), .B2(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_46), .A2(n_50), .B1(n_321), .B2(n_478), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_47), .A2(n_255), .B1(n_310), .B2(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_48), .A2(n_216), .B1(n_505), .B2(n_645), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_49), .A2(n_263), .B1(n_407), .B2(n_408), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_51), .A2(n_179), .B1(n_405), .B2(n_621), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_52), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_53), .A2(n_221), .B1(n_638), .B2(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_54), .A2(n_155), .B1(n_640), .B2(n_755), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_55), .A2(n_177), .B1(n_547), .B2(n_548), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_56), .A2(n_215), .B1(n_645), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_57), .A2(n_163), .B1(n_392), .B2(n_415), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_58), .A2(n_261), .B1(n_333), .B2(n_338), .Y(n_610) );
OAI22x1_ASAP7_75t_SL g632 ( .A1(n_59), .A2(n_633), .B1(n_655), .B2(n_656), .Y(n_632) );
INVx1_ASAP7_75t_L g655 ( .A(n_59), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_60), .A2(n_114), .B1(n_478), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_61), .A2(n_79), .B1(n_320), .B2(n_325), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_62), .A2(n_225), .B1(n_368), .B2(n_608), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_63), .A2(n_213), .B1(n_638), .B2(n_640), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_64), .A2(n_122), .B1(n_333), .B2(n_664), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_66), .A2(n_71), .B1(n_353), .B2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_68), .A2(n_150), .B1(n_548), .B2(n_717), .Y(n_716) );
AOI222xp33_ASAP7_75t_L g612 ( .A1(n_69), .A2(n_73), .B1(n_258), .B2(n_389), .C1(n_613), .C2(n_614), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_74), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_75), .A2(n_240), .B1(n_648), .B2(n_690), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g270 ( .A1(n_76), .A2(n_271), .B1(n_280), .B2(n_700), .C(n_710), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_77), .A2(n_208), .B1(n_345), .B2(n_347), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_78), .A2(n_209), .B1(n_392), .B2(n_415), .Y(n_414) );
AOI222xp33_ASAP7_75t_L g628 ( .A1(n_80), .A2(n_159), .B1(n_231), .B2(n_321), .C1(n_478), .C2(n_613), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_81), .A2(n_146), .B1(n_503), .B2(n_559), .Y(n_558) );
INVx3_ASAP7_75t_L g297 ( .A(n_82), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_83), .A2(n_157), .B1(n_385), .B2(n_386), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_84), .B(n_419), .Y(n_418) );
XNOR2x2_ASAP7_75t_L g410 ( .A(n_85), .B(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_86), .A2(n_252), .B1(n_577), .B2(n_578), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_88), .A2(n_232), .B1(n_388), .B2(n_417), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_89), .A2(n_158), .B1(n_401), .B2(n_402), .Y(n_448) );
INVx1_ASAP7_75t_L g513 ( .A(n_90), .Y(n_513) );
OA22x2_ASAP7_75t_L g595 ( .A1(n_91), .A2(n_596), .B1(n_597), .B2(n_615), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_91), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_92), .A2(n_109), .B1(n_372), .B2(n_580), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_93), .A2(n_130), .B1(n_550), .B2(n_551), .Y(n_549) );
AO22x2_ASAP7_75t_L g676 ( .A1(n_94), .A2(n_677), .B1(n_678), .B2(n_694), .Y(n_676) );
INVx1_ASAP7_75t_L g694 ( .A(n_94), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_95), .B(n_480), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_96), .A2(n_187), .B1(n_550), .B2(n_574), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_97), .A2(n_129), .B1(n_391), .B2(n_392), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_98), .A2(n_156), .B1(n_580), .B2(n_581), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_99), .A2(n_119), .B1(n_550), .B2(n_574), .Y(n_573) );
OA22x2_ASAP7_75t_L g735 ( .A1(n_101), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_101), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_102), .A2(n_234), .B1(n_352), .B2(n_356), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_103), .A2(n_131), .B1(n_653), .B2(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_104), .A2(n_124), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx1_ASAP7_75t_SL g298 ( .A(n_105), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_105), .B(n_127), .Y(n_709) );
INVx2_ASAP7_75t_L g276 ( .A(n_107), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_108), .A2(n_168), .B1(n_402), .B2(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_110), .A2(n_256), .B1(n_398), .B2(n_399), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_111), .A2(n_166), .B1(n_468), .B2(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_112), .A2(n_223), .B1(n_388), .B2(n_389), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_113), .A2(n_123), .B1(n_559), .B2(n_682), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_115), .A2(n_167), .B1(n_405), .B2(n_652), .Y(n_670) );
OA22x2_ASAP7_75t_L g485 ( .A1(n_116), .A2(n_486), .B1(n_487), .B2(n_514), .Y(n_485) );
INVx1_ASAP7_75t_L g514 ( .A(n_116), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_121), .A2(n_233), .B1(n_356), .B2(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_125), .A2(n_217), .B1(n_332), .B2(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_126), .A2(n_170), .B1(n_365), .B2(n_493), .Y(n_671) );
AO22x2_ASAP7_75t_L g300 ( .A1(n_127), .A2(n_210), .B1(n_297), .B2(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_132), .B(n_584), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_133), .A2(n_203), .B1(n_463), .B2(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_134), .A2(n_257), .B1(n_477), .B2(n_478), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_135), .A2(n_194), .B1(n_321), .B2(n_478), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_136), .A2(n_198), .B1(n_401), .B2(n_402), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_137), .A2(n_183), .B1(n_356), .B2(n_545), .Y(n_544) );
OA22x2_ASAP7_75t_L g285 ( .A1(n_139), .A2(n_286), .B1(n_287), .B2(n_373), .Y(n_285) );
INVx1_ASAP7_75t_L g373 ( .A(n_139), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_140), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_141), .A2(n_160), .B1(n_404), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_142), .A2(n_180), .B1(n_345), .B2(n_602), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_144), .A2(n_154), .B1(n_372), .B2(n_652), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_147), .A2(n_192), .B1(n_347), .B2(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_148), .A2(n_262), .B1(n_320), .B2(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g299 ( .A(n_149), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_151), .B(n_394), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_152), .A2(n_182), .B1(n_642), .B2(n_758), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_153), .A2(n_712), .B1(n_713), .B2(n_732), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_153), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_161), .A2(n_174), .B1(n_425), .B2(n_426), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_162), .B(n_440), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_164), .A2(n_171), .B1(n_398), .B2(n_399), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_165), .A2(n_246), .B1(n_492), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_169), .A2(n_191), .B1(n_457), .B2(n_459), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_175), .A2(n_265), .B1(n_401), .B2(n_402), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_176), .A2(n_248), .B1(n_398), .B2(n_399), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_178), .A2(n_212), .B1(n_550), .B2(n_551), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_181), .A2(n_244), .B1(n_685), .B2(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_184), .B(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_189), .A2(n_196), .B1(n_310), .B2(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_190), .A2(n_220), .B1(n_719), .B2(n_749), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_193), .A2(n_266), .B1(n_461), .B2(n_463), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_195), .A2(n_204), .B1(n_310), .B2(n_315), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_197), .B(n_291), .Y(n_561) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_199), .A2(n_211), .B1(n_493), .B2(n_523), .Y(n_522) );
XNOR2x1_ASAP7_75t_L g453 ( .A(n_200), .B(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_202), .A2(n_224), .B1(n_391), .B2(n_392), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_205), .A2(n_268), .B1(n_473), .B2(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_206), .A2(n_226), .B1(n_425), .B2(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_214), .B(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_219), .Y(n_590) );
AND2x4_ASAP7_75t_L g278 ( .A(n_222), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g704 ( .A(n_222), .Y(n_704) );
AO21x1_ASAP7_75t_L g769 ( .A1(n_222), .A2(n_274), .B(n_770), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_228), .A2(n_254), .B1(n_407), .B2(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g279 ( .A(n_229), .Y(n_279) );
AND2x2_ASAP7_75t_R g734 ( .A(n_229), .B(n_704), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_235), .B(n_290), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_238), .A2(n_247), .B1(n_338), .B2(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_241), .A2(n_253), .B1(n_321), .B2(n_326), .Y(n_586) );
INVxp67_ASAP7_75t_L g275 ( .A(n_242), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_243), .Y(n_535) );
INVx1_ASAP7_75t_L g509 ( .A(n_249), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_251), .A2(n_264), .B1(n_344), .B2(n_347), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_260), .B(n_636), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_279), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g770 ( .A(n_279), .Y(n_770) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_568), .Y(n_280) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_281), .A2(n_568), .B(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_428), .B1(n_566), .B2(n_567), .Y(n_281) );
INVx1_ASAP7_75t_L g566 ( .A(n_282), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_374), .B2(n_375), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_342), .Y(n_287) );
NAND4xp25_ASAP7_75t_SL g288 ( .A(n_289), .B(n_309), .C(n_319), .D(n_331), .Y(n_288) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx3_ASAP7_75t_SL g394 ( .A(n_292), .Y(n_394) );
INVx4_ASAP7_75t_SL g419 ( .A(n_292), .Y(n_419) );
INVx4_ASAP7_75t_SL g584 ( .A(n_292), .Y(n_584) );
INVx6_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_302), .Y(n_293) );
AND2x4_ASAP7_75t_L g317 ( .A(n_294), .B(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g339 ( .A(n_294), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g386 ( .A(n_294), .B(n_340), .Y(n_386) );
AND2x2_ASAP7_75t_L g392 ( .A(n_294), .B(n_318), .Y(n_392) );
AND2x2_ASAP7_75t_L g436 ( .A(n_294), .B(n_318), .Y(n_436) );
AND2x4_ASAP7_75t_L g440 ( .A(n_294), .B(n_302), .Y(n_440) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_300), .Y(n_294) );
INVx2_ASAP7_75t_L g314 ( .A(n_295), .Y(n_314) );
AND2x2_ASAP7_75t_L g323 ( .A(n_295), .B(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_295), .Y(n_330) );
OAI22x1_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B1(n_298), .B2(n_299), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g301 ( .A(n_297), .Y(n_301) );
INVx2_ASAP7_75t_L g305 ( .A(n_297), .Y(n_305) );
INVx1_ASAP7_75t_L g308 ( .A(n_297), .Y(n_308) );
AND2x2_ASAP7_75t_L g313 ( .A(n_300), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g324 ( .A(n_300), .Y(n_324) );
BUFx2_ASAP7_75t_L g366 ( .A(n_300), .Y(n_366) );
AND2x4_ASAP7_75t_L g346 ( .A(n_302), .B(n_323), .Y(n_346) );
AND2x4_ASAP7_75t_L g355 ( .A(n_302), .B(n_350), .Y(n_355) );
AND2x2_ASAP7_75t_L g369 ( .A(n_302), .B(n_313), .Y(n_369) );
AND2x6_ASAP7_75t_L g401 ( .A(n_302), .B(n_313), .Y(n_401) );
AND2x2_ASAP7_75t_L g407 ( .A(n_302), .B(n_323), .Y(n_407) );
AND2x2_ASAP7_75t_L g446 ( .A(n_302), .B(n_350), .Y(n_446) );
AND2x4_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g312 ( .A(n_304), .B(n_306), .Y(n_312) );
AND2x2_ASAP7_75t_L g329 ( .A(n_304), .B(n_307), .Y(n_329) );
INVx1_ASAP7_75t_L g336 ( .A(n_304), .Y(n_336) );
INVxp67_ASAP7_75t_L g318 ( .A(n_306), .Y(n_318) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g335 ( .A(n_307), .B(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx3_ASAP7_75t_L g559 ( .A(n_311), .Y(n_559) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_311), .Y(n_756) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x2_ASAP7_75t_L g322 ( .A(n_312), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g372 ( .A(n_312), .B(n_350), .Y(n_372) );
AND2x4_ASAP7_75t_L g388 ( .A(n_312), .B(n_323), .Y(n_388) );
AND2x2_ASAP7_75t_L g391 ( .A(n_312), .B(n_313), .Y(n_391) );
AND2x2_ASAP7_75t_L g415 ( .A(n_312), .B(n_313), .Y(n_415) );
AND2x2_ASAP7_75t_L g426 ( .A(n_312), .B(n_350), .Y(n_426) );
AND2x2_ASAP7_75t_L g362 ( .A(n_313), .B(n_335), .Y(n_362) );
AND2x2_ASAP7_75t_L g398 ( .A(n_313), .B(n_335), .Y(n_398) );
AND2x4_ASAP7_75t_L g350 ( .A(n_314), .B(n_324), .Y(n_350) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_SL g475 ( .A(n_316), .Y(n_475) );
INVx1_ASAP7_75t_L g503 ( .A(n_316), .Y(n_503) );
INVx2_ASAP7_75t_L g640 ( .A(n_316), .Y(n_640) );
INVx2_ASAP7_75t_L g666 ( .A(n_316), .Y(n_666) );
INVx2_ASAP7_75t_L g682 ( .A(n_316), .Y(n_682) );
INVx6_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g508 ( .A(n_320), .Y(n_508) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx5_ASAP7_75t_L g477 ( .A(n_322), .Y(n_477) );
INVx2_ASAP7_75t_L g725 ( .A(n_322), .Y(n_725) );
BUFx3_ASAP7_75t_L g759 ( .A(n_322), .Y(n_759) );
AND2x2_ASAP7_75t_L g334 ( .A(n_323), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g385 ( .A(n_323), .B(n_335), .Y(n_385) );
BUFx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx3_ASAP7_75t_L g643 ( .A(n_327), .Y(n_643) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx12f_ASAP7_75t_L g478 ( .A(n_328), .Y(n_478) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x4_ASAP7_75t_L g349 ( .A(n_329), .B(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g365 ( .A(n_329), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_SL g389 ( .A(n_329), .B(n_330), .Y(n_389) );
AND2x4_ASAP7_75t_L g399 ( .A(n_329), .B(n_366), .Y(n_399) );
AND2x4_ASAP7_75t_L g408 ( .A(n_329), .B(n_350), .Y(n_408) );
AND2x2_ASAP7_75t_SL g417 ( .A(n_329), .B(n_330), .Y(n_417) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_334), .Y(n_539) );
INVx3_ASAP7_75t_L g557 ( .A(n_334), .Y(n_557) );
AND2x4_ASAP7_75t_L g358 ( .A(n_335), .B(n_350), .Y(n_358) );
AND2x6_ASAP7_75t_L g402 ( .A(n_335), .B(n_350), .Y(n_402) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_336), .Y(n_341) );
BUFx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
BUFx6f_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
BUFx4f_ASAP7_75t_L g473 ( .A(n_339), .Y(n_473) );
INVx2_ASAP7_75t_L g506 ( .A(n_339), .Y(n_506) );
INVx1_ASAP7_75t_L g589 ( .A(n_339), .Y(n_589) );
BUFx3_ASAP7_75t_L g664 ( .A(n_339), .Y(n_664) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND4xp25_ASAP7_75t_L g342 ( .A(n_343), .B(n_351), .C(n_359), .D(n_367), .Y(n_342) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx6_ASAP7_75t_L g458 ( .A(n_346), .Y(n_458) );
BUFx3_ASAP7_75t_L g600 ( .A(n_346), .Y(n_600) );
INVx2_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_SL g548 ( .A(n_348), .Y(n_548) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g581 ( .A(n_349), .Y(n_581) );
BUFx3_ASAP7_75t_L g602 ( .A(n_349), .Y(n_602) );
BUFx2_ASAP7_75t_SL g743 ( .A(n_349), .Y(n_743) );
BUFx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
INVx3_ASAP7_75t_L g404 ( .A(n_354), .Y(n_404) );
INVx4_ASAP7_75t_L g425 ( .A(n_354), .Y(n_425) );
INVx2_ASAP7_75t_SL g470 ( .A(n_354), .Y(n_470) );
INVx3_ASAP7_75t_SL g621 ( .A(n_354), .Y(n_621) );
INVx2_ASAP7_75t_L g652 ( .A(n_354), .Y(n_652) );
INVx8_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g463 ( .A(n_357), .Y(n_463) );
INVx2_ASAP7_75t_L g578 ( .A(n_357), .Y(n_578) );
INVx2_ASAP7_75t_L g608 ( .A(n_357), .Y(n_608) );
INVx2_ASAP7_75t_L g690 ( .A(n_357), .Y(n_690) );
INVx2_ASAP7_75t_L g749 ( .A(n_357), .Y(n_749) );
INVx8_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g467 ( .A(n_362), .Y(n_467) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_362), .Y(n_550) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g574 ( .A(n_364), .Y(n_574) );
INVx2_ASAP7_75t_L g606 ( .A(n_364), .Y(n_606) );
INVx2_ASAP7_75t_L g650 ( .A(n_364), .Y(n_650) );
INVx5_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g468 ( .A(n_365), .Y(n_468) );
BUFx2_ASAP7_75t_L g523 ( .A(n_365), .Y(n_523) );
BUFx3_ASAP7_75t_L g551 ( .A(n_365), .Y(n_551) );
BUFx3_ASAP7_75t_L g648 ( .A(n_368), .Y(n_648) );
BUFx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx3_ASAP7_75t_L g462 ( .A(n_369), .Y(n_462) );
BUFx2_ASAP7_75t_L g545 ( .A(n_369), .Y(n_545) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g730 ( .A(n_371), .Y(n_730) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_372), .Y(n_405) );
BUFx3_ASAP7_75t_L g459 ( .A(n_372), .Y(n_459) );
INVx2_ASAP7_75t_L g531 ( .A(n_372), .Y(n_531) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B1(n_409), .B2(n_427), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NOR2x1_ASAP7_75t_L g382 ( .A(n_383), .B(n_395), .Y(n_382) );
NAND4xp25_ASAP7_75t_L g383 ( .A(n_384), .B(n_387), .C(n_390), .D(n_393), .Y(n_383) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_388), .Y(n_614) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_394), .Y(n_480) );
INVx2_ASAP7_75t_L g753 ( .A(n_394), .Y(n_753) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_403), .C(n_406), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_400), .Y(n_396) );
INVx1_ASAP7_75t_L g526 ( .A(n_401), .Y(n_526) );
INVx2_ASAP7_75t_L g499 ( .A(n_405), .Y(n_499) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_405), .Y(n_747) );
INVx1_ASAP7_75t_SL g427 ( .A(n_409), .Y(n_427) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_420), .Y(n_411) );
NAND4xp25_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .C(n_416), .D(n_418), .Y(n_412) );
BUFx2_ASAP7_75t_L g636 ( .A(n_419), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .C(n_423), .D(n_424), .Y(n_420) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_425), .Y(n_717) );
INVx2_ASAP7_75t_L g746 ( .A(n_425), .Y(n_746) );
INVx1_ASAP7_75t_L g567 ( .A(n_428), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_483), .B1(n_564), .B2(n_565), .Y(n_428) );
INVx1_ASAP7_75t_L g565 ( .A(n_429), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B1(n_451), .B2(n_481), .Y(n_429) );
OA22x2_ASAP7_75t_L g569 ( .A1(n_430), .A2(n_431), .B1(n_570), .B2(n_591), .Y(n_569) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
XOR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_450), .Y(n_431) );
NAND2x1_ASAP7_75t_SL g432 ( .A(n_433), .B(n_442), .Y(n_432) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_434), .B(n_438), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_441), .Y(n_438) );
INVx2_ASAP7_75t_SL g534 ( .A(n_440), .Y(n_534) );
BUFx2_ASAP7_75t_L g613 ( .A(n_440), .Y(n_613) );
NOR2x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_447), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_453), .Y(n_482) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_471), .Y(n_454) );
NAND4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_460), .C(n_464), .D(n_469), .Y(n_455) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g547 ( .A(n_458), .Y(n_547) );
INVx3_ASAP7_75t_L g580 ( .A(n_458), .Y(n_580) );
INVx1_ASAP7_75t_SL g693 ( .A(n_458), .Y(n_693) );
INVx2_ASAP7_75t_L g742 ( .A(n_458), .Y(n_742) );
INVx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g496 ( .A(n_462), .Y(n_496) );
INVx2_ASAP7_75t_L g577 ( .A(n_462), .Y(n_577) );
INVx2_ASAP7_75t_SL g719 ( .A(n_462), .Y(n_719) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g493 ( .A(n_467), .Y(n_493) );
INVx1_ASAP7_75t_L g605 ( .A(n_467), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .C(n_476), .D(n_479), .Y(n_471) );
INVx2_ASAP7_75t_L g512 ( .A(n_478), .Y(n_512) );
INVx3_ASAP7_75t_L g511 ( .A(n_480), .Y(n_511) );
INVxp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g564 ( .A(n_483), .Y(n_564) );
AOI22x1_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_515), .B2(n_516), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_500), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_494), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_497), .Y(n_494) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_507), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g686 ( .A(n_506), .Y(n_686) );
OAI222xp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_510), .B2(n_511), .C1(n_512), .C2(n_513), .Y(n_507) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OA22x2_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_541), .B1(n_562), .B2(n_563), .Y(n_516) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_517), .Y(n_563) );
XNOR2x1_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
NAND2x1p5_ASAP7_75t_L g519 ( .A(n_520), .B(n_532), .Y(n_519) );
NOR2x1_ASAP7_75t_L g520 ( .A(n_521), .B(n_527), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_524), .Y(n_521) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g553 ( .A(n_531), .Y(n_553) );
NOR2x1_ASAP7_75t_L g532 ( .A(n_533), .B(n_537), .Y(n_532) );
OAI21xp5_ASAP7_75t_SL g533 ( .A1(n_534), .A2(n_535), .B(n_536), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
BUFx6f_ASAP7_75t_SL g645 ( .A(n_539), .Y(n_645) );
INVx1_ASAP7_75t_L g562 ( .A(n_541), .Y(n_562) );
NOR2xp67_ASAP7_75t_L g542 ( .A(n_543), .B(n_554), .Y(n_542) );
NAND4xp25_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .C(n_549), .D(n_552), .Y(n_543) );
NAND4xp25_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .C(n_560), .D(n_561), .Y(n_554) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx4_ASAP7_75t_L g763 ( .A(n_557), .Y(n_763) );
INVx1_ASAP7_75t_L g639 ( .A(n_559), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_569), .A2(n_592), .B1(n_698), .B2(n_699), .Y(n_568) );
INVx2_ASAP7_75t_L g699 ( .A(n_569), .Y(n_699) );
INVx1_ASAP7_75t_SL g591 ( .A(n_570), .Y(n_591) );
XNOR2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_590), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_582), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .C(n_576), .D(n_579), .Y(n_572) );
NAND4xp25_ASAP7_75t_SL g582 ( .A(n_583), .B(n_585), .C(n_586), .D(n_587), .Y(n_582) );
INVx2_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g698 ( .A(n_592), .Y(n_698) );
AOI22xp5_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_657), .B1(n_658), .B2(n_697), .Y(n_592) );
INVx1_ASAP7_75t_SL g697 ( .A(n_593), .Y(n_697) );
XNOR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_632), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_616), .B1(n_630), .B2(n_631), .Y(n_594) );
INVx1_ASAP7_75t_L g630 ( .A(n_595), .Y(n_630) );
INVx2_ASAP7_75t_L g615 ( .A(n_597), .Y(n_615) );
NAND4xp75_ASAP7_75t_L g597 ( .A(n_598), .B(n_603), .C(n_609), .D(n_612), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_602), .Y(n_653) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_SL g631 ( .A(n_616), .Y(n_631) );
XOR2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_629), .Y(n_616) );
NAND4xp75_ASAP7_75t_L g617 ( .A(n_618), .B(n_622), .C(n_625), .D(n_628), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx2_ASAP7_75t_SL g656 ( .A(n_633), .Y(n_656) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_646), .Y(n_633) );
NAND4xp25_ASAP7_75t_SL g634 ( .A(n_635), .B(n_637), .C(n_641), .D(n_644), .Y(n_634) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND4xp25_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .C(n_651), .D(n_654), .Y(n_646) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_676), .B1(n_695), .B2(n_696), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_660), .Y(n_695) );
INVx1_ASAP7_75t_L g675 ( .A(n_661), .Y(n_675) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_662), .B(n_669), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .C(n_667), .D(n_668), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .C(n_672), .D(n_673), .Y(n_669) );
INVx4_ASAP7_75t_L g696 ( .A(n_676), .Y(n_696) );
INVx2_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_687), .Y(n_678) );
NAND4xp25_ASAP7_75t_SL g679 ( .A(n_680), .B(n_681), .C(n_683), .D(n_684), .Y(n_679) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND4xp25_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .C(n_691), .D(n_692), .Y(n_687) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_703), .B(n_706), .Y(n_766) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
OAI222xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_733), .B1(n_735), .B2(n_736), .C1(n_764), .C2(n_767), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_720), .C(n_727), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
NAND4xp25_ASAP7_75t_SL g720 ( .A(n_721), .B(n_722), .C(n_723), .D(n_726), .Y(n_720) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_731), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NOR2x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_750), .Y(n_738) );
NAND4xp25_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .C(n_744), .D(n_748), .Y(n_739) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND4xp25_ASAP7_75t_SL g750 ( .A(n_751), .B(n_754), .C(n_757), .D(n_760), .Y(n_750) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
BUFx4f_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
BUFx6f_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
CKINVDCx6p67_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_769), .Y(n_768) );
endmodule