module fake_aes_6491_n_21 (n_1, n_2, n_4, n_3, n_5, n_0, n_21);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_21;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_6;
wire n_7;
OR2x6_ASAP7_75t_L g6 ( .A(n_1), .B(n_4), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
INVx3_ASAP7_75t_L g8 ( .A(n_1), .Y(n_8) );
BUFx2_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
NOR2xp33_ASAP7_75t_L g10 ( .A(n_8), .B(n_2), .Y(n_10) );
AND2x6_ASAP7_75t_L g11 ( .A(n_8), .B(n_5), .Y(n_11) );
AND2x4_ASAP7_75t_SL g12 ( .A(n_10), .B(n_6), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_13), .B(n_9), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_15), .B(n_14), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_15), .A2(n_6), .B(n_7), .Y(n_17) );
NOR2xp67_ASAP7_75t_L g18 ( .A(n_17), .B(n_3), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_16), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AOI22xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_18), .B1(n_11), .B2(n_6), .Y(n_21) );
endmodule