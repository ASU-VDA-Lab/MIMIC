module real_jpeg_31490_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g121 ( 
.A(n_0),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_0),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_0),
.Y(n_187)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_0),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_140),
.B1(n_143),
.B2(n_144),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_1),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_1),
.A2(n_143),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_1),
.A2(n_143),
.B1(n_520),
.B2(n_522),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_2),
.A2(n_123),
.B1(n_124),
.B2(n_129),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_2),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_2),
.A2(n_123),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_2),
.A2(n_123),
.B1(n_512),
.B2(n_514),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_3),
.A2(n_62),
.B1(n_293),
.B2(n_297),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_3),
.A2(n_62),
.B1(n_383),
.B2(n_385),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_3),
.A2(n_62),
.B1(n_437),
.B2(n_441),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_5),
.A2(n_171),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_5),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_5),
.A2(n_175),
.B1(n_397),
.B2(n_507),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_6),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_6),
.A2(n_78),
.B1(n_257),
.B2(n_260),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_6),
.A2(n_78),
.B1(n_365),
.B2(n_366),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_6),
.A2(n_78),
.B1(n_397),
.B2(n_400),
.Y(n_396)
);

OAI22x1_ASAP7_75t_SL g51 ( 
.A1(n_7),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_7),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_7),
.A2(n_54),
.B1(n_112),
.B2(n_116),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_7),
.A2(n_54),
.B1(n_274),
.B2(n_277),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_7),
.A2(n_54),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_8),
.A2(n_179),
.B1(n_181),
.B2(n_184),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_8),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_8),
.A2(n_184),
.B1(n_500),
.B2(n_501),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_9),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_11),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_11),
.Y(n_180)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_11),
.Y(n_371)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_12),
.Y(n_197)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_12),
.Y(n_200)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_12),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_13),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_13),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_13),
.A2(n_242),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_13),
.A2(n_242),
.B1(n_314),
.B2(n_317),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_13),
.A2(n_242),
.B1(n_532),
.B2(n_536),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_14),
.Y(n_561)
);

OAI32xp33_ASAP7_75t_L g575 ( 
.A1(n_14),
.A2(n_493),
.A3(n_559),
.B1(n_569),
.B2(n_573),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_15),
.B(n_38),
.Y(n_160)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_15),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_15),
.B(n_69),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_15),
.A2(n_286),
.B1(n_404),
.B2(n_407),
.Y(n_403)
);

OAI32xp33_ASAP7_75t_L g411 ( 
.A1(n_15),
.A2(n_343),
.A3(n_412),
.B1(n_415),
.B2(n_422),
.Y(n_411)
);

OAI21xp33_ASAP7_75t_L g452 ( 
.A1(n_15),
.A2(n_176),
.B(n_372),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_16),
.B(n_561),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_17),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_17),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_18),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_18),
.Y(n_409)
);

OAI331xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_493),
.A3(n_559),
.B1(n_562),
.B2(n_568),
.B3(n_569),
.C1(n_570),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_20),
.A2(n_571),
.B(n_575),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_325),
.B(n_489),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_262),
.B(n_302),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_23),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_167),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_24),
.B(n_168),
.C(n_564),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_70),
.C(n_117),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_25),
.A2(n_26),
.B1(n_71),
.B2(n_72),
.Y(n_266)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_60),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_27),
.B(n_530),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_51),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g255 ( 
.A1(n_28),
.A2(n_61),
.B1(n_69),
.B2(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_28),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_28),
.B(n_256),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

AOI22x1_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_30),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_31),
.Y(n_518)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_33),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_33),
.Y(n_166)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_36),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_45),
.B2(n_49),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_48),
.Y(n_535)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_51),
.B(n_69),
.Y(n_281)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g536 ( 
.A(n_53),
.Y(n_536)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_59),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_59),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_69),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_68),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_69),
.B(n_531),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_81),
.B(n_108),
.Y(n_72)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_73),
.Y(n_290)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_77),
.Y(n_296)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22x1_ASAP7_75t_L g247 ( 
.A1(n_81),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_247)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_81),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_81),
.A2(n_108),
.B(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_82),
.B(n_111),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_82),
.A2(n_109),
.B1(n_251),
.B2(n_519),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_95),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_89),
.B2(n_93),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_89),
.B1(n_93),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_85),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_85),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_85),
.Y(n_399)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_85),
.Y(n_509)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_88),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_91),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_92),
.Y(n_219)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_99),
.B1(n_102),
.B2(n_107),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_98),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_98),
.Y(n_301)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_107),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_109),
.Y(n_249)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_111),
.Y(n_248)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_114),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_114),
.Y(n_522)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_115),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_117),
.A2(n_118),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_146),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_119),
.A2(n_146),
.B1(n_147),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_119),
.Y(n_309)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_133),
.B2(n_138),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_120),
.A2(n_133),
.B1(n_435),
.B2(n_443),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_122),
.Y(n_232)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_127),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_128),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_128),
.Y(n_378)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_132),
.Y(n_319)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_133),
.B(n_374),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g525 ( 
.A1(n_133),
.A2(n_178),
.B(n_526),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

INVx8_ASAP7_75t_L g429 ( 
.A(n_137),
.Y(n_429)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_139),
.A2(n_176),
.B1(n_233),
.B2(n_313),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_142),
.Y(n_460)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI32xp33_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_151),
.A3(n_156),
.B1(n_160),
.B2(n_161),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_160),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_229),
.Y(n_167)
);

XOR2x2_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_188),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_169),
.B(n_189),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_176),
.B1(n_177),
.B2(n_185),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_170),
.A2(n_176),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_171),
.Y(n_346)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_176),
.A2(n_364),
.B(n_372),
.Y(n_363)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_180),
.Y(n_336)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_185),
.Y(n_373)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_187),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_213),
.B1(n_220),
.B2(n_227),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_190),
.A2(n_213),
.B1(n_227),
.B2(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_SL g272 ( 
.A(n_190),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g395 ( 
.A1(n_190),
.A2(n_227),
.B1(n_382),
.B2(n_396),
.Y(n_395)
);

OAI21xp33_ASAP7_75t_SL g472 ( 
.A1(n_190),
.A2(n_355),
.B(n_396),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_190),
.A2(n_220),
.B1(n_227),
.B2(n_506),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_205),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_194),
.B1(n_198),
.B2(n_201),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVx3_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

OAI22x1_ASAP7_75t_L g205 ( 
.A1(n_198),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_203),
.Y(n_276)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_204),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_219),
.Y(n_384)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_225),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_226),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_226),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_227),
.A2(n_382),
.B(n_387),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_227),
.B(n_286),
.Y(n_447)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_228),
.A2(n_272),
.B1(n_273),
.B2(n_279),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_228),
.B(n_273),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g498 ( 
.A1(n_228),
.A2(n_272),
.B1(n_499),
.B2(n_505),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g564 ( 
.A(n_229),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_246),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_230),
.B(n_247),
.C(n_255),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_237),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_237),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx2_ASAP7_75t_R g526 ( 
.A(n_236),
.Y(n_526)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_241),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_241),
.Y(n_500)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_255),
.Y(n_246)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_249),
.A2(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_249),
.B(n_286),
.Y(n_380)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_263),
.B(n_491),
.C(n_492),
.Y(n_490)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.C(n_269),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_304)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_280),
.C(n_288),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_288),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_272),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_272),
.B(n_273),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_281),
.B(n_541),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_286),
.B(n_287),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_286),
.B(n_343),
.Y(n_342)
);

OAI21xp33_ASAP7_75t_SL g357 ( 
.A1(n_286),
.A2(n_342),
.B(n_358),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_286),
.B(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_286),
.B(n_455),
.Y(n_454)
);

AOI22x1_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_289),
.A2(n_291),
.B1(n_511),
.B2(n_519),
.Y(n_510)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_300),
.Y(n_414)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_303),
.B(n_305),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.C(n_310),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_306),
.B(n_483),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_308),
.A2(n_310),
.B1(n_311),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_308),
.Y(n_484)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_320),
.C(n_322),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_312),
.A2(n_320),
.B1(n_321),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_312),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_313),
.A2(n_427),
.B(n_430),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_319),
.Y(n_442)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XOR2x2_ASAP7_75t_L g467 ( 
.A(n_322),
.B(n_468),
.Y(n_467)
);

AOI31xp67_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_476),
.A3(n_485),
.B(n_486),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

AOI211x1_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_431),
.B(n_463),
.C(n_465),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_388),
.B(n_389),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_329),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_362),
.Y(n_329)
);

NOR2x1_ASAP7_75t_SL g388 ( 
.A(n_330),
.B(n_362),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_354),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_331),
.B(n_354),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_341),
.B1(n_345),
.B2(n_347),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_337),
.Y(n_332)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_333),
.Y(n_365)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_344),
.Y(n_425)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2x1_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_379),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_391),
.C(n_392),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_364),
.Y(n_443)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_368),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_380),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_381),
.Y(n_391)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_390),
.B(n_393),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_410),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_402),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g474 ( 
.A(n_395),
.B(n_410),
.C(n_475),
.Y(n_474)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_402),
.Y(n_475)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx5_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx8_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_409),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_426),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_411),
.B(n_426),
.Y(n_473)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx2_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx3_ASAP7_75t_SL g423 ( 
.A(n_424),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_428),
.Y(n_427)
);

INVx5_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_430),
.A2(n_436),
.B(n_449),
.Y(n_448)
);

AOI21xp33_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_445),
.B(n_462),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_444),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_434),
.B(n_444),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

BUFx2_ASAP7_75t_SL g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_446),
.A2(n_451),
.B(n_461),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_447),
.B(n_448),
.Y(n_461)
);

INVx8_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_459),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_474),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_474),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_471),
.C(n_481),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_473),
.Y(n_481)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_482),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_480),
.B(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_482),
.Y(n_488)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_493),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_557),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_547),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g558 ( 
.A(n_495),
.B(n_547),
.Y(n_558)
);

XOR2x2_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_539),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_523),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_498),
.B(n_510),
.Y(n_497)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

BUFx4f_ASAP7_75t_SL g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

XNOR2x1_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_528),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_527),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_525),
.A2(n_529),
.B1(n_537),
.B2(n_538),
.Y(n_528)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_525),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_525),
.A2(n_527),
.B1(n_538),
.B2(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_527),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_529),
.Y(n_537)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_542),
.C(n_545),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_540),
.A2(n_543),
.B1(n_544),
.B2(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_540),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_551),
.Y(n_550)
);

MAJx2_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_553),
.C(n_555),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_549),
.A2(n_550),
.B1(n_555),
.B2(n_567),
.Y(n_566)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_554),
.B(n_566),
.Y(n_565)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_555),
.Y(n_567)
);

INVxp33_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_562),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_560),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_565),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_563),
.B(n_565),
.Y(n_574)
);

NOR3xp33_ASAP7_75t_L g571 ( 
.A(n_568),
.B(n_569),
.C(n_572),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);


endmodule