module fake_jpeg_26142_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_9),
.B(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_20),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_16),
.B(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_1),
.B(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_1),
.Y(n_46)
);

AO22x2_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_18),
.B1(n_20),
.B2(n_3),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_37),
.Y(n_38)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_43),
.B1(n_38),
.B2(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_48),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_17),
.B(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_23),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_50),
.C(n_21),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_24),
.B1(n_12),
.B2(n_17),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_52),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_32),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_64),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_44),
.B1(n_48),
.B2(n_11),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_56),
.B1(n_64),
.B2(n_59),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_3),
.B(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_50),
.Y(n_67)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_63),
.C(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_70),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_38),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_52),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_53),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_78),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_79),
.B1(n_14),
.B2(n_13),
.Y(n_89)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_72),
.B(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_88),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_69),
.B1(n_67),
.B2(n_55),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_89),
.B1(n_11),
.B2(n_13),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_77),
.Y(n_88)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_93),
.Y(n_94)
);

AOI21x1_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_82),
.B(n_14),
.Y(n_92)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_91),
.A2(n_85),
.B1(n_84),
.B2(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_97),
.Y(n_98)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

OAI31xp33_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_4),
.A3(n_6),
.B(n_7),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_99),
.A2(n_100),
.B(n_8),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_7),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_102),
.Y(n_103)
);

AOI221xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_100),
.B1(n_95),
.B2(n_10),
.C(n_8),
.Y(n_104)
);


endmodule