module fake_jpeg_17467_n_184 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_14),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_35),
.Y(n_42)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_2),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_20),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_17),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_21),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_28),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_52),
.B(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_2),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_65),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_17),
.B1(n_16),
.B2(n_31),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_20),
.B1(n_17),
.B2(n_32),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_20),
.B1(n_32),
.B2(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_61),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_38),
.B1(n_30),
.B2(n_16),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_54),
.B1(n_38),
.B2(n_23),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_70),
.B1(n_75),
.B2(n_26),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_15),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_68),
.B(n_81),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_23),
.B1(n_34),
.B2(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_15),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_22),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_80),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_23),
.B1(n_22),
.B2(n_18),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_34),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_39),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_45),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_56),
.B(n_62),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_77),
.B(n_4),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_39),
.A3(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_64),
.B(n_61),
.C(n_76),
.D(n_66),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_94),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_40),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_95),
.C(n_99),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_45),
.B1(n_50),
.B2(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_50),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_45),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_63),
.B1(n_60),
.B2(n_80),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_27),
.C(n_24),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_59),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_85),
.C(n_95),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_114),
.A3(n_115),
.B1(n_86),
.B2(n_89),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_116),
.B(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_67),
.B1(n_76),
.B2(n_70),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_89),
.B(n_72),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_121),
.B(n_123),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_5),
.B(n_7),
.Y(n_139)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_126),
.C(n_127),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_90),
.B(n_83),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_128),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_83),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_102),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_102),
.C(n_99),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_129),
.C(n_130),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_98),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_122),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_93),
.C(n_92),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_88),
.C(n_100),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_135),
.B(n_138),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_142),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_133),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_145),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

OAI322xp33_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_100),
.A3(n_123),
.B1(n_111),
.B2(n_115),
.C1(n_122),
.C2(n_27),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_150),
.B(n_122),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_156),
.B(n_159),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_127),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_144),
.C(n_149),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_148),
.A2(n_117),
.B(n_110),
.Y(n_156)
);

OA21x2_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_126),
.B(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_157),
.B(n_144),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_130),
.B(n_110),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_5),
.C(n_7),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_7),
.Y(n_166)
);

XOR2x1_ASAP7_75t_SL g161 ( 
.A(n_153),
.B(n_150),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_168),
.B(n_8),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_158),
.B1(n_151),
.B2(n_155),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_162),
.B(n_163),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_8),
.C(n_10),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_25),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_172),
.Y(n_175)
);

OAI221xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_11),
.B1(n_165),
.B2(n_174),
.C(n_172),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_8),
.C(n_9),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_173),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_169),
.A2(n_165),
.B(n_10),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_11),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_170),
.C(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_176),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_181),
.Y(n_184)
);


endmodule