module fake_jpeg_3473_n_367 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_367);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_367;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_10),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_4),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_54),
.Y(n_145)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_55),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_93),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_58),
.Y(n_168)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_61),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_19),
.B(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_62),
.B(n_94),
.Y(n_176)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_8),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_65),
.B(n_87),
.Y(n_173)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_30),
.B(n_8),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_97),
.Y(n_114)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_32),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_73),
.Y(n_169)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_74),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_23),
.B(n_27),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_79),
.B(n_88),
.Y(n_172)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_23),
.B(n_8),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_89),
.B(n_90),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_91),
.B(n_92),
.Y(n_175)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_102),
.Y(n_125)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_96),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_27),
.B(n_11),
.Y(n_97)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_41),
.B1(n_34),
.B2(n_35),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_100),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_30),
.A2(n_2),
.B(n_6),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_36),
.C(n_28),
.Y(n_119)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_18),
.B(n_6),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_104),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_106),
.Y(n_146)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_41),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_108),
.Y(n_126)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_25),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_110),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_20),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_34),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_62),
.B(n_107),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_112),
.B(n_126),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g184 ( 
.A1(n_116),
.A2(n_174),
.B(n_170),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_65),
.A2(n_34),
.B1(n_18),
.B2(n_36),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_117),
.A2(n_147),
.B1(n_150),
.B2(n_165),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_119),
.B(n_130),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_33),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_28),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_140),
.B(n_143),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_97),
.A2(n_33),
.B1(n_50),
.B2(n_48),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_141),
.A2(n_154),
.B1(n_160),
.B2(n_165),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_79),
.B(n_52),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_57),
.A2(n_52),
.B1(n_50),
.B2(n_48),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_75),
.B(n_44),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_148),
.B(n_149),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_43),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_87),
.A2(n_44),
.B1(n_43),
.B2(n_37),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_37),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_153),
.B(n_175),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_84),
.A2(n_29),
.B1(n_35),
.B2(n_24),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_99),
.A2(n_24),
.B1(n_7),
.B2(n_13),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_166),
.B1(n_171),
.B2(n_168),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_14),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_159),
.B(n_164),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_100),
.A2(n_1),
.B1(n_16),
.B2(n_104),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_69),
.B(n_1),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_93),
.A2(n_63),
.B1(n_86),
.B2(n_91),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_80),
.A2(n_85),
.B1(n_82),
.B2(n_70),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_90),
.A2(n_75),
.B1(n_47),
.B2(n_73),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_170),
.A2(n_132),
.B1(n_167),
.B2(n_175),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_78),
.A2(n_84),
.B1(n_57),
.B2(n_55),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_62),
.A2(n_88),
.B1(n_97),
.B2(n_23),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_176),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_180),
.B(n_182),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_112),
.B(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_188),
.Y(n_232)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_114),
.B(n_173),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_190),
.B(n_198),
.Y(n_246)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_191),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_192),
.B(n_205),
.Y(n_256)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_193),
.Y(n_269)
);

BUFx2_ASAP7_75t_SL g194 ( 
.A(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_194),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_195),
.B(n_203),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_197),
.B(n_199),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_137),
.B(n_145),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_115),
.B(n_125),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_207),
.Y(n_236)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_133),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_167),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_216),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_SL g209 ( 
.A1(n_160),
.A2(n_171),
.B(n_150),
.C(n_116),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_SL g260 ( 
.A1(n_209),
.A2(n_210),
.B(n_225),
.C(n_211),
.Y(n_260)
);

BUFx8_ASAP7_75t_L g211 ( 
.A(n_131),
.Y(n_211)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_144),
.A2(n_133),
.B1(n_128),
.B2(n_138),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_213),
.A2(n_222),
.B1(n_229),
.B2(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_127),
.B(n_128),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_217),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_178),
.B1(n_231),
.B2(n_179),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_127),
.B(n_118),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_113),
.A2(n_121),
.B(n_151),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_182),
.B(n_203),
.C(n_190),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_152),
.B(n_139),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_231),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_113),
.B(n_152),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_177),
.A2(n_124),
.B1(n_135),
.B2(n_121),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_177),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_224),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_120),
.B(n_129),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_131),
.B(n_120),
.C(n_129),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_226),
.Y(n_262)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_135),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_158),
.B(n_131),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_230),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_158),
.A2(n_87),
.B1(n_166),
.B2(n_107),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_202),
.B1(n_188),
.B2(n_204),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_171),
.A2(n_157),
.B1(n_94),
.B2(n_155),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_157),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_241),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_L g275 ( 
.A1(n_242),
.A2(n_260),
.B(n_232),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_247),
.A2(n_250),
.B1(n_252),
.B2(n_268),
.Y(n_292)
);

OA22x2_ASAP7_75t_SL g248 ( 
.A1(n_209),
.A2(n_180),
.B1(n_195),
.B2(n_215),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_248),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_195),
.A2(n_181),
.B1(n_198),
.B2(n_217),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_212),
.A2(n_184),
.B1(n_214),
.B2(n_220),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_251),
.A2(n_246),
.B1(n_237),
.B2(n_238),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_206),
.A2(n_191),
.B1(n_226),
.B2(n_193),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_189),
.B(n_200),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_196),
.B(n_183),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_233),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_185),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_211),
.B(n_207),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_271),
.B(n_289),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_186),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_261),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_278),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_250),
.C(n_261),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_281),
.C(n_282),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_275),
.A2(n_296),
.B1(n_236),
.B2(n_253),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_244),
.B(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_276),
.B(n_287),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_261),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_257),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_237),
.B(n_238),
.C(n_262),
.Y(n_281)
);

XOR2x2_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_292),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_258),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_249),
.B(n_263),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_252),
.B(n_268),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_293),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_232),
.A2(n_235),
.B(n_248),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_232),
.C(n_239),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_295),
.C(n_253),
.Y(n_304)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_243),
.Y(n_291)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_260),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_256),
.A2(n_241),
.B1(n_260),
.B2(n_243),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_294),
.A2(n_245),
.B1(n_270),
.B2(n_284),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_269),
.B(n_260),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_269),
.A2(n_234),
.B1(n_240),
.B2(n_255),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_299),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_276),
.B(n_266),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_311),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_281),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_270),
.A2(n_245),
.B1(n_264),
.B2(n_292),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_310),
.B1(n_271),
.B2(n_278),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_296),
.Y(n_309)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_309),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_290),
.B(n_284),
.CI(n_282),
.CON(n_311),
.SN(n_311)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_288),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_314),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_279),
.B(n_280),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_320),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_308),
.B(n_293),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_316),
.A2(n_312),
.B(n_313),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_322),
.C(n_324),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_314),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_318),
.B(n_319),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_305),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_298),
.A2(n_294),
.B1(n_285),
.B2(n_289),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_274),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_282),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_295),
.C(n_273),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_304),
.C(n_301),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_298),
.A2(n_283),
.B1(n_277),
.B2(n_272),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_309),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_287),
.Y(n_329)
);

OA21x2_ASAP7_75t_SL g340 ( 
.A1(n_329),
.A2(n_286),
.B(n_300),
.Y(n_340)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_331),
.A2(n_333),
.B1(n_335),
.B2(n_336),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_337),
.Y(n_348)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_328),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_297),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_326),
.C(n_322),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_340),
.B(n_341),
.Y(n_344)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_317),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_347),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_343),
.B(n_345),
.Y(n_352)
);

AOI321xp33_ASAP7_75t_L g345 ( 
.A1(n_331),
.A2(n_307),
.A3(n_321),
.B1(n_301),
.B2(n_324),
.C(n_316),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_330),
.B(n_304),
.Y(n_347)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_338),
.Y(n_349)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_349),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_297),
.C(n_295),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_350),
.B(n_332),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_344),
.A2(n_333),
.B1(n_335),
.B2(n_325),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_348),
.Y(n_359)
);

OAI221xp5_ASAP7_75t_L g358 ( 
.A1(n_355),
.A2(n_347),
.B1(n_346),
.B2(n_343),
.C(n_350),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_334),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_356),
.B(n_334),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_354),
.B(n_349),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_357),
.A2(n_358),
.B(n_352),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_359),
.A2(n_337),
.B(n_300),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_360),
.B(n_356),
.C(n_310),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_361),
.A2(n_351),
.B(n_336),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_362),
.B(n_363),
.C(n_360),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_364),
.A2(n_365),
.B(n_351),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_366),
.A2(n_302),
.B(n_306),
.Y(n_367)
);


endmodule