module fake_jpeg_3092_n_281 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_49),
.Y(n_89)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_44),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_24),
.B(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_51),
.Y(n_120)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_26),
.B(n_22),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_54),
.B(n_60),
.Y(n_113)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_26),
.B(n_1),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_32),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_14),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_27),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_27),
.B(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_67),
.B(n_71),
.Y(n_100)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_17),
.B(n_2),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_58),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_79),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_L g78 ( 
.A(n_18),
.B(n_2),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_5),
.B1(n_8),
.B2(n_11),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_95),
.B(n_98),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_39),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_107),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_50),
.A2(n_21),
.B1(n_38),
.B2(n_37),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_101),
.A2(n_117),
.B1(n_56),
.B2(n_72),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_62),
.A2(n_39),
.B1(n_31),
.B2(n_21),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_103),
.A2(n_93),
.B1(n_120),
.B2(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_31),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_63),
.B(n_48),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_108),
.Y(n_154)
);

NAND2xp67_ASAP7_75t_SL g112 ( 
.A(n_80),
.B(n_38),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_55),
.B(n_36),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_57),
.A2(n_37),
.B1(n_36),
.B2(n_8),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_58),
.B(n_3),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_124),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_45),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_122),
.A2(n_118),
.B1(n_121),
.B2(n_104),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_46),
.B(n_77),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_111),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_133),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_110),
.B(n_87),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_154),
.B(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_68),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_138),
.B(n_139),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_59),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_142),
.B(n_143),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_81),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_147),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_146),
.A2(n_164),
.B1(n_161),
.B2(n_157),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_75),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_152),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_51),
.B1(n_77),
.B2(n_42),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_150),
.A2(n_151),
.B1(n_163),
.B2(n_156),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_104),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_89),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_114),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_157),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_160),
.Y(n_194)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_162),
.Y(n_186)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_120),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_83),
.C(n_123),
.Y(n_179)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_97),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_117),
.B1(n_122),
.B2(n_114),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_166),
.A2(n_183),
.B1(n_185),
.B2(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_172),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_153),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_137),
.B(n_134),
.C(n_132),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_83),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_141),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_165),
.C(n_161),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_96),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_156),
.A2(n_96),
.B1(n_123),
.B2(n_151),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_135),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_190),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_158),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_160),
.B1(n_149),
.B2(n_128),
.Y(n_193)
);

AO22x1_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_188),
.B1(n_178),
.B2(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_194),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_210),
.C(n_211),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_177),
.B(n_144),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_179),
.C(n_191),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_172),
.A2(n_126),
.B1(n_162),
.B2(n_167),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_208),
.B1(n_212),
.B2(n_216),
.Y(n_218)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_174),
.C(n_178),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_178),
.C(n_188),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_183),
.B1(n_175),
.B2(n_184),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_171),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_169),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_176),
.B1(n_168),
.B2(n_182),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_212),
.B1(n_202),
.B2(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_226),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_216),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_222),
.B(n_214),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_205),
.Y(n_238)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_186),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_193),
.Y(n_230)
);

OAI21x1_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_233),
.B(n_195),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_210),
.C(n_200),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_231),
.B(n_195),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_193),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_232),
.B(n_199),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_236),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_234),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_217),
.C(n_229),
.Y(n_251)
);

OAI322xp33_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_240),
.A3(n_227),
.B1(n_226),
.B2(n_223),
.C1(n_230),
.C2(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_205),
.C(n_206),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_214),
.B(n_206),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_245),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_233),
.B1(n_225),
.B2(n_219),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_231),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_251),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_252),
.A2(n_254),
.B1(n_243),
.B2(n_242),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_221),
.B1(n_218),
.B2(n_220),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_246),
.A2(n_218),
.B1(n_220),
.B2(n_217),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_241),
.B1(n_242),
.B2(n_247),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_189),
.C(n_191),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_256),
.B(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_261),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_257),
.B(n_255),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_254),
.A2(n_240),
.B1(n_204),
.B2(n_193),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_249),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_170),
.B(n_252),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_256),
.B(n_170),
.Y(n_268)
);

NAND4xp25_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_257),
.C(n_250),
.D(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_267),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_270),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_260),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_263),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_273),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_260),
.C(n_258),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_266),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_272),
.C(n_275),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_271),
.A2(n_262),
.B(n_273),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_279),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_278),
.Y(n_281)
);


endmodule