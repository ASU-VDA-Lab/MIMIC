module real_aes_6213_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_148;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_0), .B(n_110), .C(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g449 ( .A(n_0), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_1), .A2(n_137), .B(n_141), .C(n_236), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_2), .A2(n_173), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g470 ( .A(n_3), .Y(n_470) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_4), .A2(n_457), .B1(n_737), .B2(n_740), .C1(n_743), .C2(n_744), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_5), .B(n_213), .Y(n_270) );
AOI21xp33_ASAP7_75t_L g497 ( .A1(n_6), .A2(n_173), .B(n_498), .Y(n_497) );
AND2x6_ASAP7_75t_L g137 ( .A(n_7), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g196 ( .A(n_8), .Y(n_196) );
INVx1_ASAP7_75t_L g107 ( .A(n_9), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_9), .B(n_40), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_10), .A2(n_172), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_11), .B(n_149), .Y(n_240) );
INVx1_ASAP7_75t_L g502 ( .A(n_12), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_13), .B(n_207), .Y(n_525) );
INVx1_ASAP7_75t_L g157 ( .A(n_14), .Y(n_157) );
INVx1_ASAP7_75t_L g547 ( .A(n_15), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_16), .A2(n_147), .B(n_221), .C(n_223), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_17), .B(n_213), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_18), .B(n_481), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_19), .B(n_173), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_20), .B(n_186), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_21), .A2(n_207), .B(n_208), .C(n_210), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_22), .B(n_213), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_23), .B(n_149), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_24), .A2(n_181), .B(n_223), .C(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_25), .B(n_149), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g253 ( .A(n_26), .Y(n_253) );
INVx1_ASAP7_75t_L g145 ( .A(n_27), .Y(n_145) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_28), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_29), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_30), .B(n_149), .Y(n_471) );
INVx1_ASAP7_75t_L g179 ( .A(n_31), .Y(n_179) );
INVx1_ASAP7_75t_L g492 ( .A(n_32), .Y(n_492) );
INVx2_ASAP7_75t_L g135 ( .A(n_33), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_34), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_35), .A2(n_207), .B(n_266), .C(n_268), .Y(n_265) );
INVxp67_ASAP7_75t_L g180 ( .A(n_36), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_37), .A2(n_141), .B(n_144), .C(n_152), .Y(n_140) );
CKINVDCx14_ASAP7_75t_R g264 ( .A(n_38), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_39), .A2(n_137), .B(n_141), .C(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_40), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g491 ( .A(n_41), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_42), .A2(n_194), .B(n_195), .C(n_197), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_43), .B(n_149), .Y(n_537) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_44), .A2(n_47), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_44), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_45), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_46), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_47), .Y(n_123) );
INVx1_ASAP7_75t_L g205 ( .A(n_48), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_49), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_50), .B(n_173), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_51), .A2(n_141), .B1(n_210), .B2(n_490), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_52), .A2(n_102), .B1(n_114), .B2(n_747), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_53), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_54), .Y(n_467) );
CKINVDCx14_ASAP7_75t_R g192 ( .A(n_55), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_56), .A2(n_194), .B(n_268), .C(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_57), .Y(n_540) );
INVx1_ASAP7_75t_L g499 ( .A(n_58), .Y(n_499) );
INVx1_ASAP7_75t_L g138 ( .A(n_59), .Y(n_138) );
INVx1_ASAP7_75t_L g156 ( .A(n_60), .Y(n_156) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_61), .A2(n_90), .B1(n_738), .B2(n_739), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_61), .Y(n_738) );
INVx1_ASAP7_75t_SL g267 ( .A(n_62), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_63), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_64), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_65), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g256 ( .A(n_66), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_SL g480 ( .A1(n_67), .A2(n_268), .B(n_481), .C(n_482), .Y(n_480) );
INVxp67_ASAP7_75t_L g483 ( .A(n_68), .Y(n_483) );
INVx1_ASAP7_75t_L g113 ( .A(n_69), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_70), .A2(n_173), .B(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_71), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_72), .A2(n_173), .B(n_218), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_73), .Y(n_495) );
INVx1_ASAP7_75t_L g534 ( .A(n_74), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_75), .A2(n_172), .B(n_174), .Y(n_171) );
CKINVDCx16_ASAP7_75t_R g139 ( .A(n_76), .Y(n_139) );
INVx1_ASAP7_75t_L g219 ( .A(n_77), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_78), .A2(n_137), .B(n_141), .C(n_536), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_79), .A2(n_173), .B(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g222 ( .A(n_80), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_81), .B(n_146), .Y(n_516) );
INVx2_ASAP7_75t_L g154 ( .A(n_82), .Y(n_154) );
INVx1_ASAP7_75t_L g237 ( .A(n_83), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_84), .B(n_481), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_85), .A2(n_137), .B(n_141), .C(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g110 ( .A(n_86), .Y(n_110) );
OR2x2_ASAP7_75t_L g446 ( .A(n_86), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g736 ( .A(n_86), .B(n_448), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_87), .A2(n_141), .B(n_255), .C(n_258), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_88), .B(n_153), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_89), .Y(n_474) );
CKINVDCx14_ASAP7_75t_R g739 ( .A(n_90), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_91), .A2(n_137), .B(n_141), .C(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_92), .Y(n_529) );
INVx1_ASAP7_75t_L g479 ( .A(n_93), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_94), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_95), .B(n_146), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_96), .B(n_161), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_97), .B(n_161), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_98), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g209 ( .A(n_99), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_100), .A2(n_173), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g747 ( .A(n_104), .Y(n_747) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g734 ( .A(n_110), .B(n_448), .Y(n_734) );
NOR2x2_ASAP7_75t_L g744 ( .A(n_110), .B(n_447), .Y(n_744) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_455), .Y(n_114) );
BUFx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g746 ( .A(n_118), .Y(n_746) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_443), .B(n_451), .Y(n_120) );
XNOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
INVx1_ASAP7_75t_SL g735 ( .A(n_125), .Y(n_735) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_125), .A2(n_459), .B1(n_732), .B2(n_741), .Y(n_740) );
OR5x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_337), .C(n_401), .D(n_417), .E(n_432), .Y(n_125) );
NAND4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_271), .C(n_298), .D(n_321), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_214), .B(n_225), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_163), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx3_ASAP7_75t_SL g248 ( .A(n_130), .Y(n_248) );
AND2x4_ASAP7_75t_L g284 ( .A(n_130), .B(n_273), .Y(n_284) );
OR2x2_ASAP7_75t_L g294 ( .A(n_130), .B(n_250), .Y(n_294) );
OR2x2_ASAP7_75t_L g340 ( .A(n_130), .B(n_166), .Y(n_340) );
AND2x2_ASAP7_75t_L g354 ( .A(n_130), .B(n_249), .Y(n_354) );
AND2x2_ASAP7_75t_L g397 ( .A(n_130), .B(n_287), .Y(n_397) );
AND2x2_ASAP7_75t_L g404 ( .A(n_130), .B(n_261), .Y(n_404) );
AND2x2_ASAP7_75t_L g423 ( .A(n_130), .B(n_313), .Y(n_423) );
AND2x2_ASAP7_75t_L g441 ( .A(n_130), .B(n_283), .Y(n_441) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_158), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_139), .B(n_140), .C(n_153), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_132), .A2(n_234), .B(n_235), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_132), .A2(n_253), .B(n_254), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_132), .A2(n_467), .B(n_468), .Y(n_466) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_132), .A2(n_183), .B1(n_489), .B2(n_493), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_132), .A2(n_534), .B(n_535), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
AND2x4_ASAP7_75t_L g173 ( .A(n_133), .B(n_137), .Y(n_173) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g151 ( .A(n_134), .Y(n_151) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g142 ( .A(n_135), .Y(n_142) );
INVx1_ASAP7_75t_L g211 ( .A(n_135), .Y(n_211) );
INVx1_ASAP7_75t_L g143 ( .A(n_136), .Y(n_143) );
INVx3_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_136), .Y(n_182) );
INVx1_ASAP7_75t_L g481 ( .A(n_136), .Y(n_481) );
BUFx3_ASAP7_75t_L g152 ( .A(n_137), .Y(n_152) );
INVx4_ASAP7_75t_SL g183 ( .A(n_137), .Y(n_183) );
INVx5_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx3_ASAP7_75t_L g198 ( .A(n_142), .Y(n_198) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_142), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_148), .C(n_150), .Y(n_144) );
OAI22xp33_ASAP7_75t_L g178 ( .A1(n_146), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_146), .A2(n_470), .B(n_471), .C(n_472), .Y(n_469) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_147), .B(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_147), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_147), .B(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
INVx4_ASAP7_75t_L g207 ( .A(n_149), .Y(n_207) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_151), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_153), .A2(n_190), .B(n_199), .Y(n_189) );
INVx1_ASAP7_75t_L g232 ( .A(n_153), .Y(n_232) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_153), .A2(n_542), .B(n_548), .Y(n_541) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AND2x2_ASAP7_75t_L g162 ( .A(n_154), .B(n_155), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx3_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_160), .B(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_160), .A2(n_252), .B(n_259), .Y(n_251) );
NOR2xp33_ASAP7_75t_SL g518 ( .A(n_160), .B(n_519), .Y(n_518) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_161), .A2(n_477), .B(n_484), .Y(n_476) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g169 ( .A(n_162), .Y(n_169) );
INVx1_ASAP7_75t_L g406 ( .A(n_163), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_188), .Y(n_163) );
AND2x2_ASAP7_75t_L g316 ( .A(n_164), .B(n_249), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_164), .B(n_336), .Y(n_335) );
AOI32xp33_ASAP7_75t_L g349 ( .A1(n_164), .A2(n_350), .A3(n_353), .B1(n_355), .B2(n_359), .Y(n_349) );
AND2x2_ASAP7_75t_L g419 ( .A(n_164), .B(n_313), .Y(n_419) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g283 ( .A(n_166), .B(n_250), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_166), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g325 ( .A(n_166), .B(n_272), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_166), .B(n_404), .Y(n_403) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_184), .Y(n_166) );
INVx1_ASAP7_75t_L g288 ( .A(n_167), .Y(n_288) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_167), .A2(n_533), .B(n_539), .Y(n_532) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_SL g512 ( .A1(n_168), .A2(n_513), .B(n_514), .Y(n_512) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_169), .A2(n_466), .B(n_473), .Y(n_465) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_169), .A2(n_488), .B(n_494), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_169), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_171), .A2(n_185), .B(n_288), .Y(n_287) );
BUFx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_183), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_SL g191 ( .A1(n_176), .A2(n_183), .B(n_192), .C(n_193), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_SL g204 ( .A1(n_176), .A2(n_183), .B(n_205), .C(n_206), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_SL g218 ( .A1(n_176), .A2(n_183), .B(n_219), .C(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_176), .A2(n_183), .B(n_264), .C(n_265), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_176), .A2(n_183), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_176), .A2(n_183), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_176), .A2(n_183), .B(n_544), .C(n_545), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_181), .B(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_181), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_181), .B(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g239 ( .A(n_182), .Y(n_239) );
OAI22xp5_ASAP7_75t_SL g490 ( .A1(n_182), .A2(n_239), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g258 ( .A(n_183), .Y(n_258) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_187), .B(n_260), .Y(n_259) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_187), .A2(n_521), .B(n_528), .Y(n_520) );
AND2x2_ASAP7_75t_L g290 ( .A(n_188), .B(n_229), .Y(n_290) );
AND2x2_ASAP7_75t_L g366 ( .A(n_188), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g438 ( .A(n_188), .Y(n_438) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_200), .Y(n_188) );
OR2x2_ASAP7_75t_L g228 ( .A(n_189), .B(n_201), .Y(n_228) );
AND2x2_ASAP7_75t_L g245 ( .A(n_189), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_189), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g297 ( .A(n_189), .Y(n_297) );
AND2x2_ASAP7_75t_L g324 ( .A(n_189), .B(n_201), .Y(n_324) );
BUFx3_ASAP7_75t_L g327 ( .A(n_189), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_189), .B(n_302), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_189), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g241 ( .A(n_197), .Y(n_241) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g223 ( .A(n_198), .Y(n_223) );
INVx2_ASAP7_75t_L g278 ( .A(n_200), .Y(n_278) );
AND2x2_ASAP7_75t_L g296 ( .A(n_200), .B(n_276), .Y(n_296) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g307 ( .A(n_201), .B(n_216), .Y(n_307) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_201), .Y(n_320) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_212), .Y(n_201) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_202), .A2(n_217), .B(n_224), .Y(n_216) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_202), .A2(n_262), .B(n_270), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_207), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g472 ( .A(n_210), .Y(n_472) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_213), .A2(n_497), .B(n_503), .Y(n_496) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_215), .B(n_327), .Y(n_377) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_SL g246 ( .A(n_216), .Y(n_246) );
NAND3xp33_ASAP7_75t_L g295 ( .A(n_216), .B(n_296), .C(n_297), .Y(n_295) );
OR2x2_ASAP7_75t_L g303 ( .A(n_216), .B(n_276), .Y(n_303) );
AND2x2_ASAP7_75t_L g323 ( .A(n_216), .B(n_276), .Y(n_323) );
AND2x2_ASAP7_75t_L g367 ( .A(n_216), .B(n_231), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_244), .B(n_247), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_227), .B(n_229), .Y(n_226) );
AND2x2_ASAP7_75t_L g442 ( .A(n_227), .B(n_367), .Y(n_442) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_228), .A2(n_340), .B1(n_382), .B2(n_384), .Y(n_381) );
OR2x2_ASAP7_75t_L g388 ( .A(n_228), .B(n_303), .Y(n_388) );
OR2x2_ASAP7_75t_L g412 ( .A(n_228), .B(n_413), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_228), .B(n_332), .Y(n_425) );
AND2x2_ASAP7_75t_L g318 ( .A(n_229), .B(n_319), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_229), .A2(n_391), .B(n_406), .Y(n_405) );
AOI32xp33_ASAP7_75t_L g426 ( .A1(n_229), .A2(n_316), .A3(n_427), .B1(n_429), .B2(n_430), .Y(n_426) );
OR2x2_ASAP7_75t_L g437 ( .A(n_229), .B(n_438), .Y(n_437) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g305 ( .A(n_230), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_230), .B(n_319), .Y(n_384) );
BUFx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx4_ASAP7_75t_L g276 ( .A(n_231), .Y(n_276) );
AND2x2_ASAP7_75t_L g342 ( .A(n_231), .B(n_307), .Y(n_342) );
AND3x2_ASAP7_75t_L g351 ( .A(n_231), .B(n_245), .C(n_352), .Y(n_351) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_242), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_232), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_232), .B(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_232), .B(n_540), .Y(n_539) );
O2A1O1Ixp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_240), .C(n_241), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_238), .A2(n_241), .B(n_256), .C(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_241), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_241), .A2(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g277 ( .A(n_246), .B(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_246), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_246), .B(n_276), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
AND2x2_ASAP7_75t_L g272 ( .A(n_248), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g312 ( .A(n_248), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g330 ( .A(n_248), .B(n_261), .Y(n_330) );
AND2x2_ASAP7_75t_L g348 ( .A(n_248), .B(n_250), .Y(n_348) );
OR2x2_ASAP7_75t_L g362 ( .A(n_248), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g408 ( .A(n_248), .B(n_336), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_249), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_261), .Y(n_249) );
AND2x2_ASAP7_75t_L g309 ( .A(n_250), .B(n_287), .Y(n_309) );
OR2x2_ASAP7_75t_L g363 ( .A(n_250), .B(n_287), .Y(n_363) );
AND2x2_ASAP7_75t_L g416 ( .A(n_250), .B(n_273), .Y(n_416) );
INVx2_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
BUFx2_ASAP7_75t_L g314 ( .A(n_251), .Y(n_314) );
AND2x2_ASAP7_75t_L g336 ( .A(n_251), .B(n_261), .Y(n_336) );
INVx2_ASAP7_75t_L g273 ( .A(n_261), .Y(n_273) );
INVx1_ASAP7_75t_L g293 ( .A(n_261), .Y(n_293) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_269), .Y(n_526) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_274), .B(n_279), .C(n_291), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_272), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g435 ( .A(n_272), .Y(n_435) );
AND2x2_ASAP7_75t_L g313 ( .A(n_273), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_276), .B(n_277), .Y(n_285) );
INVx1_ASAP7_75t_L g370 ( .A(n_276), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_276), .B(n_297), .Y(n_394) );
AND2x2_ASAP7_75t_L g410 ( .A(n_276), .B(n_324), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_277), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g301 ( .A(n_278), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_285), .B1(n_286), .B2(n_289), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_282), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_283), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g308 ( .A(n_284), .B(n_309), .Y(n_308) );
AOI221xp5_ASAP7_75t_SL g373 ( .A1(n_284), .A2(n_326), .B1(n_374), .B2(n_379), .C(n_381), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_284), .B(n_347), .Y(n_380) );
INVx1_ASAP7_75t_L g440 ( .A(n_286), .Y(n_440) );
BUFx3_ASAP7_75t_L g347 ( .A(n_287), .Y(n_347) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI21xp33_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_294), .B(n_295), .Y(n_291) );
INVx1_ASAP7_75t_L g356 ( .A(n_293), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_293), .B(n_347), .Y(n_400) );
INVx1_ASAP7_75t_L g357 ( .A(n_294), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_294), .B(n_347), .Y(n_358) );
INVxp67_ASAP7_75t_L g378 ( .A(n_296), .Y(n_378) );
AND2x2_ASAP7_75t_L g319 ( .A(n_297), .B(n_320), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_304), .B(n_308), .C(n_310), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_SL g333 ( .A(n_301), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_302), .B(n_333), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_302), .B(n_324), .Y(n_375) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_305), .A2(n_311), .B1(n_315), .B2(n_317), .Y(n_310) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g326 ( .A(n_307), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g371 ( .A(n_307), .B(n_372), .Y(n_371) );
OAI21xp33_ASAP7_75t_L g374 ( .A1(n_309), .A2(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_313), .A2(n_322), .B1(n_325), .B2(n_326), .C(n_328), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_313), .B(n_347), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_313), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g429 ( .A(n_319), .Y(n_429) );
INVxp67_ASAP7_75t_L g352 ( .A(n_320), .Y(n_352) );
INVx1_ASAP7_75t_L g359 ( .A(n_322), .Y(n_359) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g398 ( .A(n_323), .B(n_327), .Y(n_398) );
INVx1_ASAP7_75t_L g372 ( .A(n_327), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_327), .B(n_342), .Y(n_402) );
OAI32xp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .A3(n_333), .B1(n_334), .B2(n_335), .Y(n_328) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_SL g341 ( .A(n_336), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_336), .B(n_368), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_336), .B(n_397), .Y(n_428) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_336), .B(n_347), .Y(n_436) );
NAND5xp2_ASAP7_75t_L g337 ( .A(n_338), .B(n_360), .C(n_373), .D(n_385), .E(n_386), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B1(n_343), .B2(n_345), .C(n_349), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp33_ASAP7_75t_SL g364 ( .A(n_344), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_347), .B(n_416), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_348), .A2(n_361), .B1(n_364), .B2(n_368), .Y(n_360) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
OAI211xp5_ASAP7_75t_SL g355 ( .A1(n_351), .A2(n_356), .B(n_357), .C(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g383 ( .A(n_363), .Y(n_383) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_372), .B(n_421), .Y(n_431) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI222xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B1(n_391), .B2(n_395), .C1(n_398), .C2(n_399), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_405), .B2(n_407), .C(n_409), .Y(n_401) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B(n_414), .Y(n_409) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g421 ( .A(n_413), .Y(n_421) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B1(n_422), .B2(n_424), .C(n_426), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_436), .B(n_437), .C(n_439), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g454 ( .A(n_446), .Y(n_454) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_451), .B(n_456), .C(n_745), .Y(n_455) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_732), .B1(n_735), .B2(n_736), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR4x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_621), .C(n_681), .D(n_708), .Y(n_459) );
NAND4xp25_ASAP7_75t_SL g460 ( .A(n_461), .B(n_569), .C(n_600), .D(n_617), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_504), .B(n_506), .C(n_549), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_485), .Y(n_462) );
INVx1_ASAP7_75t_L g611 ( .A(n_463), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_463), .A2(n_652), .B1(n_700), .B2(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_475), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_464), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g562 ( .A(n_464), .B(n_487), .Y(n_562) );
AND2x2_ASAP7_75t_L g604 ( .A(n_464), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_464), .B(n_505), .Y(n_616) );
INVx1_ASAP7_75t_L g656 ( .A(n_464), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_464), .B(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g584 ( .A(n_465), .B(n_487), .Y(n_584) );
INVx3_ASAP7_75t_L g588 ( .A(n_465), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_465), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g675 ( .A(n_475), .B(n_496), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_475), .B(n_588), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_475), .B(n_703), .Y(n_702) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g505 ( .A(n_476), .B(n_487), .Y(n_505) );
INVx1_ASAP7_75t_L g557 ( .A(n_476), .Y(n_557) );
BUFx2_ASAP7_75t_L g561 ( .A(n_476), .Y(n_561) );
AND2x2_ASAP7_75t_L g605 ( .A(n_476), .B(n_486), .Y(n_605) );
OR2x2_ASAP7_75t_L g644 ( .A(n_476), .B(n_486), .Y(n_644) );
AND2x2_ASAP7_75t_L g669 ( .A(n_476), .B(n_496), .Y(n_669) );
AND2x2_ASAP7_75t_L g728 ( .A(n_476), .B(n_558), .Y(n_728) );
INVx1_ASAP7_75t_L g703 ( .A(n_485), .Y(n_703) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_486), .B(n_496), .Y(n_589) );
AND2x2_ASAP7_75t_L g599 ( .A(n_486), .B(n_588), .Y(n_599) );
BUFx2_ASAP7_75t_L g610 ( .A(n_486), .Y(n_610) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g632 ( .A(n_487), .B(n_496), .Y(n_632) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_487), .Y(n_687) );
AND2x2_ASAP7_75t_SL g504 ( .A(n_496), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_SL g558 ( .A(n_496), .Y(n_558) );
BUFx2_ASAP7_75t_L g583 ( .A(n_496), .Y(n_583) );
INVx2_ASAP7_75t_L g602 ( .A(n_496), .Y(n_602) );
AND2x2_ASAP7_75t_L g664 ( .A(n_496), .B(n_588), .Y(n_664) );
AOI321xp33_ASAP7_75t_L g683 ( .A1(n_504), .A2(n_684), .A3(n_685), .B1(n_686), .B2(n_688), .C(n_689), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_505), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_505), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g677 ( .A(n_505), .B(n_656), .Y(n_677) );
AND2x2_ASAP7_75t_L g710 ( .A(n_505), .B(n_602), .Y(n_710) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_530), .Y(n_507) );
OR2x2_ASAP7_75t_L g612 ( .A(n_508), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g564 ( .A(n_511), .Y(n_564) );
AND2x2_ASAP7_75t_L g574 ( .A(n_511), .B(n_532), .Y(n_574) );
AND2x2_ASAP7_75t_L g579 ( .A(n_511), .B(n_554), .Y(n_579) );
INVx1_ASAP7_75t_L g596 ( .A(n_511), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_511), .B(n_577), .Y(n_615) );
AND2x2_ASAP7_75t_L g620 ( .A(n_511), .B(n_553), .Y(n_620) );
OR2x2_ASAP7_75t_L g652 ( .A(n_511), .B(n_641), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_511), .B(n_565), .Y(n_691) );
AND2x2_ASAP7_75t_L g725 ( .A(n_511), .B(n_551), .Y(n_725) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_518), .Y(n_511) );
INVx1_ASAP7_75t_L g552 ( .A(n_520), .Y(n_552) );
INVx2_ASAP7_75t_L g567 ( .A(n_520), .Y(n_567) );
AND2x2_ASAP7_75t_L g607 ( .A(n_520), .B(n_578), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_520), .B(n_554), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_526), .Y(n_523) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g713 ( .A(n_531), .B(n_564), .Y(n_713) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_541), .Y(n_531) );
INVx2_ASAP7_75t_L g554 ( .A(n_532), .Y(n_554) );
AND2x2_ASAP7_75t_L g707 ( .A(n_532), .B(n_567), .Y(n_707) );
AND2x2_ASAP7_75t_L g553 ( .A(n_541), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g568 ( .A(n_541), .Y(n_568) );
INVx1_ASAP7_75t_L g578 ( .A(n_541), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_555), .B1(n_559), .B2(n_563), .Y(n_549) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_550), .A2(n_668), .B1(n_705), .B2(n_706), .Y(n_704) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g619 ( .A(n_552), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_553), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g614 ( .A(n_554), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_554), .B(n_567), .Y(n_641) );
INVx1_ASAP7_75t_L g657 ( .A(n_554), .Y(n_657) );
AND2x2_ASAP7_75t_L g598 ( .A(n_556), .B(n_599), .Y(n_598) );
INVx3_ASAP7_75t_SL g637 ( .A(n_556), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_556), .B(n_562), .Y(n_714) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g723 ( .A(n_559), .Y(n_723) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_560), .B(n_656), .Y(n_698) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx3_ASAP7_75t_SL g603 ( .A(n_562), .Y(n_603) );
NAND2x1_ASAP7_75t_SL g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g624 ( .A(n_564), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g631 ( .A(n_564), .B(n_568), .Y(n_631) );
AND2x2_ASAP7_75t_L g636 ( .A(n_564), .B(n_577), .Y(n_636) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_564), .Y(n_685) );
OAI311xp33_ASAP7_75t_L g708 ( .A1(n_565), .A2(n_709), .A3(n_711), .B1(n_712), .C1(n_722), .Y(n_708) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g721 ( .A(n_566), .B(n_594), .Y(n_721) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
AND2x2_ASAP7_75t_L g577 ( .A(n_567), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g625 ( .A(n_567), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g680 ( .A(n_567), .Y(n_680) );
INVx1_ASAP7_75t_L g573 ( .A(n_568), .Y(n_573) );
INVx1_ASAP7_75t_L g593 ( .A(n_568), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_568), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g626 ( .A(n_568), .Y(n_626) );
AOI221xp5_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_572), .B1(n_580), .B2(n_585), .C(n_590), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_575), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx4_ASAP7_75t_L g594 ( .A(n_574), .Y(n_594) );
AND2x2_ASAP7_75t_L g688 ( .A(n_574), .B(n_607), .Y(n_688) );
AND2x2_ASAP7_75t_L g695 ( .A(n_574), .B(n_577), .Y(n_695) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_577), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g606 ( .A(n_579), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_582), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g731 ( .A(n_584), .B(n_675), .Y(n_731) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g716 ( .A(n_588), .B(n_644), .Y(n_716) );
OAI211xp5_ASAP7_75t_L g681 ( .A1(n_589), .A2(n_682), .B(n_683), .C(n_696), .Y(n_681) );
AOI21xp33_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_595), .B(n_597), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp67_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g660 ( .A(n_594), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g689 ( .A1(n_595), .A2(n_690), .B1(n_691), .B2(n_692), .C(n_693), .Y(n_689) );
AND2x2_ASAP7_75t_L g666 ( .A(n_596), .B(n_607), .Y(n_666) );
AND2x2_ASAP7_75t_L g719 ( .A(n_596), .B(n_614), .Y(n_719) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_599), .B(n_637), .Y(n_661) );
O2A1O1Ixp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_604), .B(n_606), .C(n_608), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g647 ( .A(n_602), .B(n_605), .Y(n_647) );
OR2x2_ASAP7_75t_L g690 ( .A(n_602), .B(n_644), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_603), .B(n_669), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_603), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g634 ( .A(n_604), .Y(n_634) );
INVx1_ASAP7_75t_L g700 ( .A(n_607), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .B1(n_615), .B2(n_616), .Y(n_608) );
INVx1_ASAP7_75t_L g623 ( .A(n_609), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_610), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g686 ( .A(n_611), .B(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g672 ( .A(n_613), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_614), .B(n_700), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_615), .A2(n_674), .B1(n_676), .B2(n_678), .Y(n_673) );
INVx1_ASAP7_75t_L g682 ( .A(n_618), .Y(n_682) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AND2x2_ASAP7_75t_L g724 ( .A(n_619), .B(n_719), .Y(n_724) );
AOI222xp33_ASAP7_75t_L g653 ( .A1(n_620), .A2(n_654), .B1(n_657), .B2(n_658), .C1(n_661), .C2(n_662), .Y(n_653) );
NAND4xp25_ASAP7_75t_SL g621 ( .A(n_622), .B(n_642), .C(n_653), .D(n_665), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_627), .B2(n_632), .C(n_633), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_625), .B(n_660), .Y(n_659) );
INVxp67_ASAP7_75t_L g651 ( .A(n_626), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_627), .A2(n_697), .B1(n_699), .B2(n_701), .C(n_704), .Y(n_696) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g639 ( .A(n_631), .B(n_640), .Y(n_639) );
OAI21xp33_ASAP7_75t_L g693 ( .A1(n_632), .A2(n_694), .B(n_695), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B1(n_637), .B2(n_638), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI21xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B(n_648), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g684 ( .A(n_655), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_656), .B(n_675), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_656), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_660), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g692 ( .A(n_664), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_670), .B2(n_672), .C(n_673), .Y(n_665) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g712 ( .A1(n_675), .A2(n_713), .B1(n_714), .B2(n_715), .C1(n_717), .C2(n_720), .Y(n_712) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_679), .B(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g711 ( .A(n_685), .Y(n_711) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVxp33_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_725), .B2(n_726), .C(n_729), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g742 ( .A(n_736), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_737), .Y(n_743) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
endmodule