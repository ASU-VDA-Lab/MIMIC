module fake_jpeg_31734_n_112 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_112);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_20),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_19),
.Y(n_37)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_8),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_2),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_18),
.B1(n_19),
.B2(n_15),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_39),
.A2(n_27),
.B1(n_28),
.B2(n_9),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_15),
.B1(n_22),
.B2(n_21),
.Y(n_42)
);

OA21x2_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_46),
.B(n_52),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_22),
.B1(n_21),
.B2(n_12),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_45),
.B1(n_52),
.B2(n_29),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_23),
.B1(n_17),
.B2(n_14),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_26),
.A2(n_23),
.B1(n_17),
.B2(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_5),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_48),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_43),
.B1(n_56),
.B2(n_66),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_32),
.B1(n_36),
.B2(n_28),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_67),
.B1(n_69),
.B2(n_59),
.Y(n_81)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_59),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_34),
.B(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_9),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_2),
.Y(n_66)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_62),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_34),
.B1(n_27),
.B2(n_11),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_73),
.B(n_69),
.C(n_57),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_43),
.B1(n_50),
.B2(n_11),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_53),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_67),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_84),
.B1(n_86),
.B2(n_69),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_87),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_57),
.B(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_89),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_69),
.B(n_65),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_96),
.B1(n_84),
.B2(n_76),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_75),
.C(n_74),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_75),
.C(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_99),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_84),
.B(n_71),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_55),
.B(n_77),
.Y(n_105)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_98),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_103),
.B(n_105),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_93),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_100),
.B1(n_97),
.B2(n_58),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_72),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_109),
.B(n_80),
.C(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_80),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_68),
.C(n_72),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_72),
.Y(n_112)
);


endmodule