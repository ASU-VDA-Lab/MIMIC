module fake_jpeg_3287_n_657 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_657);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_657;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_19),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_58),
.Y(n_161)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_59),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_60),
.Y(n_175)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_63),
.B(n_123),
.Y(n_225)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_64),
.Y(n_220)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

CKINVDCx9p33_ASAP7_75t_R g179 ( 
.A(n_65),
.Y(n_179)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_67),
.B(n_80),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_68),
.B(n_128),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_70),
.Y(n_197)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_71),
.Y(n_183)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_72),
.B(n_73),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_74),
.Y(n_189)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_75),
.Y(n_230)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_76),
.Y(n_188)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_78),
.Y(n_185)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_79),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_2),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_22),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_89),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_21),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_82),
.A2(n_100),
.B1(n_57),
.B2(n_56),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_24),
.B(n_3),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_83),
.B(n_84),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_24),
.B(n_4),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_85),
.Y(n_224)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_86),
.B(n_88),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_4),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_91),
.Y(n_209)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_92),
.B(n_96),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_94),
.Y(n_234)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_97),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_98),
.Y(n_169)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_99),
.B(n_101),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_27),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_104),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_28),
.Y(n_111)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_30),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g168 ( 
.A(n_112),
.B(n_131),
.Y(n_168)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_40),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_113),
.B(n_115),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_28),
.Y(n_114)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_38),
.B(n_6),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_117),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_43),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_30),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_121),
.B(n_124),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g122 ( 
.A(n_35),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g233 ( 
.A(n_122),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_37),
.B(n_6),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_125),
.Y(n_215)
);

BUFx8_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

BUFx16f_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_22),
.B(n_8),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_37),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_130),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_37),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_44),
.Y(n_132)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_132),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_135),
.A2(n_165),
.B1(n_208),
.B2(n_226),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_63),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_136),
.B(n_182),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_46),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_140),
.B(n_160),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_65),
.A2(n_33),
.B1(n_55),
.B2(n_50),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_145),
.A2(n_151),
.B1(n_171),
.B2(n_178),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_73),
.B(n_46),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_146),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_57),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_147),
.B(n_149),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_56),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_82),
.A2(n_53),
.B1(n_44),
.B2(n_55),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_60),
.B(n_51),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_155),
.B(n_172),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_32),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_61),
.A2(n_53),
.B1(n_44),
.B2(n_45),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_69),
.B(n_50),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_166),
.B(n_170),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_74),
.B(n_50),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_65),
.A2(n_55),
.B1(n_48),
.B2(n_36),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_94),
.B(n_39),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_87),
.A2(n_39),
.B1(n_51),
.B2(n_45),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_173),
.A2(n_223),
.B1(n_200),
.B2(n_201),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_23),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_174),
.B(n_177),
.Y(n_246)
);

HAxp5_ASAP7_75t_SL g176 ( 
.A(n_126),
.B(n_23),
.CON(n_176),
.SN(n_176)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_176),
.A2(n_66),
.B(n_168),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_48),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_126),
.A2(n_48),
.B1(n_36),
.B2(n_33),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_95),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_62),
.B(n_36),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_184),
.B(n_190),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_71),
.B(n_33),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_76),
.B(n_32),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_192),
.B(n_202),
.Y(n_268)
);

AO22x1_ASAP7_75t_SL g194 ( 
.A1(n_90),
.A2(n_53),
.B1(n_32),
.B2(n_11),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_194),
.B(n_228),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_130),
.A2(n_53),
.B1(n_10),
.B2(n_11),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_196),
.A2(n_161),
.B1(n_220),
.B2(n_197),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_93),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_200),
.A2(n_201),
.B1(n_161),
.B2(n_231),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_102),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_78),
.B(n_13),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_108),
.B(n_13),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_203),
.B(n_232),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_103),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_208),
.A2(n_226),
.B1(n_215),
.B2(n_187),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_105),
.B(n_14),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_210),
.B(n_213),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_109),
.B(n_14),
.C(n_16),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_212),
.B(n_169),
.C(n_207),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_110),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_111),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_218),
.B(n_227),
.Y(n_287)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_120),
.Y(n_221)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_114),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_118),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_125),
.B(n_17),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_97),
.B(n_66),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_59),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_231),
.B(n_216),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_127),
.B(n_122),
.Y(n_232)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_235),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_236),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_166),
.A2(n_170),
.B1(n_151),
.B2(n_194),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_238),
.A2(n_244),
.B1(n_259),
.B2(n_270),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_233),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_239),
.B(n_247),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_240),
.Y(n_340)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_137),
.Y(n_245)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_245),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_205),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_160),
.B(n_228),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_248),
.B(n_256),
.C(n_261),
.Y(n_337)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_249),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_250),
.B(n_278),
.Y(n_342)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_252),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_140),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_253),
.B(n_262),
.Y(n_330)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_254),
.Y(n_352)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_255),
.Y(n_358)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_214),
.B(n_148),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_168),
.A2(n_176),
.B(n_146),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_257),
.A2(n_211),
.B(n_150),
.Y(n_329)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_137),
.Y(n_258)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_258),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_165),
.A2(n_151),
.B1(n_136),
.B2(n_194),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_156),
.Y(n_260)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_260),
.Y(n_360)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_148),
.B(n_159),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_159),
.B(n_186),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_263),
.A2(n_284),
.B1(n_288),
.B2(n_301),
.Y(n_325)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_183),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_167),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_265),
.Y(n_348)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_156),
.Y(n_266)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_266),
.Y(n_369)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_183),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_267),
.Y(n_334)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_179),
.Y(n_269)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_269),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_151),
.A2(n_225),
.B1(n_182),
.B2(n_143),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_167),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_271),
.B(n_290),
.Y(n_385)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_167),
.Y(n_272)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_272),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_229),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_273),
.B(n_285),
.Y(n_363)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_209),
.Y(n_275)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_275),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_157),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_159),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_229),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_280),
.B(n_289),
.Y(n_349)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_157),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_281),
.Y(n_365)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_158),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_283),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_206),
.A2(n_225),
.B1(n_222),
.B2(n_139),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_220),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_220),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_286),
.B(n_291),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_L g288 ( 
.A1(n_213),
.A2(n_218),
.B1(n_163),
.B2(n_215),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_186),
.Y(n_289)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_158),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_163),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_292),
.B(n_294),
.Y(n_367)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_187),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_162),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_295),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_138),
.A2(n_204),
.B(n_212),
.C(n_186),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_296),
.A2(n_255),
.B(n_249),
.C(n_252),
.Y(n_376)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_188),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_298),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_209),
.Y(n_298)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_188),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_300),
.B(n_318),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_148),
.B(n_197),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_302),
.B(n_304),
.C(n_322),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_133),
.B(n_234),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_305),
.B(n_314),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_311),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_144),
.A2(n_195),
.B1(n_193),
.B2(n_154),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_133),
.A2(n_224),
.B1(n_199),
.B2(n_142),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_230),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_312),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_142),
.A2(n_195),
.B1(n_144),
.B2(n_193),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_230),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_154),
.A2(n_191),
.B1(n_189),
.B2(n_162),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_313),
.A2(n_317),
.B1(n_152),
.B2(n_134),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_141),
.B(n_199),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_153),
.A2(n_198),
.B1(n_224),
.B2(n_234),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_L g378 ( 
.A1(n_315),
.A2(n_240),
.B1(n_269),
.B2(n_273),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_141),
.B(n_150),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_319),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_L g317 ( 
.A1(n_189),
.A2(n_191),
.B1(n_217),
.B2(n_221),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_153),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_150),
.B(n_217),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_198),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_321),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_150),
.B(n_175),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_175),
.B(n_211),
.C(n_185),
.Y(n_322)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_164),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_323),
.B(n_240),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_329),
.B(n_368),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_L g397 ( 
.A1(n_338),
.A2(n_285),
.B1(n_260),
.B2(n_281),
.Y(n_397)
);

AOI32xp33_ASAP7_75t_L g344 ( 
.A1(n_303),
.A2(n_181),
.A3(n_134),
.B1(n_180),
.B2(n_164),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_344),
.A2(n_356),
.B(n_379),
.C(n_337),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_248),
.B(n_185),
.C(n_181),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_346),
.B(n_361),
.C(n_258),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_180),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_351),
.B(n_355),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_299),
.B(n_152),
.Y(n_355)
);

AOI32xp33_ASAP7_75t_L g356 ( 
.A1(n_309),
.A2(n_181),
.A3(n_299),
.B1(n_268),
.B2(n_282),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_248),
.B(n_251),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_380),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_253),
.C(n_256),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_244),
.A2(n_309),
.B1(n_259),
.B2(n_301),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_362),
.A2(n_294),
.B1(n_283),
.B2(n_266),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_257),
.A2(n_293),
.B(n_274),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_270),
.A2(n_287),
.B1(n_279),
.B2(n_256),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_373),
.A2(n_383),
.B1(n_311),
.B2(n_323),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_374),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_376),
.B(n_288),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_242),
.A2(n_237),
.B1(n_246),
.B2(n_319),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_377),
.A2(n_373),
.B1(n_330),
.B2(n_385),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_378),
.A2(n_286),
.B1(n_265),
.B2(n_272),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_241),
.A2(n_296),
.B(n_253),
.Y(n_379)
);

OAI32xp33_ASAP7_75t_L g380 ( 
.A1(n_262),
.A2(n_261),
.A3(n_302),
.B1(n_316),
.B2(n_322),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_320),
.B(n_312),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_381),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_261),
.A2(n_262),
.B1(n_302),
.B2(n_277),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_243),
.B(n_292),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_267),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_359),
.B(n_318),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_386),
.B(n_395),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_356),
.B(n_235),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_387),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_389),
.A2(n_397),
.B1(n_340),
.B2(n_382),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_390),
.A2(n_365),
.B(n_353),
.Y(n_475)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_391),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_367),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_413),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_379),
.B(n_254),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_327),
.B(n_310),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_396),
.B(n_412),
.Y(n_448)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_398),
.Y(n_462)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_399),
.Y(n_467)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_243),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g457 ( 
.A(n_403),
.B(n_411),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_331),
.A2(n_317),
.B1(n_291),
.B2(n_285),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_404),
.A2(n_340),
.B1(n_370),
.B2(n_366),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_405),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_345),
.B(n_245),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_406),
.B(n_409),
.Y(n_439)
);

NOR2x1_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_297),
.Y(n_407)
);

NOR2x1_ASAP7_75t_L g446 ( 
.A(n_407),
.B(n_363),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_348),
.Y(n_408)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_345),
.B(n_264),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_423),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_367),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_343),
.B(n_298),
.C(n_300),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_414),
.B(n_417),
.Y(n_469)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_347),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_415),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_362),
.A2(n_275),
.B1(n_295),
.B2(n_325),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_416),
.A2(n_335),
.B1(n_338),
.B2(n_329),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_418),
.B(n_425),
.Y(n_471)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_419),
.Y(n_472)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_347),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_422),
.Y(n_438)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_341),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_421),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_367),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_339),
.B(n_355),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_364),
.B(n_342),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_427),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_343),
.B(n_337),
.Y(n_425)
);

BUFx5_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

INVx13_ASAP7_75t_L g463 ( 
.A(n_426),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_363),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_339),
.B(n_351),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_429),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_330),
.B(n_376),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_333),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_431),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_363),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_350),
.B(n_354),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_433),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_350),
.B(n_354),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_434),
.A2(n_444),
.B1(n_447),
.B2(n_453),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_416),
.A2(n_325),
.B1(n_335),
.B2(n_330),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_437),
.A2(n_445),
.B1(n_450),
.B2(n_418),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_406),
.Y(n_441)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_441),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_393),
.A2(n_380),
.B1(n_358),
.B2(n_336),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_446),
.A2(n_460),
.B(n_475),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_393),
.A2(n_358),
.B1(n_336),
.B2(n_344),
.Y(n_450)
);

INVxp67_ASAP7_75t_R g451 ( 
.A(n_392),
.Y(n_451)
);

FAx1_ASAP7_75t_L g513 ( 
.A(n_451),
.B(n_426),
.CI(n_341),
.CON(n_513),
.SN(n_513)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_389),
.A2(n_383),
.B1(n_346),
.B2(n_349),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_402),
.B(n_357),
.Y(n_456)
);

CKINVDCx14_ASAP7_75t_R g484 ( 
.A(n_456),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_409),
.Y(n_459)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_459),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_388),
.A2(n_332),
.B(n_324),
.Y(n_460)
);

OAI32xp33_ASAP7_75t_L g465 ( 
.A1(n_394),
.A2(n_333),
.A3(n_365),
.B1(n_382),
.B2(n_353),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_468),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_410),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g501 ( 
.A(n_466),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_396),
.B(n_401),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_432),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_474),
.B(n_422),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_443),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_476),
.B(n_486),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_425),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_477),
.B(n_487),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_411),
.C(n_403),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_478),
.B(n_488),
.C(n_492),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_449),
.Y(n_480)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_480),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_481),
.A2(n_506),
.B1(n_453),
.B2(n_472),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_401),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_483),
.B(n_494),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_438),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_485),
.B(n_496),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_473),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_471),
.B(n_394),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_423),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_473),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_489),
.B(n_504),
.Y(n_528)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_491),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_465),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_414),
.C(n_428),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_493),
.B(n_495),
.C(n_499),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_386),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_464),
.B(n_417),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_442),
.B(n_419),
.Y(n_496)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_454),
.Y(n_498)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_498),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_445),
.B(n_429),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_454),
.Y(n_500)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_500),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_440),
.B(n_388),
.C(n_430),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_502),
.B(n_507),
.Y(n_535)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_462),
.Y(n_503)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_503),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_438),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_413),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_505),
.B(n_512),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_472),
.A2(n_412),
.B1(n_390),
.B2(n_395),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_456),
.B(n_372),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_448),
.A2(n_388),
.B1(n_407),
.B2(n_431),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_508),
.A2(n_510),
.B1(n_466),
.B2(n_491),
.Y(n_521)
);

OAI22xp33_ASAP7_75t_SL g509 ( 
.A1(n_441),
.A2(n_407),
.B1(n_433),
.B2(n_391),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_509),
.A2(n_459),
.B1(n_436),
.B2(n_450),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_448),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_435),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_511),
.B(n_455),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_435),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_SL g539 ( 
.A1(n_513),
.A2(n_508),
.B(n_479),
.C(n_510),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_517),
.A2(n_521),
.B1(n_523),
.B2(n_532),
.Y(n_561)
);

NOR2x1_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_464),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_518),
.B(n_526),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_479),
.Y(n_520)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_520),
.Y(n_559)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_498),
.Y(n_524)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_524),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_514),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_525),
.B(n_531),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_514),
.A2(n_446),
.B(n_460),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_490),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_530),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_513),
.B(n_475),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_482),
.A2(n_437),
.B1(n_444),
.B2(n_452),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_513),
.A2(n_446),
.B(n_461),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_533),
.B(n_539),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_501),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_534),
.B(n_537),
.Y(n_571)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_490),
.Y(n_536)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_536),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_505),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_481),
.A2(n_451),
.B1(n_452),
.B2(n_447),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_541),
.A2(n_548),
.B1(n_420),
.B2(n_415),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_484),
.A2(n_461),
.B1(n_451),
.B2(n_439),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_542),
.A2(n_470),
.B1(n_467),
.B2(n_462),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_486),
.B(n_455),
.Y(n_546)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_546),
.Y(n_578)
);

CKINVDCx14_ASAP7_75t_R g555 ( 
.A(n_547),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_512),
.A2(n_436),
.B1(n_461),
.B2(n_439),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_538),
.B(n_493),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_551),
.B(n_528),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_532),
.A2(n_489),
.B1(n_504),
.B2(n_497),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_552),
.A2(n_565),
.B1(n_568),
.B2(n_577),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_538),
.B(n_477),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_553),
.B(n_556),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_478),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_540),
.B(n_527),
.C(n_492),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_558),
.B(n_567),
.C(n_570),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_546),
.B(n_476),
.Y(n_562)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_562),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_527),
.B(n_488),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_563),
.B(n_564),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_518),
.B(n_495),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_517),
.A2(n_497),
.B1(n_499),
.B2(n_487),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_535),
.B(n_503),
.C(n_500),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_529),
.A2(n_467),
.B1(n_470),
.B2(n_458),
.Y(n_569)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_569),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_525),
.B(n_375),
.C(n_372),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_515),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_572),
.B(n_545),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_526),
.B(n_375),
.C(n_334),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_573),
.B(n_576),
.C(n_531),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_575),
.A2(n_533),
.B1(n_515),
.B2(n_516),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_541),
.B(n_326),
.C(n_334),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_521),
.A2(n_458),
.B1(n_408),
.B2(n_366),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_581),
.Y(n_609)
);

OAI321xp33_ASAP7_75t_L g618 ( 
.A1(n_582),
.A2(n_597),
.A3(n_598),
.B1(n_600),
.B2(n_583),
.C(n_602),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_555),
.B(n_519),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_584),
.B(n_585),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_575),
.A2(n_578),
.B1(n_516),
.B2(n_561),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_586),
.A2(n_587),
.B1(n_602),
.B2(n_549),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_578),
.A2(n_528),
.B1(n_545),
.B2(n_539),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_588),
.B(n_566),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_550),
.A2(n_539),
.B(n_531),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_589),
.A2(n_599),
.B(n_577),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_571),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_590),
.B(n_593),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_551),
.B(n_567),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_591),
.B(n_595),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_559),
.A2(n_539),
.B1(n_548),
.B2(n_531),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_558),
.B(n_522),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_556),
.B(n_536),
.C(n_524),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_596),
.B(n_570),
.C(n_573),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_566),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_552),
.B(n_530),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_550),
.A2(n_544),
.B(n_543),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_562),
.B(n_549),
.Y(n_600)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_560),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_603),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_580),
.B(n_596),
.C(n_579),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_604),
.B(n_606),
.Y(n_624)
);

FAx1_ASAP7_75t_SL g605 ( 
.A(n_589),
.B(n_565),
.CI(n_574),
.CON(n_605),
.SN(n_605)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_605),
.B(n_615),
.Y(n_622)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_600),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_580),
.B(n_553),
.C(n_563),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_607),
.B(n_612),
.Y(n_633)
);

BUFx24_ASAP7_75t_SL g611 ( 
.A(n_590),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g634 ( 
.A(n_611),
.B(n_613),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_579),
.B(n_564),
.C(n_576),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_585),
.B(n_559),
.C(n_554),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_601),
.A2(n_554),
.B1(n_560),
.B2(n_557),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_SL g632 ( 
.A1(n_614),
.A2(n_619),
.B1(n_621),
.B2(n_597),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_616),
.B(n_593),
.Y(n_626)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_617),
.Y(n_623)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g631 ( 
.A1(n_618),
.A2(n_599),
.B(n_587),
.C(n_581),
.D(n_586),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_592),
.B(n_408),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_592),
.B(n_544),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_608),
.A2(n_601),
.B1(n_583),
.B2(n_598),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_625),
.A2(n_630),
.B1(n_631),
.B2(n_463),
.Y(n_643)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_626),
.B(n_628),
.Y(n_639)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_603),
.B(n_594),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g629 ( 
.A(n_612),
.B(n_594),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_629),
.B(n_632),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_615),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_634),
.B(n_610),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_635),
.B(n_640),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_622),
.A2(n_608),
.B(n_609),
.Y(n_636)
);

AOI31xp33_ASAP7_75t_L g644 ( 
.A1(n_636),
.A2(n_630),
.A3(n_623),
.B(n_638),
.Y(n_644)
);

AOI322xp5_ASAP7_75t_L g637 ( 
.A1(n_623),
.A2(n_620),
.A3(n_614),
.B1(n_605),
.B2(n_543),
.C1(n_613),
.C2(n_588),
.Y(n_637)
);

OAI221xp5_ASAP7_75t_L g649 ( 
.A1(n_637),
.A2(n_622),
.B1(n_625),
.B2(n_626),
.C(n_463),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_627),
.B(n_604),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_624),
.A2(n_605),
.B(n_607),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_641),
.B(n_642),
.C(n_629),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_628),
.B(n_326),
.C(n_371),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_643),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_644),
.A2(n_648),
.B(n_649),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_647),
.B(n_639),
.C(n_642),
.Y(n_652)
);

NOR2x1_ASAP7_75t_L g648 ( 
.A(n_636),
.B(n_633),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_646),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_651),
.B(n_652),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_650),
.B(n_639),
.C(n_645),
.Y(n_654)
);

AOI322xp5_ASAP7_75t_L g655 ( 
.A1(n_654),
.A2(n_644),
.A3(n_643),
.B1(n_463),
.B2(n_348),
.C1(n_370),
.C2(n_421),
.Y(n_655)
);

OAI321xp33_ASAP7_75t_L g656 ( 
.A1(n_655),
.A2(n_348),
.A3(n_352),
.B1(n_371),
.B2(n_653),
.C(n_557),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_656),
.Y(n_657)
);


endmodule