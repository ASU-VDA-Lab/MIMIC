module real_jpeg_4220_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_1),
.A2(n_83),
.B1(n_84),
.B2(n_88),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_1),
.A2(n_83),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_1),
.A2(n_66),
.B1(n_83),
.B2(n_335),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_1),
.A2(n_45),
.B1(n_83),
.B2(n_319),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_2),
.A2(n_86),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_2),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_2),
.A2(n_193),
.B1(n_258),
.B2(n_263),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_2),
.A2(n_162),
.B1(n_193),
.B2(n_318),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g417 ( 
.A1(n_2),
.A2(n_149),
.B1(n_193),
.B2(n_418),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_3),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_4),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_4),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_4),
.A2(n_258),
.B1(n_276),
.B2(n_294),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_4),
.A2(n_126),
.B1(n_276),
.B2(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_4),
.A2(n_192),
.B1(n_276),
.B2(n_412),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_5),
.A2(n_143),
.B1(n_148),
.B2(n_151),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_5),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_151),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_5),
.A2(n_151),
.B1(n_204),
.B2(n_208),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_5),
.A2(n_151),
.B1(n_294),
.B2(n_366),
.Y(n_365)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_6),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_7),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_7),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_8),
.A2(n_69),
.B1(n_70),
.B2(n_74),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_8),
.A2(n_38),
.B1(n_69),
.B2(n_170),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_8),
.A2(n_69),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_9),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_9),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_9),
.A2(n_102),
.B1(n_241),
.B2(n_244),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_9),
.A2(n_102),
.B1(n_170),
.B2(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_9),
.A2(n_95),
.B1(n_102),
.B2(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_48),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_10),
.A2(n_42),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_10),
.A2(n_42),
.B1(n_400),
.B2(n_402),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_11),
.A2(n_35),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_12),
.Y(n_384)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_12),
.Y(n_388)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_13),
.Y(n_89)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_13),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_13),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_13),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_13),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_13),
.Y(n_413)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_15),
.A2(n_164),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_15),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_15),
.B(n_251),
.C(n_254),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_15),
.B(n_134),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_15),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_15),
.B(n_77),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_15),
.B(n_326),
.Y(n_325)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_16),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_226),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_224),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_195),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_20),
.B(n_195),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_115),
.C(n_166),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_21),
.A2(n_22),
.B1(n_115),
.B2(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_78),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_23),
.A2(n_24),
.B(n_80),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_24),
.A2(n_79),
.B1(n_80),
.B2(n_114),
.Y(n_78)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_24),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_24),
.A2(n_40),
.B1(n_114),
.B2(n_429),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B(n_34),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_25),
.A2(n_34),
.B1(n_169),
.B2(n_173),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_25),
.A2(n_257),
.B(n_265),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_25),
.A2(n_238),
.B(n_265),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_25),
.A2(n_394),
.B1(n_395),
.B2(n_398),
.Y(n_393)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_26),
.B(n_268),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_26),
.A2(n_299),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_26),
.A2(n_334),
.B1(n_365),
.B2(n_367),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_26),
.A2(n_399),
.B1(n_435),
.B2(n_436),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_31),
.Y(n_174)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_33),
.Y(n_267)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_33),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_37),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_38),
.Y(n_287)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_39),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_40),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_51),
.B1(n_68),
.B2(n_77),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_41),
.A2(n_51),
.B1(n_77),
.B2(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_46),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_46),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_46),
.Y(n_245)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_47),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_47),
.Y(n_139)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_47),
.Y(n_182)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_47),
.Y(n_279)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_51),
.A2(n_68),
.B1(n_77),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_51),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_51),
.B(n_240),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_63),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_62),
.Y(n_178)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_63),
.A2(n_273),
.B(n_280),
.Y(n_272)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_73),
.Y(n_243)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_73),
.Y(n_249)
);

AOI32xp33_ASAP7_75t_L g340 ( 
.A1(n_74),
.A2(n_121),
.A3(n_325),
.B1(n_341),
.B2(n_344),
.Y(n_340)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_76),
.Y(n_237)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_77),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_77),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_100),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_90),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_82),
.Y(n_201)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_90),
.B(n_101),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_90),
.Y(n_202)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_98),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_94),
.Y(n_218)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_94),
.Y(n_330)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_100),
.A2(n_202),
.B(n_439),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_108),
.Y(n_100)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_106),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_106),
.B(n_238),
.Y(n_391)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_108),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_108),
.A2(n_410),
.B(n_414),
.Y(n_409)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_115),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_158),
.B(n_165),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_159),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_134),
.B1(n_141),
.B2(n_152),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_118),
.A2(n_323),
.B(n_327),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_118),
.B(n_361),
.Y(n_360)
);

AOI22x1_ASAP7_75t_L g440 ( 
.A1(n_118),
.A2(n_134),
.B1(n_361),
.B2(n_441),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_118),
.A2(n_327),
.B(n_457),
.Y(n_456)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_119),
.A2(n_142),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_119),
.A2(n_187),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_119),
.A2(n_187),
.B1(n_357),
.B2(n_417),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_134),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_126),
.B1(n_129),
.B2(n_131),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_126),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_130),
.Y(n_346)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_133),
.Y(n_221)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

AO22x2_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_SL g323 ( 
.A1(n_144),
.A2(n_238),
.B(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_147),
.Y(n_343)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_147),
.Y(n_359)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_147),
.Y(n_380)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_147),
.Y(n_390)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_161),
.A2(n_211),
.B(n_212),
.Y(n_210)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_166),
.B(n_443),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_183),
.C(n_188),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_167),
.B(n_427),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_168),
.B(n_175),
.Y(n_451)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_169),
.Y(n_435)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_171),
.Y(n_264)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_171),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_172),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_172),
.Y(n_297)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_176),
.Y(n_433)
);

NAND2xp33_ASAP7_75t_SL g344 ( 
.A(n_177),
.B(n_345),
.Y(n_344)
);

INVx4_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_181),
.Y(n_320)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_183),
.B(n_188),
.Y(n_427)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_184),
.Y(n_441)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_187),
.B(n_328),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_187),
.A2(n_357),
.B(n_360),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B(n_194),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_189),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_189),
.A2(n_190),
.B1(n_202),
.B2(n_439),
.Y(n_438)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_194),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_209),
.B2(n_223),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_202),
.B(n_238),
.Y(n_363)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_213),
.B1(n_214),
.B2(n_222),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_211),
.A2(n_235),
.B(n_239),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_211),
.A2(n_212),
.B1(n_273),
.B2(n_317),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_211),
.A2(n_239),
.B(n_317),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_211),
.A2(n_212),
.B1(n_420),
.B2(n_433),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_212),
.A2(n_280),
.B(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_217),
.Y(n_418)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI311xp33_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_423),
.A3(n_459),
.B1(n_477),
.C1(n_478),
.Y(n_227)
);

AOI21x1_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_371),
.B(n_422),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_348),
.B(n_370),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_311),
.B(n_347),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_283),
.B(n_310),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_255),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_233),
.B(n_255),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_246),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_234),
.A2(n_246),
.B1(n_247),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_234),
.Y(n_308)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

OAI21xp33_ASAP7_75t_SL g410 ( 
.A1(n_238),
.A2(n_391),
.B(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_270),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_271),
.C(n_282),
.Y(n_312)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_262),
.Y(n_337)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_281),
.B2(n_282),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_303),
.B(n_309),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_291),
.B(n_302),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_290),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_289),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_301),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_301),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_298),
.B(n_300),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_296),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_300),
.A2(n_333),
.B(n_338),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_307),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_313),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_331),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_321),
.B2(n_322),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_321),
.C(n_331),
.Y(n_349)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx5_ASAP7_75t_SL g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_328),
.Y(n_361)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_340),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_340),
.Y(n_354)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_SL g338 ( 
.A(n_339),
.Y(n_338)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_349),
.B(n_350),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_355),
.B2(n_369),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_354),
.C(n_369),
.Y(n_372)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_355),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_362),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_356),
.B(n_363),
.C(n_364),
.Y(n_404)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_365),
.Y(n_394)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_372),
.B(n_373),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_407),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_404),
.B1(n_405),
.B2(n_406),
.Y(n_374)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_392),
.B2(n_393),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_377),
.B(n_392),
.Y(n_455)
);

OAI32xp33_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_381),
.A3(n_383),
.B1(n_385),
.B2(n_391),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_389),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_397),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_404),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_404),
.B(n_405),
.C(n_407),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_409),
.B1(n_415),
.B2(n_421),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_408),
.B(n_416),
.C(n_419),
.Y(n_468)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_415),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_419),
.Y(n_415)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_417),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_445),
.Y(n_423)
);

A2O1A1Ixp33_ASAP7_75t_SL g478 ( 
.A1(n_424),
.A2(n_445),
.B(n_479),
.C(n_482),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_442),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_425),
.B(n_442),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.C(n_430),
.Y(n_425)
);

FAx1_ASAP7_75t_SL g458 ( 
.A(n_426),
.B(n_428),
.CI(n_430),
.CON(n_458),
.SN(n_458)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_437),
.C(n_440),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_449),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_432),
.B(n_434),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_437),
.A2(n_438),
.B1(n_440),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_440),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_458),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_458),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_451),
.C(n_452),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_447),
.A2(n_448),
.B1(n_451),
.B2(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_451),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_470),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.C(n_456),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_453),
.A2(n_454),
.B1(n_456),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_456),
.Y(n_465)
);

BUFx24_ASAP7_75t_SL g483 ( 
.A(n_458),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_472),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_461),
.A2(n_480),
.B(n_481),
.Y(n_479)
);

NOR2x1_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_469),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_469),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.C(n_468),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_475),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_466),
.A2(n_467),
.B1(n_468),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_468),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_474),
.Y(n_480)
);


endmodule