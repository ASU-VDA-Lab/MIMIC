module fake_jpeg_21358_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_14),
.B1(n_17),
.B2(n_15),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_30),
.B1(n_26),
.B2(n_16),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_13),
.B1(n_16),
.B2(n_12),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

AND2x6_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_24),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_21),
.B(n_35),
.C(n_29),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_35),
.B(n_12),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_30),
.B1(n_34),
.B2(n_31),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_20),
.B(n_11),
.Y(n_55)
);

OAI22x1_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_40),
.B1(n_44),
.B2(n_43),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_51),
.B1(n_42),
.B2(n_31),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_22),
.C(n_10),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_19),
.C(n_11),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_10),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_50),
.B(n_49),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_2),
.B(n_3),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_57),
.B1(n_11),
.B2(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_46),
.Y(n_64)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_66),
.A3(n_67),
.B1(n_8),
.B2(n_2),
.C1(n_63),
.C2(n_19),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

AOI322xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_20),
.A3(n_19),
.B1(n_7),
.B2(n_6),
.C1(n_8),
.C2(n_4),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_2),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_70),
.B(n_71),
.Y(n_72)
);


endmodule