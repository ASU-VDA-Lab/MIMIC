module real_jpeg_3473_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_1),
.A2(n_52),
.B1(n_54),
.B2(n_58),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_58),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_1),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_331)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_44),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_3),
.A2(n_44),
.B1(n_63),
.B2(n_64),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_3),
.A2(n_44),
.B1(n_52),
.B2(n_54),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_4),
.B(n_63),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_4),
.B(n_165),
.Y(n_202)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_4),
.A2(n_29),
.B(n_30),
.C(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_4),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_4),
.B(n_35),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_215),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_4),
.B(n_49),
.C(n_52),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_215),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_4),
.B(n_92),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_4),
.B(n_81),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_5),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_124),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_124),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_5),
.A2(n_52),
.B1(n_54),
.B2(n_124),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_66),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_66),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_7),
.A2(n_52),
.B1(n_54),
.B2(n_66),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_56),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_8),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_8),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_10),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_164),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_164),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_10),
.A2(n_52),
.B1(n_54),
.B2(n_164),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_102),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_102),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_14),
.A2(n_52),
.B1(n_54),
.B2(n_102),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_15),
.A2(n_41),
.B1(n_63),
.B2(n_64),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_15),
.A2(n_41),
.B1(n_52),
.B2(n_54),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_328),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_315),
.B(n_327),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_140),
.B(n_312),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_127),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_103),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_23),
.B(n_103),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_84),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_59),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_25),
.A2(n_26),
.B(n_45),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_25),
.B(n_59),
.C(n_84),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_45),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_27),
.A2(n_42),
.B1(n_43),
.B2(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_27),
.A2(n_40),
.B1(n_42),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_27),
.A2(n_42),
.B1(n_78),
.B2(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_27),
.A2(n_181),
.B(n_183),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_27),
.A2(n_183),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_28),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_28),
.A2(n_35),
.B1(n_182),
.B2(n_199),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_28),
.A2(n_35),
.B(n_319),
.Y(n_318)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B(n_34),
.C(n_35),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

AO22x2_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_35)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_30),
.A2(n_31),
.B1(n_70),
.B2(n_72),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g185 ( 
.A1(n_30),
.A2(n_64),
.A3(n_70),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_31),
.B(n_72),
.Y(n_187)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_35),
.B(n_161),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_37),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_36),
.A2(n_39),
.B(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_37),
.B(n_260),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_42),
.A2(n_120),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_42),
.A2(n_160),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_51),
.B1(n_55),
.B2(n_57),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_46),
.A2(n_51),
.B1(n_55),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_46),
.A2(n_51),
.B1(n_208),
.B2(n_242),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_46),
.A2(n_210),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_47),
.A2(n_81),
.B1(n_97),
.B2(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_47),
.A2(n_81),
.B1(n_118),
.B2(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_47),
.A2(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_47),
.B(n_211),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_51),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_51),
.A2(n_231),
.B(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_52),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_52),
.B(n_271),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_75),
.B2(n_83),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_60),
.A2(n_61),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_SL g138 ( 
.A(n_61),
.B(n_76),
.C(n_80),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_61),
.B(n_131),
.C(n_138),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_69),
.B2(n_74),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_69),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_64),
.B1(n_70),
.B2(n_72),
.Y(n_73)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_64),
.A2(n_67),
.B(n_215),
.C(n_224),
.Y(n_223)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_67),
.A2(n_122),
.B(n_125),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_67),
.A2(n_69),
.B1(n_74),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_68),
.A2(n_123),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_68),
.A2(n_165),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_68),
.A2(n_165),
.B1(n_322),
.B2(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_69),
.A2(n_99),
.B(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_70),
.Y(n_72)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_79),
.A2(n_80),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_80),
.B(n_132),
.C(n_136),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_81),
.B(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_88),
.B(n_98),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_86),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_95),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_88),
.B1(n_98),
.B2(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_87),
.A2(n_88),
.B1(n_95),
.B2(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_92),
.B(n_93),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_89),
.A2(n_92),
.B1(n_115),
.B2(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_89),
.A2(n_215),
.B(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_90),
.A2(n_91),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_90),
.A2(n_91),
.B1(n_190),
.B2(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_90),
.B(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_90),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_90),
.A2(n_91),
.B1(n_246),
.B2(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_91),
.A2(n_205),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_91),
.B(n_219),
.Y(n_248)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_92),
.A2(n_218),
.B(n_275),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_95),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.C(n_110),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_105),
.B1(n_109),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_119),
.C(n_121),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_112),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_121),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_126),
.B(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_127),
.A2(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_139),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_128),
.B(n_139),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_138),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_133),
.Y(n_321)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_137),
.Y(n_319)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_166),
.B(n_311),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_142),
.B(n_145),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_158),
.C(n_162),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_153),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_154),
.B(n_156),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_192),
.B(n_310),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_168),
.B(n_170),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.C(n_177),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_171),
.B(n_175),
.Y(n_295)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_177),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_184),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_178),
.B(n_180),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_184),
.B(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_185),
.A2(n_188),
.B1(n_189),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI31xp33_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_292),
.A3(n_302),
.B(n_307),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_236),
.B(n_291),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_220),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_195),
.B(n_220),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_206),
.C(n_212),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_196),
.B(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_201),
.C(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_206),
.B(n_212),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_216),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_232),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_221),
.B(n_233),
.C(n_235),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_222),
.B(n_227),
.C(n_228),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_286),
.B(n_290),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_255),
.B(n_285),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_249),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_249),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.C(n_244),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_245),
.B1(n_264),
.B2(n_266),
.Y(n_263)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_253),
.C(n_254),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_267),
.B(n_284),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_263),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_263),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_278),
.B(n_283),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_273),
.B(n_277),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_276),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_275),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_281),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_289),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_296),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.C(n_300),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_306),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_326),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_326),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_325),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_320),
.B1(n_323),
.B2(n_324),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_323),
.C(n_325),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_333),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);


endmodule