module real_aes_8486_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_501, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_501;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_330;
wire n_388;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_434;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_288;
wire n_150;
wire n_147;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_484;
wire n_326;
wire n_492;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_SL g235 ( .A1(n_0), .A2(n_236), .B(n_237), .C(n_241), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_1), .B(n_230), .Y(n_243) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
AOI221xp5_ASAP7_75t_L g134 ( .A1(n_3), .A2(n_31), .B1(n_135), .B2(n_138), .C(n_141), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_4), .B(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_5), .A2(n_224), .B(n_326), .Y(n_325) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_6), .A2(n_197), .B(n_283), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g114 ( .A1(n_7), .A2(n_66), .B1(n_115), .B2(n_120), .C(n_124), .Y(n_114) );
INVx1_ASAP7_75t_L g142 ( .A(n_8), .Y(n_142) );
AOI221xp5_ASAP7_75t_L g81 ( .A1(n_9), .A2(n_22), .B1(n_82), .B2(n_99), .C(n_103), .Y(n_81) );
AOI222xp33_ASAP7_75t_L g153 ( .A1(n_10), .A2(n_17), .B1(n_70), .B2(n_154), .C1(n_156), .C2(n_160), .Y(n_153) );
INVx1_ASAP7_75t_L g187 ( .A(n_11), .Y(n_187) );
AND2x6_ASAP7_75t_L g222 ( .A(n_11), .B(n_185), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_11), .B(n_487), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g300 ( .A1(n_12), .A2(n_205), .B(n_222), .C(n_301), .Y(n_300) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_13), .A2(n_25), .B1(n_88), .B2(n_93), .Y(n_96) );
INVx1_ASAP7_75t_L g202 ( .A(n_14), .Y(n_202) );
OAI22xp5_ASAP7_75t_SL g171 ( .A1(n_15), .A2(n_72), .B1(n_172), .B2(n_173), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_15), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_16), .B(n_216), .Y(n_289) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_18), .A2(n_27), .B1(n_88), .B2(n_89), .Y(n_98) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_19), .A2(n_205), .B(n_267), .C(n_272), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_20), .A2(n_205), .B(n_272), .C(n_286), .Y(n_285) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_21), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_23), .A2(n_224), .B(n_232), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_23), .A2(n_80), .B1(n_165), .B2(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_23), .Y(n_483) );
INVx2_ASAP7_75t_L g207 ( .A(n_24), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_26), .A2(n_220), .B(n_251), .C(n_252), .Y(n_250) );
OAI221xp5_ASAP7_75t_L g178 ( .A1(n_27), .A2(n_43), .B1(n_54), .B2(n_179), .C(n_180), .Y(n_178) );
INVxp67_ASAP7_75t_L g181 ( .A(n_27), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_28), .B(n_288), .Y(n_287) );
OAI22xp5_ASAP7_75t_SL g167 ( .A1(n_29), .A2(n_58), .B1(n_168), .B2(n_169), .Y(n_167) );
INVx1_ASAP7_75t_L g169 ( .A(n_29), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_29), .B(n_265), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_30), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_32), .B(n_216), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_33), .B(n_224), .Y(n_284) );
INVx1_ASAP7_75t_L g147 ( .A(n_34), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_35), .A2(n_220), .B(n_251), .C(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g125 ( .A(n_36), .Y(n_125) );
INVx1_ASAP7_75t_L g238 ( .A(n_37), .Y(n_238) );
INVx1_ASAP7_75t_L g104 ( .A(n_38), .Y(n_104) );
INVx1_ASAP7_75t_L g313 ( .A(n_39), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_40), .B(n_224), .Y(n_310) );
INVx1_ASAP7_75t_L g129 ( .A(n_41), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_42), .Y(n_276) );
AO22x2_ASAP7_75t_L g87 ( .A1(n_43), .A2(n_62), .B1(n_88), .B2(n_89), .Y(n_87) );
INVxp67_ASAP7_75t_L g182 ( .A(n_43), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_44), .A2(n_80), .B1(n_165), .B2(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_44), .Y(n_495) );
INVx1_ASAP7_75t_L g185 ( .A(n_45), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_46), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_47), .B(n_230), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g328 ( .A1(n_48), .A2(n_212), .B(n_271), .C(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g201 ( .A(n_49), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_50), .A2(n_80), .B1(n_164), .B2(n_165), .Y(n_79) );
INVx1_ASAP7_75t_SL g164 ( .A(n_50), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_51), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_52), .B(n_216), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_53), .B(n_217), .Y(n_302) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_54), .A2(n_68), .B1(n_88), .B2(n_93), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g233 ( .A(n_55), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_56), .B(n_255), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_57), .A2(n_205), .B(n_210), .C(n_220), .Y(n_204) );
INVx1_ASAP7_75t_L g168 ( .A(n_58), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g327 ( .A(n_59), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_60), .B(n_254), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_61), .Y(n_260) );
INVx2_ASAP7_75t_L g199 ( .A(n_63), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_64), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_65), .B(n_240), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_67), .B(n_224), .Y(n_249) );
INVx1_ASAP7_75t_L g253 ( .A(n_69), .Y(n_253) );
INVxp67_ASAP7_75t_L g330 ( .A(n_71), .Y(n_330) );
INVx1_ASAP7_75t_L g173 ( .A(n_72), .Y(n_173) );
INVx1_ASAP7_75t_L g88 ( .A(n_73), .Y(n_88) );
INVx1_ASAP7_75t_L g90 ( .A(n_73), .Y(n_90) );
INVx1_ASAP7_75t_L g211 ( .A(n_74), .Y(n_211) );
INVx1_ASAP7_75t_L g298 ( .A(n_75), .Y(n_298) );
AND2x2_ASAP7_75t_L g315 ( .A(n_76), .B(n_258), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_175), .B1(n_188), .B2(n_480), .C(n_481), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_166), .Y(n_78) );
INVx1_ASAP7_75t_L g165 ( .A(n_80), .Y(n_165) );
AND4x1_ASAP7_75t_L g80 ( .A(n_81), .B(n_114), .C(n_134), .D(n_153), .Y(n_80) );
BUFx6f_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
BUFx6f_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
AND2x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_94), .Y(n_84) );
AND2x6_ASAP7_75t_L g117 ( .A(n_85), .B(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g123 ( .A(n_85), .B(n_107), .Y(n_123) );
AND2x6_ASAP7_75t_L g155 ( .A(n_85), .B(n_150), .Y(n_155) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_91), .Y(n_85) );
AND2x2_ASAP7_75t_L g102 ( .A(n_86), .B(n_92), .Y(n_102) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g108 ( .A(n_87), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_87), .B(n_92), .Y(n_113) );
AND2x2_ASAP7_75t_L g145 ( .A(n_87), .B(n_96), .Y(n_145) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g93 ( .A(n_90), .Y(n_93) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g109 ( .A(n_92), .Y(n_109) );
INVx1_ASAP7_75t_L g159 ( .A(n_92), .Y(n_159) );
AND2x4_ASAP7_75t_L g101 ( .A(n_94), .B(n_102), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_94), .B(n_108), .Y(n_128) );
AND2x4_ASAP7_75t_L g132 ( .A(n_94), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g94 ( .A(n_95), .B(n_97), .Y(n_94) );
AND2x2_ASAP7_75t_L g107 ( .A(n_95), .B(n_98), .Y(n_107) );
OR2x2_ASAP7_75t_L g119 ( .A(n_95), .B(n_98), .Y(n_119) );
INVx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g150 ( .A(n_96), .B(n_98), .Y(n_150) );
INVx1_ASAP7_75t_L g146 ( .A(n_97), .Y(n_146) );
AND2x2_ASAP7_75t_L g158 ( .A(n_97), .B(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx1_ASAP7_75t_L g112 ( .A(n_98), .Y(n_112) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x4_ASAP7_75t_L g137 ( .A(n_102), .B(n_118), .Y(n_137) );
AND2x6_ASAP7_75t_L g140 ( .A(n_102), .B(n_107), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_105), .B1(n_110), .B2(n_111), .Y(n_103) );
BUFx2_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g152 ( .A(n_109), .Y(n_152) );
OR2x6_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g133 ( .A(n_113), .Y(n_133) );
INVx4_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx11_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_129), .B2(n_130), .Y(n_124) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_SL g130 ( .A(n_131), .Y(n_130) );
BUFx2_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B1(n_147), .B2(n_148), .Y(n_141) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x4_ASAP7_75t_L g157 ( .A(n_145), .B(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g162 ( .A(n_145), .B(n_163), .Y(n_162) );
OR2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g163 ( .A(n_159), .Y(n_163) );
BUFx4f_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
BUFx12f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g166 ( .A1(n_167), .A2(n_170), .B1(n_171), .B2(n_174), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_167), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
AND3x1_ASAP7_75t_SL g177 ( .A(n_178), .B(n_183), .C(n_186), .Y(n_177) );
INVxp67_ASAP7_75t_L g487 ( .A(n_178), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx1_ASAP7_75t_SL g489 ( .A(n_183), .Y(n_489) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_183), .A2(n_225), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g499 ( .A(n_183), .Y(n_499) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_184), .B(n_187), .Y(n_493) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OR2x2_ASAP7_75t_SL g498 ( .A(n_186), .B(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_191), .B(n_423), .Y(n_190) );
AND4x1_ASAP7_75t_L g191 ( .A(n_192), .B(n_363), .C(n_378), .D(n_403), .Y(n_191) );
NOR2xp33_ASAP7_75t_SL g192 ( .A(n_193), .B(n_336), .Y(n_192) );
OAI21xp33_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_244), .B(n_316), .Y(n_193) );
AND2x2_ASAP7_75t_L g366 ( .A(n_194), .B(n_262), .Y(n_366) );
AND2x2_ASAP7_75t_L g379 ( .A(n_194), .B(n_261), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_194), .B(n_245), .Y(n_429) );
INVx1_ASAP7_75t_L g433 ( .A(n_194), .Y(n_433) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_229), .Y(n_194) );
INVx2_ASAP7_75t_L g350 ( .A(n_195), .Y(n_350) );
BUFx2_ASAP7_75t_L g377 ( .A(n_195), .Y(n_377) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_203), .B(n_227), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_196), .B(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_196), .B(n_260), .Y(n_259) );
AO21x2_ASAP7_75t_L g296 ( .A1(n_196), .A2(n_297), .B(n_304), .Y(n_296) );
INVx4_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_197), .A2(n_284), .B(n_285), .Y(n_283) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_197), .Y(n_324) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g306 ( .A(n_198), .Y(n_306) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
AND2x2_ASAP7_75t_SL g258 ( .A(n_199), .B(n_200), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_223), .Y(n_203) );
INVx5_ASAP7_75t_L g234 ( .A(n_205), .Y(n_234) );
AND2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_208), .Y(n_205) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_206), .Y(n_219) );
BUFx3_ASAP7_75t_L g242 ( .A(n_206), .Y(n_242) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g226 ( .A(n_207), .Y(n_226) );
INVx1_ASAP7_75t_L g292 ( .A(n_207), .Y(n_292) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_209), .Y(n_214) );
INVx3_ASAP7_75t_L g217 ( .A(n_209), .Y(n_217) );
AND2x2_ASAP7_75t_L g225 ( .A(n_209), .B(n_226), .Y(n_225) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_209), .Y(n_240) );
INVx1_ASAP7_75t_L g288 ( .A(n_209), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_215), .C(n_218), .Y(n_210) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g255 ( .A(n_214), .Y(n_255) );
INVx2_ASAP7_75t_L g236 ( .A(n_216), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_216), .B(n_330), .Y(n_329) );
INVx5_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_SL g232 ( .A1(n_221), .A2(n_233), .B(n_234), .C(n_235), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_221), .A2(n_234), .B(n_327), .C(n_328), .Y(n_326) );
INVx4_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
AND2x4_ASAP7_75t_L g224 ( .A(n_222), .B(n_225), .Y(n_224) );
BUFx3_ASAP7_75t_L g272 ( .A(n_222), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_222), .B(n_225), .Y(n_299) );
BUFx2_ASAP7_75t_L g265 ( .A(n_224), .Y(n_265) );
INVx1_ASAP7_75t_L g271 ( .A(n_226), .Y(n_271) );
AND2x2_ASAP7_75t_L g317 ( .A(n_229), .B(n_262), .Y(n_317) );
INVx2_ASAP7_75t_L g333 ( .A(n_229), .Y(n_333) );
AND2x2_ASAP7_75t_L g342 ( .A(n_229), .B(n_261), .Y(n_342) );
AND2x2_ASAP7_75t_L g421 ( .A(n_229), .B(n_350), .Y(n_421) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_243), .Y(n_229) );
INVx2_ASAP7_75t_L g251 ( .A(n_234), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx4_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_242), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_278), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_245), .B(n_348), .Y(n_386) );
INVx1_ASAP7_75t_L g474 ( .A(n_245), .Y(n_474) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_261), .Y(n_245) );
AND2x2_ASAP7_75t_L g332 ( .A(n_246), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g346 ( .A(n_246), .B(n_347), .Y(n_346) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_246), .Y(n_375) );
OR2x2_ASAP7_75t_L g407 ( .A(n_246), .B(n_349), .Y(n_407) );
AND2x2_ASAP7_75t_L g415 ( .A(n_246), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g448 ( .A(n_246), .B(n_417), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_246), .B(n_317), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_246), .B(n_377), .Y(n_473) );
AND2x2_ASAP7_75t_L g479 ( .A(n_246), .B(n_366), .Y(n_479) );
INVx5_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
BUFx2_ASAP7_75t_L g339 ( .A(n_247), .Y(n_339) );
AND2x2_ASAP7_75t_L g369 ( .A(n_247), .B(n_349), .Y(n_369) );
AND2x2_ASAP7_75t_L g402 ( .A(n_247), .B(n_362), .Y(n_402) );
AND2x2_ASAP7_75t_L g422 ( .A(n_247), .B(n_262), .Y(n_422) );
AND2x2_ASAP7_75t_L g456 ( .A(n_247), .B(n_322), .Y(n_456) );
OR2x6_ASAP7_75t_L g247 ( .A(n_248), .B(n_259), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_250), .B(n_258), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_256), .C(n_257), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_254), .A2(n_257), .B(n_313), .C(n_314), .Y(n_312) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g274 ( .A(n_258), .Y(n_274) );
INVx1_ASAP7_75t_L g277 ( .A(n_258), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_258), .A2(n_310), .B(n_311), .Y(n_309) );
AND2x4_ASAP7_75t_L g362 ( .A(n_261), .B(n_333), .Y(n_362) );
AND2x2_ASAP7_75t_L g373 ( .A(n_261), .B(n_369), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_261), .B(n_349), .Y(n_412) );
INVx2_ASAP7_75t_L g427 ( .A(n_261), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_261), .B(n_361), .Y(n_450) );
AND2x2_ASAP7_75t_L g469 ( .A(n_261), .B(n_421), .Y(n_469) );
INVx5_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_262), .Y(n_368) );
AND2x2_ASAP7_75t_L g376 ( .A(n_262), .B(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g417 ( .A(n_262), .B(n_333), .Y(n_417) );
OR2x6_ASAP7_75t_L g262 ( .A(n_263), .B(n_275), .Y(n_262) );
AOI21xp5_ASAP7_75t_SL g263 ( .A1(n_264), .A2(n_266), .B(n_273), .Y(n_263) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_265), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B(n_270), .Y(n_267) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_293), .Y(n_279) );
AND2x2_ASAP7_75t_L g340 ( .A(n_280), .B(n_323), .Y(n_340) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_281), .B(n_296), .Y(n_320) );
OR2x2_ASAP7_75t_L g353 ( .A(n_281), .B(n_323), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_281), .B(n_323), .Y(n_358) );
AND2x2_ASAP7_75t_L g385 ( .A(n_281), .B(n_322), .Y(n_385) );
AND2x2_ASAP7_75t_L g437 ( .A(n_281), .B(n_295), .Y(n_437) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_282), .B(n_307), .Y(n_345) );
AND2x2_ASAP7_75t_L g381 ( .A(n_282), .B(n_296), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_289), .B(n_290), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_290), .A2(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_293), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g371 ( .A(n_294), .B(n_353), .Y(n_371) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_307), .Y(n_294) );
OAI322xp33_ASAP7_75t_L g336 ( .A1(n_295), .A2(n_337), .A3(n_341), .B1(n_343), .B2(n_346), .C1(n_351), .C2(n_359), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_295), .B(n_322), .Y(n_344) );
OR2x2_ASAP7_75t_L g354 ( .A(n_295), .B(n_308), .Y(n_354) );
AND2x2_ASAP7_75t_L g356 ( .A(n_295), .B(n_308), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_295), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_295), .B(n_323), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_295), .B(n_452), .Y(n_451) );
INVx5_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_296), .B(n_340), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_300), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_307), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g334 ( .A(n_307), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_307), .B(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g396 ( .A(n_307), .B(n_323), .Y(n_396) );
AOI211xp5_ASAP7_75t_SL g424 ( .A1(n_307), .A2(n_425), .B(n_428), .C(n_440), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_307), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g462 ( .A(n_307), .B(n_437), .Y(n_462) );
INVx5_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g390 ( .A(n_308), .B(n_323), .Y(n_390) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_308), .Y(n_399) );
AND2x2_ASAP7_75t_L g439 ( .A(n_308), .B(n_437), .Y(n_439) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_308), .B(n_340), .Y(n_470) );
AND2x2_ASAP7_75t_L g477 ( .A(n_308), .B(n_436), .Y(n_477) );
OR2x6_ASAP7_75t_L g308 ( .A(n_309), .B(n_315), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_332), .B2(n_334), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_317), .B(n_339), .Y(n_387) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g335 ( .A(n_320), .Y(n_335) );
OR2x2_ASAP7_75t_L g395 ( .A(n_320), .B(n_396), .Y(n_395) );
OAI221xp5_ASAP7_75t_SL g443 ( .A1(n_320), .A2(n_444), .B1(n_446), .B2(n_447), .C(n_449), .Y(n_443) );
INVx2_ASAP7_75t_L g382 ( .A(n_321), .Y(n_382) );
AND2x2_ASAP7_75t_L g355 ( .A(n_322), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g445 ( .A(n_322), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_322), .B(n_437), .Y(n_458) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVxp67_ASAP7_75t_L g400 ( .A(n_323), .Y(n_400) );
AND2x2_ASAP7_75t_L g436 ( .A(n_323), .B(n_437), .Y(n_436) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B(n_331), .Y(n_323) );
AND2x2_ASAP7_75t_L g438 ( .A(n_332), .B(n_377), .Y(n_438) );
AND2x2_ASAP7_75t_L g348 ( .A(n_333), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_333), .B(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_SL g419 ( .A(n_335), .B(n_382), .Y(n_419) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g425 ( .A(n_338), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
OR2x2_ASAP7_75t_L g411 ( .A(n_339), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g476 ( .A(n_339), .B(n_421), .Y(n_476) );
INVx2_ASAP7_75t_L g409 ( .A(n_340), .Y(n_409) );
NAND4xp25_ASAP7_75t_SL g472 ( .A(n_341), .B(n_473), .C(n_474), .D(n_475), .Y(n_472) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_342), .B(n_406), .Y(n_441) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_SL g478 ( .A(n_345), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g440 ( .A1(n_346), .A2(n_409), .B(n_413), .C(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g435 ( .A(n_348), .B(n_427), .Y(n_435) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_349), .Y(n_361) );
INVx1_ASAP7_75t_L g416 ( .A(n_349), .Y(n_416) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_350), .Y(n_393) );
AOI211xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B(n_355), .C(n_357), .Y(n_351) );
AND2x2_ASAP7_75t_L g372 ( .A(n_352), .B(n_356), .Y(n_372) );
OAI322xp33_ASAP7_75t_SL g410 ( .A1(n_352), .A2(n_411), .A3(n_413), .B1(n_414), .B2(n_418), .C1(n_419), .C2(n_420), .Y(n_410) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g432 ( .A(n_354), .B(n_358), .Y(n_432) );
INVx1_ASAP7_75t_L g413 ( .A(n_356), .Y(n_413) );
INVx1_ASAP7_75t_SL g431 ( .A(n_358), .Y(n_431) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
AOI222xp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_370), .B1(n_372), .B2(n_373), .C1(n_374), .C2(n_501), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_365), .B(n_367), .Y(n_364) );
OAI322xp33_ASAP7_75t_L g453 ( .A1(n_365), .A2(n_427), .A3(n_432), .B1(n_454), .B2(n_455), .C1(n_457), .C2(n_458), .Y(n_453) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_366), .A2(n_380), .B1(n_404), .B2(n_408), .C(n_410), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OAI222xp33_ASAP7_75t_L g383 ( .A1(n_371), .A2(n_384), .B1(n_386), .B2(n_387), .C1(n_388), .C2(n_391), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_373), .A2(n_380), .B1(n_450), .B2(n_451), .Y(n_449) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
AOI211xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B(n_383), .C(n_394), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_380), .A2(n_417), .B(n_460), .C(n_463), .Y(n_459) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
AND2x2_ASAP7_75t_L g389 ( .A(n_381), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g452 ( .A(n_385), .Y(n_452) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_392), .B(n_417), .Y(n_446) );
BUFx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI21xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B(n_401), .Y(n_394) );
OAI221xp5_ASAP7_75t_SL g463 ( .A1(n_395), .A2(n_464), .B1(n_465), .B2(n_466), .C(n_467), .Y(n_463) );
INVxp33_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_399), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_406), .B(n_417), .Y(n_457) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AND2x2_ASAP7_75t_L g468 ( .A(n_421), .B(n_427), .Y(n_468) );
AND4x1_ASAP7_75t_L g423 ( .A(n_424), .B(n_442), .C(n_459), .D(n_471), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI221xp5_ASAP7_75t_SL g428 ( .A1(n_429), .A2(n_430), .B1(n_432), .B2(n_433), .C(n_434), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B1(n_438), .B2(n_439), .Y(n_434) );
INVx1_ASAP7_75t_L g464 ( .A(n_435), .Y(n_464) );
INVx1_ASAP7_75t_SL g454 ( .A(n_439), .Y(n_454) );
NOR2xp33_ASAP7_75t_SL g442 ( .A(n_443), .B(n_453), .Y(n_442) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_455), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_462), .A2(n_468), .B1(n_469), .B2(n_470), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_477), .B1(n_478), .B2(n_479), .Y(n_471) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI322xp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .A3(n_484), .B1(n_488), .B2(n_490), .C1(n_494), .C2(n_496), .Y(n_481) );
CKINVDCx14_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
endmodule