module real_aes_11524_n_329 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_329);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_329;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_1797;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1835;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_1787;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_399;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1802;
wire n_397;
wire n_1056;
wire n_1083;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_1352;
wire n_729;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g1194 ( .A(n_0), .Y(n_1194) );
INVx1_ASAP7_75t_L g925 ( .A(n_1), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_2), .A2(n_83), .B1(n_419), .B2(n_427), .Y(n_418) );
INVx1_ASAP7_75t_L g520 ( .A(n_2), .Y(n_520) );
INVx1_ASAP7_75t_L g1556 ( .A(n_3), .Y(n_1556) );
INVx1_ASAP7_75t_L g1440 ( .A(n_4), .Y(n_1440) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_4), .A2(n_127), .B1(n_1467), .B2(n_1468), .Y(n_1466) );
INVx1_ASAP7_75t_L g1413 ( .A(n_5), .Y(n_1413) );
INVx1_ASAP7_75t_L g1788 ( .A(n_6), .Y(n_1788) );
AOI22xp33_ASAP7_75t_L g1803 ( .A1(n_6), .A2(n_93), .B1(n_844), .B2(n_1804), .Y(n_1803) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_7), .A2(n_82), .B1(n_587), .B2(n_589), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_7), .A2(n_82), .B1(n_596), .B2(n_608), .C(n_610), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g904 ( .A1(n_8), .A2(n_241), .B1(n_561), .B2(n_564), .C(n_905), .Y(n_904) );
OAI22xp33_ASAP7_75t_L g913 ( .A1(n_8), .A2(n_90), .B1(n_738), .B2(n_740), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g1794 ( .A1(n_9), .A2(n_99), .B1(n_993), .B2(n_1795), .Y(n_1794) );
AOI22xp33_ASAP7_75t_SL g1801 ( .A1(n_9), .A2(n_99), .B1(n_799), .B2(n_1233), .Y(n_1801) );
INVx1_ASAP7_75t_L g1097 ( .A(n_10), .Y(n_1097) );
OAI211xp5_ASAP7_75t_SL g1117 ( .A1(n_10), .A2(n_589), .B(n_1118), .C(n_1124), .Y(n_1117) );
AOI221xp5_ASAP7_75t_L g832 ( .A1(n_11), .A2(n_271), .B1(n_498), .B2(n_564), .C(n_725), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_11), .A2(n_271), .B1(n_844), .B2(n_845), .Y(n_843) );
INVx1_ASAP7_75t_L g776 ( .A(n_12), .Y(n_776) );
AOI22xp33_ASAP7_75t_SL g792 ( .A1(n_12), .A2(n_260), .B1(n_793), .B2(n_795), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g1091 ( .A(n_13), .Y(n_1091) );
AO221x2_ASAP7_75t_L g1554 ( .A1(n_14), .A2(n_253), .B1(n_1531), .B2(n_1553), .C(n_1555), .Y(n_1554) );
OAI22xp33_ASAP7_75t_L g1041 ( .A1(n_15), .A2(n_63), .B1(n_419), .B2(n_427), .Y(n_1041) );
OAI22xp33_ASAP7_75t_L g1047 ( .A1(n_15), .A2(n_170), .B1(n_345), .B2(n_1027), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_16), .Y(n_688) );
CKINVDCx16_ASAP7_75t_R g1576 ( .A(n_17), .Y(n_1576) );
AOI21xp5_ASAP7_75t_L g1450 ( .A1(n_18), .A2(n_560), .B(n_561), .Y(n_1450) );
INVx1_ASAP7_75t_L g1453 ( .A(n_18), .Y(n_1453) );
XNOR2xp5_ASAP7_75t_L g651 ( .A(n_19), .B(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g1796 ( .A1(n_20), .A2(n_77), .B1(n_993), .B2(n_1797), .Y(n_1796) );
INVxp67_ASAP7_75t_SL g1816 ( .A(n_20), .Y(n_1816) );
INVx1_ASAP7_75t_L g1038 ( .A(n_21), .Y(n_1038) );
OAI222xp33_ASAP7_75t_L g1044 ( .A1(n_21), .A2(n_210), .B1(n_303), .B2(n_558), .C1(n_1045), .C2(n_1046), .Y(n_1044) );
OAI222xp33_ASAP7_75t_L g1186 ( .A1(n_22), .A2(n_61), .B1(n_129), .B2(n_976), .C1(n_1187), .C2(n_1190), .Y(n_1186) );
INVx1_ASAP7_75t_L g1207 ( .A(n_22), .Y(n_1207) );
CKINVDCx5p33_ASAP7_75t_R g1269 ( .A(n_23), .Y(n_1269) );
AOI22xp33_ASAP7_75t_SL g989 ( .A1(n_24), .A2(n_114), .B1(n_790), .B2(n_990), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_24), .A2(n_114), .B1(n_1000), .B2(n_1001), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g817 ( .A1(n_25), .A2(n_182), .B1(n_757), .B2(n_818), .C(n_819), .Y(n_817) );
INVx1_ASAP7_75t_L g852 ( .A(n_25), .Y(n_852) );
INVx1_ASAP7_75t_L g971 ( .A(n_26), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_26), .A2(n_306), .B1(n_723), .B2(n_725), .Y(n_996) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_27), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g518 ( .A(n_27), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g1094 ( .A(n_28), .Y(n_1094) );
CKINVDCx5p33_ASAP7_75t_R g752 ( .A(n_29), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g1242 ( .A1(n_30), .A2(n_140), .B1(n_1010), .B2(n_1011), .Y(n_1242) );
AOI22xp33_ASAP7_75t_SL g1259 ( .A1(n_30), .A2(n_140), .B1(n_763), .B2(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g336 ( .A(n_31), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g1445 ( .A(n_32), .Y(n_1445) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_33), .A2(n_98), .B1(n_409), .B2(n_1040), .Y(n_1039) );
AOI22xp33_ASAP7_75t_SL g1058 ( .A1(n_33), .A2(n_98), .B1(n_995), .B2(n_1000), .Y(n_1058) );
INVx1_ASAP7_75t_L g928 ( .A(n_34), .Y(n_928) );
OAI211xp5_ASAP7_75t_SL g950 ( .A1(n_34), .A2(n_589), .B(n_951), .C(n_956), .Y(n_950) );
AOI21xp33_ASAP7_75t_L g1438 ( .A1(n_35), .A2(n_498), .B(n_564), .Y(n_1438) );
INVx1_ASAP7_75t_L g1464 ( .A(n_35), .Y(n_1464) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_36), .A2(n_143), .B1(n_815), .B2(n_816), .Y(n_814) );
INVx1_ASAP7_75t_L g853 ( .A(n_36), .Y(n_853) );
INVxp67_ASAP7_75t_SL g1789 ( .A(n_37), .Y(n_1789) );
OAI22xp33_ASAP7_75t_L g1810 ( .A1(n_37), .A2(n_163), .B1(n_976), .B2(n_1187), .Y(n_1810) );
INVx1_ASAP7_75t_L g1478 ( .A(n_38), .Y(n_1478) );
AOI22xp33_ASAP7_75t_L g1506 ( .A1(n_38), .A2(n_196), .B1(n_723), .B2(n_1054), .Y(n_1506) );
INVx1_ASAP7_75t_L g1289 ( .A(n_39), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_39), .A2(n_263), .B1(n_1314), .B2(n_1317), .Y(n_1313) );
INVx1_ASAP7_75t_L g1049 ( .A(n_40), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_40), .A2(n_208), .B1(n_669), .B2(n_1075), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_41), .A2(n_132), .B1(n_1054), .B2(n_1216), .Y(n_1503) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_41), .A2(n_132), .B1(n_596), .B2(n_793), .Y(n_1509) );
CKINVDCx5p33_ASAP7_75t_R g1444 ( .A(n_42), .Y(n_1444) );
AOI22x1_ASAP7_75t_SL g1029 ( .A1(n_43), .A2(n_1030), .B1(n_1076), .B2(n_1077), .Y(n_1029) );
INVx1_ASAP7_75t_L g1076 ( .A(n_43), .Y(n_1076) );
INVx1_ASAP7_75t_L g1372 ( .A(n_44), .Y(n_1372) );
XNOR2xp5_ASAP7_75t_L g1080 ( .A(n_45), .B(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g877 ( .A(n_46), .Y(n_877) );
OAI221xp5_ASAP7_75t_L g887 ( .A1(n_46), .A2(n_587), .B1(n_712), .B2(n_888), .C(n_894), .Y(n_887) );
INVx1_ASAP7_75t_L g1142 ( .A(n_47), .Y(n_1142) );
OAI221xp5_ASAP7_75t_L g1159 ( .A1(n_47), .A2(n_589), .B1(n_1160), .B2(n_1165), .C(n_1170), .Y(n_1159) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_48), .A2(n_221), .B1(n_646), .B2(n_649), .Y(n_935) );
INVx1_ASAP7_75t_L g954 ( .A(n_48), .Y(n_954) );
AOI22xp5_ASAP7_75t_L g1582 ( .A1(n_49), .A2(n_304), .B1(n_1531), .B2(n_1553), .Y(n_1582) );
INVx1_ASAP7_75t_L g983 ( .A(n_50), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_50), .A2(n_167), .B1(n_993), .B2(n_995), .Y(n_992) );
INVx1_ASAP7_75t_L g721 ( .A(n_51), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g735 ( .A1(n_51), .A2(n_113), .B1(n_649), .B2(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g1303 ( .A(n_52), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_52), .A2(n_252), .B1(n_669), .B2(n_1075), .Y(n_1329) );
INVx1_ASAP7_75t_L g1305 ( .A(n_53), .Y(n_1305) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_53), .A2(n_286), .B1(n_1035), .B2(n_1067), .Y(n_1328) );
INVx1_ASAP7_75t_L g1211 ( .A(n_54), .Y(n_1211) );
AOI22xp33_ASAP7_75t_SL g1230 ( .A1(n_54), .A2(n_97), .B1(n_596), .B2(n_1231), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_55), .A2(n_328), .B1(n_669), .B2(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g702 ( .A(n_55), .Y(n_702) );
INVx1_ASAP7_75t_L g547 ( .A(n_56), .Y(n_547) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_56), .A2(n_228), .B1(n_596), .B2(n_598), .C(n_601), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_57), .B(n_811), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_58), .Y(n_1089) );
OAI22xp33_ASAP7_75t_L g748 ( .A1(n_59), .A2(n_291), .B1(n_695), .B2(n_696), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_59), .A2(n_291), .B1(n_469), .B2(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g1294 ( .A(n_60), .Y(n_1294) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_60), .A2(n_305), .B1(n_1019), .B2(n_1300), .Y(n_1299) );
AOI22xp33_ASAP7_75t_SL g1215 ( .A1(n_61), .A2(n_282), .B1(n_1003), .B2(n_1216), .Y(n_1215) );
AOI22xp33_ASAP7_75t_L g1502 ( .A1(n_62), .A2(n_177), .B1(n_993), .B2(n_1169), .Y(n_1502) );
AOI22xp33_ASAP7_75t_L g1508 ( .A1(n_62), .A2(n_177), .B1(n_684), .B2(n_1233), .Y(n_1508) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_63), .A2(n_124), .B1(n_1054), .B2(n_1060), .Y(n_1059) );
CKINVDCx5p33_ASAP7_75t_R g1136 ( .A(n_64), .Y(n_1136) );
INVxp33_ASAP7_75t_SL g1346 ( .A(n_65), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_65), .A2(n_318), .B1(n_1387), .B2(n_1389), .Y(n_1386) );
AOI22xp33_ASAP7_75t_SL g1053 ( .A1(n_66), .A2(n_136), .B1(n_564), .B2(n_1054), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_66), .A2(n_136), .B1(n_1067), .B2(n_1068), .Y(n_1066) );
OAI22xp33_ASAP7_75t_L g1104 ( .A1(n_67), .A2(n_319), .B1(n_883), .B2(n_884), .Y(n_1104) );
INVx1_ASAP7_75t_L g1126 ( .A(n_67), .Y(n_1126) );
INVx1_ASAP7_75t_L g1161 ( .A(n_68), .Y(n_1161) );
OAI22xp33_ASAP7_75t_L g1174 ( .A1(n_68), .A2(n_153), .B1(n_646), .B2(n_649), .Y(n_1174) );
INVx1_ASAP7_75t_L g932 ( .A(n_69), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_69), .A2(n_207), .B1(n_576), .B2(n_582), .Y(n_940) );
INVx1_ASAP7_75t_L g1479 ( .A(n_70), .Y(n_1479) );
AOI22xp33_ASAP7_75t_L g1505 ( .A1(n_70), .A2(n_152), .B1(n_892), .B2(n_993), .Y(n_1505) );
CKINVDCx5p33_ASAP7_75t_R g664 ( .A(n_71), .Y(n_664) );
INVxp67_ASAP7_75t_SL g1365 ( .A(n_72), .Y(n_1365) );
AOI221xp5_ASAP7_75t_L g1401 ( .A1(n_72), .A2(n_321), .B1(n_1402), .B2(n_1403), .C(n_1404), .Y(n_1401) );
INVx1_ASAP7_75t_L g1103 ( .A(n_73), .Y(n_1103) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_73), .A2(n_272), .B1(n_576), .B2(n_582), .Y(n_1108) );
XNOR2x2_ASAP7_75t_L g535 ( .A(n_74), .B(n_536), .Y(n_535) );
INVxp67_ASAP7_75t_SL g1783 ( .A(n_75), .Y(n_1783) );
AOI22xp33_ASAP7_75t_L g1806 ( .A1(n_75), .A2(n_233), .B1(n_881), .B2(n_1233), .Y(n_1806) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_76), .Y(n_563) );
INVxp33_ASAP7_75t_L g1815 ( .A(n_77), .Y(n_1815) );
BUFx2_ASAP7_75t_L g361 ( .A(n_78), .Y(n_361) );
BUFx2_ASAP7_75t_L g459 ( .A(n_78), .Y(n_459) );
INVx1_ASAP7_75t_L g530 ( .A(n_78), .Y(n_530) );
OR2x2_ASAP7_75t_L g1353 ( .A(n_78), .B(n_574), .Y(n_1353) );
AOI22xp33_ASAP7_75t_SL g1056 ( .A1(n_79), .A2(n_217), .B1(n_995), .B2(n_1057), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_79), .A2(n_217), .B1(n_1064), .B2(n_1065), .Y(n_1063) );
INVx1_ASAP7_75t_L g1431 ( .A(n_80), .Y(n_1431) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_80), .A2(n_116), .B1(n_670), .B2(n_1065), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_81), .A2(n_313), .B1(n_596), .B2(n_793), .Y(n_988) );
AOI22xp33_ASAP7_75t_SL g1002 ( .A1(n_81), .A2(n_313), .B1(n_723), .B2(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g398 ( .A(n_83), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_84), .A2(n_325), .B1(n_1057), .B2(n_1312), .Y(n_1311) );
AOI22xp33_ASAP7_75t_SL g1322 ( .A1(n_84), .A2(n_325), .B1(n_1323), .B2(n_1324), .Y(n_1322) );
INVx1_ASAP7_75t_L g1166 ( .A(n_85), .Y(n_1166) );
OAI22xp33_ASAP7_75t_L g1175 ( .A1(n_85), .A2(n_178), .B1(n_738), .B2(n_740), .Y(n_1175) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_86), .A2(n_144), .B1(n_974), .B2(n_976), .Y(n_973) );
OAI22xp33_ASAP7_75t_L g1017 ( .A1(n_86), .A2(n_144), .B1(n_1018), .B2(n_1019), .Y(n_1017) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_87), .Y(n_545) );
INVx1_ASAP7_75t_L g1145 ( .A(n_88), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_88), .A2(n_94), .B1(n_576), .B2(n_582), .Y(n_1150) );
OAI221xp5_ASAP7_75t_L g1348 ( .A1(n_89), .A2(n_169), .B1(n_1349), .B2(n_1354), .C(n_1356), .Y(n_1348) );
OAI22xp5_ASAP7_75t_L g1392 ( .A1(n_89), .A2(n_169), .B1(n_1393), .B2(n_1396), .Y(n_1392) );
INVx1_ASAP7_75t_L g901 ( .A(n_90), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g1798 ( .A1(n_91), .A2(n_185), .B1(n_723), .B2(n_1799), .Y(n_1798) );
INVxp67_ASAP7_75t_SL g1809 ( .A(n_91), .Y(n_1809) );
INVx1_ASAP7_75t_L g1291 ( .A(n_92), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_92), .A2(n_110), .B1(n_1206), .B2(n_1319), .Y(n_1318) );
INVxp33_ASAP7_75t_L g1785 ( .A(n_93), .Y(n_1785) );
INVx1_ASAP7_75t_L g1144 ( .A(n_94), .Y(n_1144) );
AO221x1_ASAP7_75t_L g1264 ( .A1(n_95), .A2(n_181), .B1(n_560), .B2(n_561), .C(n_1004), .Y(n_1264) );
INVx1_ASAP7_75t_L g1273 ( .A(n_95), .Y(n_1273) );
INVx1_ASAP7_75t_L g1202 ( .A(n_96), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_96), .A2(n_199), .B1(n_1011), .B2(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1205 ( .A(n_97), .Y(n_1205) );
XNOR2x2_ASAP7_75t_L g1281 ( .A(n_100), .B(n_1282), .Y(n_1281) );
CKINVDCx16_ASAP7_75t_R g1578 ( .A(n_101), .Y(n_1578) );
AO22x2_ASAP7_75t_L g1181 ( .A1(n_102), .A2(n_1182), .B1(n_1183), .B2(n_1234), .Y(n_1181) );
INVxp67_ASAP7_75t_SL g1182 ( .A(n_102), .Y(n_1182) );
INVx1_ASAP7_75t_L g927 ( .A(n_103), .Y(n_927) );
OAI221xp5_ASAP7_75t_L g941 ( .A1(n_103), .A2(n_587), .B1(n_942), .B2(n_945), .C(n_949), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_104), .A2(n_257), .B1(n_793), .B2(n_1244), .Y(n_1243) );
AOI221xp5_ASAP7_75t_L g1261 ( .A1(n_104), .A2(n_257), .B1(n_498), .B2(n_564), .C(n_905), .Y(n_1261) );
AOI22xp5_ASAP7_75t_L g1829 ( .A1(n_105), .A2(n_1830), .B1(n_1831), .B2(n_1832), .Y(n_1829) );
CKINVDCx5p33_ASAP7_75t_R g1831 ( .A(n_105), .Y(n_1831) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_106), .A2(n_183), .B1(n_1216), .B2(n_1224), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_106), .A2(n_183), .B1(n_596), .B2(n_793), .Y(n_1226) );
OAI22xp33_ASAP7_75t_L g685 ( .A1(n_107), .A2(n_176), .B1(n_625), .B2(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g730 ( .A(n_107), .Y(n_730) );
INVx1_ASAP7_75t_L g1139 ( .A(n_108), .Y(n_1139) );
CKINVDCx5p33_ASAP7_75t_R g871 ( .A(n_109), .Y(n_871) );
INVx1_ASAP7_75t_L g1285 ( .A(n_110), .Y(n_1285) );
OA22x2_ASAP7_75t_L g358 ( .A1(n_111), .A2(n_359), .B1(n_533), .B2(n_534), .Y(n_358) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_111), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g1552 ( .A1(n_112), .A2(n_298), .B1(n_1531), .B2(n_1553), .Y(n_1552) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_113), .A2(n_279), .B1(n_561), .B2(n_723), .C(n_724), .Y(n_722) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_115), .Y(n_764) );
INVx1_ASAP7_75t_L g1432 ( .A(n_116), .Y(n_1432) );
INVx1_ASAP7_75t_L g1494 ( .A(n_117), .Y(n_1494) );
AOI22xp33_ASAP7_75t_SL g1511 ( .A1(n_117), .A2(n_288), .B1(n_596), .B2(n_1231), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_118), .A2(n_146), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
INVx1_ASAP7_75t_L g1022 ( .A(n_118), .Y(n_1022) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_119), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g1592 ( .A1(n_120), .A2(n_122), .B1(n_1547), .B2(n_1550), .Y(n_1592) );
INVx1_ASAP7_75t_L g774 ( .A(n_121), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_121), .A2(n_264), .B1(n_790), .B2(n_791), .Y(n_789) );
INVx1_ASAP7_75t_L g716 ( .A(n_123), .Y(n_716) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_123), .A2(n_279), .B1(n_738), .B2(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g1034 ( .A(n_124), .Y(n_1034) );
AOI22xp5_ASAP7_75t_L g1593 ( .A1(n_125), .A2(n_309), .B1(n_1525), .B2(n_1594), .Y(n_1593) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_126), .Y(n_399) );
INVx1_ASAP7_75t_L g1436 ( .A(n_127), .Y(n_1436) );
CKINVDCx5p33_ASAP7_75t_R g1449 ( .A(n_128), .Y(n_1449) );
INVx1_ASAP7_75t_L g1209 ( .A(n_129), .Y(n_1209) );
XOR2xp5_ASAP7_75t_L g1332 ( .A(n_130), .B(n_1333), .Y(n_1332) );
AO221x2_ASAP7_75t_L g1524 ( .A1(n_131), .A2(n_192), .B1(n_1525), .B2(n_1531), .C(n_1532), .Y(n_1524) );
INVx1_ASAP7_75t_L g1530 ( .A(n_133), .Y(n_1530) );
INVx1_ASAP7_75t_L g1677 ( .A(n_134), .Y(n_1677) );
OAI22xp33_ASAP7_75t_L g882 ( .A1(n_135), .A2(n_307), .B1(n_883), .B2(n_884), .Y(n_882) );
INVx1_ASAP7_75t_L g907 ( .A(n_135), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g1581 ( .A1(n_137), .A2(n_317), .B1(n_1547), .B2(n_1550), .Y(n_1581) );
INVx1_ASAP7_75t_L g1489 ( .A(n_138), .Y(n_1489) );
AOI22xp33_ASAP7_75t_L g1512 ( .A1(n_138), .A2(n_175), .B1(n_641), .B2(n_684), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_139), .A2(n_324), .B1(n_683), .B2(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g890 ( .A(n_139), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_141), .A2(n_283), .B1(n_720), .B2(n_815), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_141), .A2(n_283), .B1(n_603), .B2(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g781 ( .A(n_142), .Y(n_781) );
INVx1_ASAP7_75t_L g849 ( .A(n_143), .Y(n_849) );
INVx1_ASAP7_75t_L g1786 ( .A(n_145), .Y(n_1786) );
INVx1_ASAP7_75t_L g1023 ( .A(n_146), .Y(n_1023) );
INVx1_ASAP7_75t_L g922 ( .A(n_147), .Y(n_922) );
INVx1_ASAP7_75t_L g1528 ( .A(n_148), .Y(n_1528) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_148), .B(n_1538), .Y(n_1541) );
AOI221xp5_ASAP7_75t_L g1446 ( .A1(n_149), .A2(n_281), .B1(n_1000), .B2(n_1447), .C(n_1448), .Y(n_1446) );
INVx1_ASAP7_75t_L g1456 ( .A(n_149), .Y(n_1456) );
INVx1_ASAP7_75t_L g878 ( .A(n_150), .Y(n_878) );
OAI211xp5_ASAP7_75t_SL g898 ( .A1(n_150), .A2(n_589), .B(n_899), .C(n_906), .Y(n_898) );
INVx2_ASAP7_75t_L g348 ( .A(n_151), .Y(n_348) );
INVx1_ASAP7_75t_L g1482 ( .A(n_152), .Y(n_1482) );
INVx1_ASAP7_75t_L g1167 ( .A(n_153), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_154), .A2(n_243), .B1(n_1000), .B2(n_1220), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_154), .A2(n_243), .B1(n_1011), .B2(n_1228), .Y(n_1227) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_155), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_156), .A2(n_320), .B1(n_681), .B2(n_684), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_156), .A2(n_320), .B1(n_695), .B2(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g417 ( .A(n_157), .Y(n_417) );
BUFx3_ASAP7_75t_L g433 ( .A(n_157), .Y(n_433) );
INVx1_ASAP7_75t_L g903 ( .A(n_158), .Y(n_903) );
OAI22xp33_ASAP7_75t_L g912 ( .A1(n_158), .A2(n_241), .B1(n_649), .B2(n_736), .Y(n_912) );
INVx1_ASAP7_75t_L g831 ( .A(n_159), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_159), .A2(n_235), .B1(n_629), .B2(n_634), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_160), .Y(n_445) );
INVx1_ASAP7_75t_L g1533 ( .A(n_161), .Y(n_1533) );
CKINVDCx5p33_ASAP7_75t_R g1267 ( .A(n_162), .Y(n_1267) );
INVx1_ASAP7_75t_L g1790 ( .A(n_163), .Y(n_1790) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_164), .Y(n_406) );
INVxp33_ASAP7_75t_SL g1341 ( .A(n_165), .Y(n_1341) );
AOI221xp5_ASAP7_75t_L g1380 ( .A1(n_165), .A2(n_273), .B1(n_1067), .B2(n_1381), .C(n_1383), .Y(n_1380) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_166), .A2(n_294), .B1(n_576), .B2(n_582), .Y(n_575) );
INVx1_ASAP7_75t_L g614 ( .A(n_166), .Y(n_614) );
INVx1_ASAP7_75t_L g985 ( .A(n_167), .Y(n_985) );
OAI221xp5_ASAP7_75t_L g1483 ( .A1(n_168), .A2(n_227), .B1(n_976), .B2(n_1484), .C(n_1485), .Y(n_1483) );
INVx1_ASAP7_75t_L g1492 ( .A(n_168), .Y(n_1492) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_170), .A2(n_210), .B1(n_1070), .B2(n_1072), .Y(n_1069) );
CKINVDCx5p33_ASAP7_75t_R g1252 ( .A(n_171), .Y(n_1252) );
INVx1_ASAP7_75t_L g1675 ( .A(n_172), .Y(n_1675) );
AOI22xp33_ASAP7_75t_SL g1249 ( .A1(n_173), .A2(n_326), .B1(n_641), .B2(n_799), .Y(n_1249) );
INVx1_ASAP7_75t_L g1256 ( .A(n_173), .Y(n_1256) );
AOI221xp5_ASAP7_75t_L g1123 ( .A1(n_174), .A2(n_327), .B1(n_564), .B2(n_725), .C(n_757), .Y(n_1123) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_174), .A2(n_266), .B1(n_738), .B2(n_740), .Y(n_1129) );
INVx1_ASAP7_75t_L g1490 ( .A(n_175), .Y(n_1490) );
INVx1_ASAP7_75t_L g727 ( .A(n_176), .Y(n_727) );
INVx1_ASAP7_75t_L g1164 ( .A(n_178), .Y(n_1164) );
INVx1_ASAP7_75t_L g1539 ( .A(n_179), .Y(n_1539) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_180), .Y(n_755) );
INVx1_ASAP7_75t_L g1275 ( .A(n_181), .Y(n_1275) );
INVx1_ASAP7_75t_L g850 ( .A(n_182), .Y(n_850) );
INVx1_ASAP7_75t_L g457 ( .A(n_184), .Y(n_457) );
INVx1_ASAP7_75t_L g623 ( .A(n_184), .Y(n_623) );
INVxp33_ASAP7_75t_L g1812 ( .A(n_185), .Y(n_1812) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_186), .A2(n_248), .B1(n_738), .B2(n_740), .Y(n_936) );
AOI221xp5_ASAP7_75t_L g955 ( .A1(n_186), .A2(n_221), .B1(n_561), .B2(n_897), .C(n_905), .Y(n_955) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_187), .Y(n_476) );
INVx1_ASAP7_75t_L g1565 ( .A(n_188), .Y(n_1565) );
INVx1_ASAP7_75t_L g828 ( .A(n_189), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_189), .A2(n_231), .B1(n_603), .B2(n_673), .Y(n_847) );
CKINVDCx5p33_ASAP7_75t_R g766 ( .A(n_190), .Y(n_766) );
INVx1_ASAP7_75t_L g1374 ( .A(n_191), .Y(n_1374) );
XOR2x2_ASAP7_75t_L g745 ( .A(n_192), .B(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_193), .A2(n_302), .B1(n_596), .B2(n_1246), .Y(n_1245) );
OAI221xp5_ASAP7_75t_L g1263 ( .A1(n_193), .A2(n_589), .B1(n_1264), .B2(n_1265), .C(n_1268), .Y(n_1263) );
INVx1_ASAP7_75t_L g1096 ( .A(n_194), .Y(n_1096) );
OAI221xp5_ASAP7_75t_L g1109 ( .A1(n_194), .A2(n_587), .B1(n_712), .B2(n_1110), .C(n_1116), .Y(n_1109) );
CKINVDCx5p33_ASAP7_75t_R g981 ( .A(n_195), .Y(n_981) );
INVx1_ASAP7_75t_L g1486 ( .A(n_196), .Y(n_1486) );
INVxp67_ASAP7_75t_SL g1366 ( .A(n_197), .Y(n_1366) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_197), .A2(n_275), .B1(n_1070), .B2(n_1075), .Y(n_1405) );
CKINVDCx5p33_ASAP7_75t_R g1428 ( .A(n_198), .Y(n_1428) );
INVx1_ASAP7_75t_L g1201 ( .A(n_199), .Y(n_1201) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_200), .Y(n_568) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_200), .A2(n_616), .B1(n_624), .B2(n_625), .C(n_628), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g1426 ( .A(n_201), .Y(n_1426) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_202), .A2(n_223), .B1(n_732), .B2(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g857 ( .A(n_202), .Y(n_857) );
INVx1_ASAP7_75t_L g1148 ( .A(n_203), .Y(n_1148) );
AOI22xp5_ASAP7_75t_L g1546 ( .A1(n_204), .A2(n_276), .B1(n_1547), .B2(n_1550), .Y(n_1546) );
INVx1_ASAP7_75t_L g858 ( .A(n_205), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_206), .Y(n_924) );
INVx1_ASAP7_75t_L g930 ( .A(n_207), .Y(n_930) );
INVx1_ASAP7_75t_L g1050 ( .A(n_208), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_209), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g1481 ( .A(n_211), .Y(n_1481) );
OAI22xp33_ASAP7_75t_L g1146 ( .A1(n_212), .A2(n_300), .B1(n_883), .B2(n_884), .Y(n_1146) );
INVx1_ASAP7_75t_L g1172 ( .A(n_212), .Y(n_1172) );
CKINVDCx5p33_ASAP7_75t_R g1442 ( .A(n_213), .Y(n_1442) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_214), .A2(n_292), .B1(n_1015), .B2(n_1060), .Y(n_1310) );
AOI22xp33_ASAP7_75t_SL g1326 ( .A1(n_214), .A2(n_292), .B1(n_1035), .B2(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g679 ( .A(n_215), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g713 ( .A1(n_215), .A2(n_589), .B(n_714), .C(n_726), .Y(n_713) );
CKINVDCx16_ASAP7_75t_R g1561 ( .A(n_216), .Y(n_1561) );
AOI22xp33_ASAP7_75t_L g1823 ( .A1(n_216), .A2(n_1824), .B1(n_1828), .B2(n_1833), .Y(n_1823) );
INVx1_ASAP7_75t_L g864 ( .A(n_218), .Y(n_864) );
INVx1_ASAP7_75t_L g676 ( .A(n_219), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_219), .A2(n_587), .B1(n_698), .B2(n_707), .C(n_712), .Y(n_697) );
INVx1_ASAP7_75t_L g1141 ( .A(n_220), .Y(n_1141) );
OAI221xp5_ASAP7_75t_L g1151 ( .A1(n_220), .A2(n_587), .B1(n_712), .B2(n_1152), .C(n_1156), .Y(n_1151) );
INVx1_ASAP7_75t_L g920 ( .A(n_222), .Y(n_920) );
INVx1_ASAP7_75t_L g855 ( .A(n_223), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_224), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_225), .A2(n_245), .B1(n_366), .B2(n_374), .Y(n_365) );
INVx1_ASAP7_75t_L g490 ( .A(n_225), .Y(n_490) );
INVx1_ASAP7_75t_L g869 ( .A(n_226), .Y(n_869) );
AOI21xp33_ASAP7_75t_L g896 ( .A1(n_226), .A2(n_498), .B(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g1493 ( .A(n_227), .Y(n_1493) );
AOI21xp33_ASAP7_75t_L g549 ( .A1(n_228), .A2(n_498), .B(n_550), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g663 ( .A(n_229), .Y(n_663) );
OAI221xp5_ASAP7_75t_L g749 ( .A1(n_230), .A2(n_589), .B1(n_750), .B2(n_759), .C(n_765), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g797 ( .A1(n_230), .A2(n_301), .B1(n_608), .B2(n_795), .Y(n_797) );
INVx1_ASAP7_75t_L g829 ( .A(n_231), .Y(n_829) );
OAI211xp5_ASAP7_75t_L g380 ( .A1(n_232), .A2(n_381), .B(n_386), .C(n_393), .Y(n_380) );
INVx1_ASAP7_75t_L g486 ( .A(n_232), .Y(n_486) );
INVx1_ASAP7_75t_L g1782 ( .A(n_233), .Y(n_1782) );
XNOR2xp5_ASAP7_75t_L g861 ( .A(n_234), .B(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g821 ( .A(n_235), .Y(n_821) );
INVx1_ASAP7_75t_L g1135 ( .A(n_236), .Y(n_1135) );
AOI22xp33_ASAP7_75t_SL g879 ( .A1(n_237), .A2(n_267), .B1(n_880), .B2(n_881), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_237), .A2(n_267), .B1(n_695), .B2(n_696), .Y(n_886) );
BUFx3_ASAP7_75t_L g416 ( .A(n_238), .Y(n_416) );
INVx1_ASAP7_75t_L g426 ( .A(n_238), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g1429 ( .A(n_239), .Y(n_1429) );
INVx1_ASAP7_75t_L g938 ( .A(n_240), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g1251 ( .A(n_242), .Y(n_1251) );
AO22x2_ASAP7_75t_L g1474 ( .A1(n_244), .A2(n_1475), .B1(n_1513), .B2(n_1514), .Y(n_1474) );
INVxp67_ASAP7_75t_L g1513 ( .A(n_244), .Y(n_1513) );
INVx1_ASAP7_75t_L g488 ( .A(n_245), .Y(n_488) );
XNOR2xp5_ASAP7_75t_L g915 ( .A(n_246), .B(n_916), .Y(n_915) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_247), .Y(n_344) );
INVx1_ASAP7_75t_L g532 ( .A(n_247), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_247), .B(n_308), .Y(n_574) );
AND2x2_ASAP7_75t_L g578 ( .A(n_247), .B(n_370), .Y(n_578) );
INVx1_ASAP7_75t_L g953 ( .A(n_248), .Y(n_953) );
CKINVDCx5p33_ASAP7_75t_R g1266 ( .A(n_249), .Y(n_1266) );
INVx1_ASAP7_75t_L g1681 ( .A(n_250), .Y(n_1681) );
AOI21xp33_ASAP7_75t_L g559 ( .A1(n_251), .A2(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g639 ( .A(n_251), .Y(n_639) );
INVx1_ASAP7_75t_L g1302 ( .A(n_252), .Y(n_1302) );
XNOR2xp5_ASAP7_75t_L g966 ( .A(n_253), .B(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g1566 ( .A(n_254), .Y(n_1566) );
INVx2_ASAP7_75t_L g413 ( .A(n_255), .Y(n_413) );
OR2x2_ASAP7_75t_L g638 ( .A(n_255), .B(n_623), .Y(n_638) );
INVx1_ASAP7_75t_L g1679 ( .A(n_256), .Y(n_1679) );
CKINVDCx16_ASAP7_75t_R g1563 ( .A(n_258), .Y(n_1563) );
CKINVDCx5p33_ASAP7_75t_R g1087 ( .A(n_259), .Y(n_1087) );
INVx1_ASAP7_75t_L g779 ( .A(n_260), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_261), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_262), .Y(n_467) );
INVx1_ASAP7_75t_L g1286 ( .A(n_263), .Y(n_1286) );
INVx1_ASAP7_75t_L g771 ( .A(n_264), .Y(n_771) );
INVx1_ASAP7_75t_L g1369 ( .A(n_265), .Y(n_1369) );
INVx1_ASAP7_75t_L g1119 ( .A(n_266), .Y(n_1119) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_268), .Y(n_553) );
INVx1_ASAP7_75t_L g1122 ( .A(n_269), .Y(n_1122) );
OAI22xp33_ASAP7_75t_L g1128 ( .A1(n_269), .A2(n_327), .B1(n_646), .B2(n_649), .Y(n_1128) );
INVx1_ASAP7_75t_L g1571 ( .A(n_270), .Y(n_1571) );
INVx1_ASAP7_75t_L g1100 ( .A(n_272), .Y(n_1100) );
INVxp33_ASAP7_75t_L g1344 ( .A(n_273), .Y(n_1344) );
INVx1_ASAP7_75t_L g1197 ( .A(n_274), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_274), .A2(n_285), .B1(n_993), .B2(n_1114), .Y(n_1217) );
INVxp33_ASAP7_75t_L g1360 ( .A(n_275), .Y(n_1360) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_277), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_278), .A2(n_293), .B1(n_596), .B2(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1025 ( .A(n_278), .Y(n_1025) );
AOI22x1_ASAP7_75t_L g1236 ( .A1(n_280), .A2(n_1237), .B1(n_1238), .B2(n_1276), .Y(n_1236) );
INVxp67_ASAP7_75t_SL g1276 ( .A(n_280), .Y(n_1276) );
INVx1_ASAP7_75t_L g1454 ( .A(n_281), .Y(n_1454) );
INVx1_ASAP7_75t_L g1193 ( .A(n_282), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g1793 ( .A1(n_284), .A2(n_322), .B1(n_723), .B2(n_724), .Y(n_1793) );
AOI22xp33_ASAP7_75t_L g1802 ( .A1(n_284), .A2(n_322), .B1(n_438), .B2(n_793), .Y(n_1802) );
INVx1_ASAP7_75t_L g1196 ( .A(n_285), .Y(n_1196) );
INVx1_ASAP7_75t_L g1298 ( .A(n_286), .Y(n_1298) );
INVx1_ASAP7_75t_L g1557 ( .A(n_287), .Y(n_1557) );
INVx1_ASAP7_75t_L g1499 ( .A(n_288), .Y(n_1499) );
CKINVDCx5p33_ASAP7_75t_R g1288 ( .A(n_289), .Y(n_1288) );
OAI22xp33_ASAP7_75t_L g933 ( .A1(n_290), .A2(n_312), .B1(n_883), .B2(n_884), .Y(n_933) );
INVx1_ASAP7_75t_L g959 ( .A(n_290), .Y(n_959) );
INVx1_ASAP7_75t_L g1014 ( .A(n_293), .Y(n_1014) );
INVx1_ASAP7_75t_L g611 ( .A(n_294), .Y(n_611) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_295), .Y(n_338) );
AND3x2_ASAP7_75t_L g1529 ( .A(n_295), .B(n_336), .C(n_1530), .Y(n_1529) );
NAND2xp5_ASAP7_75t_L g1536 ( .A(n_295), .B(n_336), .Y(n_1536) );
CKINVDCx5p33_ASAP7_75t_R g1106 ( .A(n_296), .Y(n_1106) );
INVx2_ASAP7_75t_L g349 ( .A(n_297), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g1138 ( .A(n_299), .Y(n_1138) );
INVx1_ASAP7_75t_L g1171 ( .A(n_300), .Y(n_1171) );
OAI221xp5_ASAP7_75t_L g768 ( .A1(n_301), .A2(n_587), .B1(n_712), .B2(n_769), .C(n_775), .Y(n_768) );
INVx1_ASAP7_75t_L g1262 ( .A(n_302), .Y(n_1262) );
CKINVDCx5p33_ASAP7_75t_R g1037 ( .A(n_303), .Y(n_1037) );
XNOR2xp5_ASAP7_75t_L g1130 ( .A(n_304), .B(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1292 ( .A(n_305), .Y(n_1292) );
INVx1_ASAP7_75t_L g978 ( .A(n_306), .Y(n_978) );
INVx1_ASAP7_75t_L g908 ( .A(n_307), .Y(n_908) );
INVx1_ASAP7_75t_L g351 ( .A(n_308), .Y(n_351) );
INVx2_ASAP7_75t_L g370 ( .A(n_308), .Y(n_370) );
AO22x2_ASAP7_75t_L g1422 ( .A1(n_309), .A2(n_1423), .B1(n_1471), .B2(n_1472), .Y(n_1422) );
INVxp67_ASAP7_75t_SL g1471 ( .A(n_309), .Y(n_1471) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_310), .Y(n_364) );
INVx1_ASAP7_75t_L g1375 ( .A(n_311), .Y(n_1375) );
INVx1_ASAP7_75t_L g957 ( .A(n_312), .Y(n_957) );
INVx1_ASAP7_75t_L g567 ( .A(n_314), .Y(n_567) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_314), .Y(n_624) );
OAI211xp5_ASAP7_75t_L g435 ( .A1(n_315), .A2(n_436), .B(n_441), .C(n_452), .Y(n_435) );
INVx1_ASAP7_75t_L g525 ( .A(n_315), .Y(n_525) );
INVx1_ASAP7_75t_L g1572 ( .A(n_316), .Y(n_1572) );
INVxp33_ASAP7_75t_SL g1337 ( .A(n_318), .Y(n_1337) );
INVx1_ASAP7_75t_L g1125 ( .A(n_319), .Y(n_1125) );
INVxp33_ASAP7_75t_SL g1362 ( .A(n_321), .Y(n_1362) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_323), .Y(n_767) );
INVx1_ASAP7_75t_L g893 ( .A(n_324), .Y(n_893) );
INVx1_ASAP7_75t_L g1257 ( .A(n_326), .Y(n_1257) );
INVx1_ASAP7_75t_L g706 ( .A(n_328), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_352), .B(n_1517), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx3_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_339), .Y(n_333) );
AND2x4_ASAP7_75t_L g1822 ( .A(n_334), .B(n_340), .Y(n_1822) );
NOR2xp33_ASAP7_75t_SL g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_SL g1827 ( .A(n_335), .Y(n_1827) );
NAND2xp5_ASAP7_75t_L g1838 ( .A(n_335), .B(n_337), .Y(n_1838) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g1826 ( .A(n_337), .B(n_1827), .Y(n_1826) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_345), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g360 ( .A(n_342), .B(n_361), .Y(n_360) );
OR2x6_ASAP7_75t_L g1028 ( .A(n_342), .B(n_361), .Y(n_1028) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g711 ( .A(n_343), .B(n_351), .Y(n_711) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g498 ( .A(n_344), .B(n_369), .Y(n_498) );
INVx8_ASAP7_75t_L g363 ( .A(n_345), .Y(n_363) );
OR2x6_ASAP7_75t_L g345 ( .A(n_346), .B(n_350), .Y(n_345) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_346), .Y(n_500) );
BUFx2_ASAP7_75t_L g948 ( .A(n_346), .Y(n_948) );
OR2x6_ASAP7_75t_L g1027 ( .A(n_346), .B(n_368), .Y(n_1027) );
INVx2_ASAP7_75t_SL g1158 ( .A(n_346), .Y(n_1158) );
INVx1_ASAP7_75t_L g1163 ( .A(n_346), .Y(n_1163) );
OR2x2_ASAP7_75t_L g1416 ( .A(n_346), .B(n_1353), .Y(n_1416) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx2_ASAP7_75t_L g373 ( .A(n_348), .Y(n_373) );
AND2x4_ASAP7_75t_L g378 ( .A(n_348), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g385 ( .A(n_348), .Y(n_385) );
INVx1_ASAP7_75t_L g392 ( .A(n_348), .Y(n_392) );
AND2x2_ASAP7_75t_L g397 ( .A(n_348), .B(n_349), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_349), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g379 ( .A(n_349), .Y(n_379) );
INVx1_ASAP7_75t_L g384 ( .A(n_349), .Y(n_384) );
INVx1_ASAP7_75t_L g401 ( .A(n_349), .Y(n_401) );
INVx1_ASAP7_75t_L g581 ( .A(n_349), .Y(n_581) );
AND2x4_ASAP7_75t_L g400 ( .A(n_350), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_351), .B(n_404), .Y(n_1019) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_351), .B(n_404), .Y(n_1046) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_1277), .B1(n_1278), .B2(n_1516), .Y(n_352) );
INVx1_ASAP7_75t_L g1516 ( .A(n_353), .Y(n_1516) );
XNOR2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_963), .Y(n_353) );
XOR2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_742), .Y(n_354) );
XNOR2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_650), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
XNOR2x1_ASAP7_75t_L g357 ( .A(n_358), .B(n_535), .Y(n_357) );
INVx1_ASAP7_75t_L g533 ( .A(n_359), .Y(n_533) );
OAI211xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B(n_407), .C(n_460), .Y(n_359) );
AND2x4_ASAP7_75t_L g493 ( .A(n_361), .B(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g642 ( .A(n_361), .B(n_643), .Y(n_642) );
AND2x4_ASAP7_75t_L g802 ( .A(n_361), .B(n_494), .Y(n_802) );
AOI211xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B(n_365), .C(n_380), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g1024 ( .A1(n_363), .A2(n_981), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_363), .A2(n_1026), .B1(n_1194), .B2(n_1211), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_363), .A2(n_1288), .B1(n_1305), .B2(n_1306), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_363), .A2(n_1306), .B1(n_1481), .B2(n_1499), .Y(n_1498) );
AOI22xp33_ASAP7_75t_L g1784 ( .A1(n_363), .A2(n_1306), .B1(n_1785), .B2(n_1786), .Y(n_1784) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_364), .A2(n_477), .B1(n_484), .B2(n_486), .Y(n_483) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_371), .Y(n_366) );
AOI322xp5_ASAP7_75t_L g393 ( .A1(n_367), .A2(n_394), .A3(n_398), .B1(n_399), .B2(n_400), .C1(n_402), .C2(n_406), .Y(n_393) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g375 ( .A(n_368), .B(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g1021 ( .A(n_368), .B(n_579), .Y(n_1021) );
AND2x4_ASAP7_75t_L g1203 ( .A(n_368), .B(n_376), .Y(n_1203) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g390 ( .A(n_370), .Y(n_390) );
INVx2_ASAP7_75t_L g506 ( .A(n_371), .Y(n_506) );
BUFx2_ASAP7_75t_L g1368 ( .A(n_371), .Y(n_1368) );
BUFx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g513 ( .A(n_372), .Y(n_513) );
INVx1_ASAP7_75t_L g541 ( .A(n_372), .Y(n_541) );
INVx1_ASAP7_75t_L g570 ( .A(n_373), .Y(n_570) );
AND2x4_ASAP7_75t_L g579 ( .A(n_373), .B(n_580), .Y(n_579) );
INVx5_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g1020 ( .A1(n_375), .A2(n_1021), .B1(n_1022), .B2(n_1023), .Y(n_1020) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_375), .A2(n_1021), .B1(n_1049), .B2(n_1050), .Y(n_1048) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g1155 ( .A(n_377), .Y(n_1155) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g509 ( .A(n_378), .Y(n_509) );
INVx3_ASAP7_75t_L g517 ( .A(n_378), .Y(n_517) );
BUFx6f_ASAP7_75t_L g763 ( .A(n_378), .Y(n_763) );
AND2x4_ASAP7_75t_L g391 ( .A(n_379), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g503 ( .A(n_383), .Y(n_503) );
INVx3_ASAP7_75t_L g548 ( .A(n_383), .Y(n_548) );
INVx2_ASAP7_75t_L g558 ( .A(n_383), .Y(n_558) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_384), .B(n_385), .Y(n_524) );
INVx1_ASAP7_75t_L g404 ( .A(n_385), .Y(n_404) );
NAND4xp25_ASAP7_75t_SL g1199 ( .A(n_386), .B(n_1200), .C(n_1204), .D(n_1210), .Y(n_1199) );
NAND4xp25_ASAP7_75t_SL g1487 ( .A(n_386), .B(n_1488), .C(n_1491), .D(n_1498), .Y(n_1487) );
NAND4xp25_ASAP7_75t_SL g1780 ( .A(n_386), .B(n_1781), .C(n_1784), .D(n_1787), .Y(n_1780) );
CKINVDCx11_ASAP7_75t_R g386 ( .A(n_387), .Y(n_386) );
AOI211xp5_ASAP7_75t_L g1013 ( .A1(n_387), .A2(n_1014), .B(n_1015), .C(n_1017), .Y(n_1013) );
NOR3xp33_ASAP7_75t_L g1043 ( .A(n_387), .B(n_1044), .C(n_1047), .Y(n_1043) );
AOI211xp5_ASAP7_75t_L g1297 ( .A1(n_387), .A2(n_1054), .B(n_1298), .C(n_1299), .Y(n_1297) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_391), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g405 ( .A(n_389), .Y(n_405) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2x1p5_ASAP7_75t_L g531 ( .A(n_390), .B(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g591 ( .A(n_391), .Y(n_591) );
BUFx6f_ASAP7_75t_L g725 ( .A(n_391), .Y(n_725) );
BUFx3_ASAP7_75t_L g905 ( .A(n_391), .Y(n_905) );
BUFx6f_ASAP7_75t_L g1004 ( .A(n_391), .Y(n_1004) );
BUFx2_ASAP7_75t_L g1497 ( .A(n_391), .Y(n_1497) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g1216 ( .A(n_395), .Y(n_1216) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_396), .Y(n_564) );
AND2x4_ASAP7_75t_L g588 ( .A(n_396), .B(n_578), .Y(n_588) );
BUFx2_ASAP7_75t_L g818 ( .A(n_396), .Y(n_818) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g551 ( .A(n_397), .Y(n_551) );
AOI322xp5_ASAP7_75t_L g441 ( .A1(n_399), .A2(n_406), .A3(n_442), .B1(n_444), .B2(n_445), .C1(n_446), .C2(n_450), .Y(n_441) );
INVx2_ASAP7_75t_L g1018 ( .A(n_400), .Y(n_1018) );
INVx2_ASAP7_75t_L g1045 ( .A(n_400), .Y(n_1045) );
INVx2_ASAP7_75t_L g1300 ( .A(n_400), .Y(n_1300) );
AOI222xp33_ASAP7_75t_L g1491 ( .A1(n_400), .A2(n_402), .B1(n_1492), .B2(n_1493), .C1(n_1494), .C2(n_1495), .Y(n_1491) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_401), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_566) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_401), .Y(n_729) );
INVx1_ASAP7_75t_L g825 ( .A(n_401), .Y(n_825) );
AOI222xp33_ASAP7_75t_L g1204 ( .A1(n_402), .A2(n_1205), .B1(n_1206), .B2(n_1207), .C1(n_1208), .C2(n_1209), .Y(n_1204) );
AOI222xp33_ASAP7_75t_L g1787 ( .A1(n_402), .A2(n_1206), .B1(n_1208), .B2(n_1788), .C1(n_1789), .C2(n_1790), .Y(n_1787) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g1271 ( .A1(n_403), .A2(n_824), .B1(n_1251), .B2(n_1252), .Y(n_1271) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI31xp33_ASAP7_75t_SL g407 ( .A1(n_408), .A2(n_418), .A3(n_435), .B(n_455), .Y(n_407) );
INVx4_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_410), .A2(n_983), .B1(n_984), .B2(n_985), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_410), .A2(n_984), .B1(n_1196), .B2(n_1197), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1287 ( .A1(n_410), .A2(n_428), .B1(n_1288), .B2(n_1289), .Y(n_1287) );
AOI22xp33_ASAP7_75t_L g1455 ( .A1(n_410), .A2(n_428), .B1(n_1426), .B2(n_1456), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1477 ( .A1(n_410), .A2(n_979), .B1(n_1478), .B2(n_1479), .Y(n_1477) );
AOI22xp33_ASAP7_75t_L g1814 ( .A1(n_410), .A2(n_984), .B1(n_1815), .B2(n_1816), .Y(n_1814) );
AND2x6_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .Y(n_410) );
AND2x4_ASAP7_75t_L g979 ( .A(n_411), .B(n_980), .Y(n_979) );
AND2x4_ASAP7_75t_L g1813 ( .A(n_411), .B(n_980), .Y(n_1813) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_412), .B(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g422 ( .A(n_413), .Y(n_422) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_413), .Y(n_430) );
AND2x2_ASAP7_75t_L g464 ( .A(n_413), .B(n_457), .Y(n_464) );
INVx2_ASAP7_75t_L g495 ( .A(n_413), .Y(n_495) );
INVx1_ASAP7_75t_L g491 ( .A(n_414), .Y(n_491) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_414), .Y(n_799) );
BUFx6f_ASAP7_75t_L g873 ( .A(n_414), .Y(n_873) );
BUFx6f_ASAP7_75t_L g881 ( .A(n_414), .Y(n_881) );
INVx2_ASAP7_75t_L g1325 ( .A(n_414), .Y(n_1325) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g474 ( .A(n_415), .Y(n_474) );
INVx1_ASAP7_75t_L g604 ( .A(n_415), .Y(n_604) );
INVx1_ASAP7_75t_L g647 ( .A(n_415), .Y(n_647) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_415), .Y(n_673) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx2_ASAP7_75t_L g434 ( .A(n_416), .Y(n_434) );
AND2x2_ASAP7_75t_L g440 ( .A(n_416), .B(n_433), .Y(n_440) );
INVx1_ASAP7_75t_L g424 ( .A(n_417), .Y(n_424) );
OR2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g444 ( .A(n_420), .Y(n_444) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g437 ( .A(n_421), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g454 ( .A(n_421), .Y(n_454) );
AND2x6_ASAP7_75t_L g984 ( .A(n_421), .B(n_443), .Y(n_984) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x6_ASAP7_75t_L g450 ( .A(n_422), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g478 ( .A(n_423), .Y(n_478) );
INVx1_ASAP7_75t_L g662 ( .A(n_423), .Y(n_662) );
BUFx2_ASAP7_75t_L g868 ( .A(n_423), .Y(n_868) );
OR2x2_ASAP7_75t_L g1410 ( .A(n_423), .B(n_638), .Y(n_1410) );
OR2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
AND2x2_ASAP7_75t_L g482 ( .A(n_424), .B(n_425), .Y(n_482) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g443 ( .A(n_426), .B(n_433), .Y(n_443) );
INVx4_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_428), .A2(n_978), .B1(n_979), .B2(n_981), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_428), .A2(n_979), .B1(n_1193), .B2(n_1194), .Y(n_1192) );
AOI221xp5_ASAP7_75t_L g1480 ( .A1(n_428), .A2(n_984), .B1(n_1481), .B2(n_1482), .C(n_1483), .Y(n_1480) );
AOI22xp33_ASAP7_75t_L g1811 ( .A1(n_428), .A2(n_1786), .B1(n_1812), .B2(n_1813), .Y(n_1811) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
AND2x2_ASAP7_75t_SL g446 ( .A(n_429), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g975 ( .A(n_429), .B(n_447), .Y(n_975) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx6_ASAP7_75t_L g600 ( .A(n_431), .Y(n_600) );
INVx2_ASAP7_75t_L g635 ( .A(n_431), .Y(n_635) );
AND2x2_ASAP7_75t_L g643 ( .A(n_431), .B(n_621), .Y(n_643) );
BUFx2_ASAP7_75t_L g844 ( .A(n_431), .Y(n_844) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g451 ( .A(n_432), .Y(n_451) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g449 ( .A(n_434), .Y(n_449) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI211xp5_ASAP7_75t_L g1808 ( .A1(n_437), .A2(n_453), .B(n_1809), .C(n_1810), .Y(n_1808) );
HB1xp67_ASAP7_75t_L g972 ( .A(n_438), .Y(n_972) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g453 ( .A(n_439), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g597 ( .A(n_439), .Y(n_597) );
INVx1_ASAP7_75t_L g657 ( .A(n_439), .Y(n_657) );
BUFx6f_ASAP7_75t_L g1073 ( .A(n_439), .Y(n_1073) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_440), .Y(n_630) );
INVx2_ASAP7_75t_L g470 ( .A(n_442), .Y(n_470) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_SL g489 ( .A(n_443), .Y(n_489) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_443), .Y(n_603) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_443), .Y(n_670) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_443), .Y(n_683) );
BUFx3_ASAP7_75t_L g880 ( .A(n_443), .Y(n_880) );
BUFx2_ASAP7_75t_L g1228 ( .A(n_443), .Y(n_1228) );
BUFx2_ASAP7_75t_L g1233 ( .A(n_443), .Y(n_1233) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_445), .A2(n_511), .B1(n_514), .B2(n_518), .Y(n_510) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g1189 ( .A(n_448), .Y(n_1189) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g618 ( .A(n_449), .Y(n_618) );
INVx3_ASAP7_75t_L g976 ( .A(n_450), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_450), .A2(n_975), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
AOI222xp33_ASAP7_75t_L g1290 ( .A1(n_450), .A2(n_1244), .B1(n_1291), .B2(n_1292), .C1(n_1293), .C2(n_1294), .Y(n_1290) );
AOI222xp33_ASAP7_75t_L g1457 ( .A1(n_450), .A2(n_1444), .B1(n_1445), .B2(n_1449), .C1(n_1458), .C2(n_1460), .Y(n_1457) );
BUFx3_ASAP7_75t_L g627 ( .A(n_451), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g1032 ( .A(n_452), .B(n_1033), .C(n_1036), .Y(n_1032) );
CKINVDCx8_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
AOI211xp5_ASAP7_75t_L g970 ( .A1(n_453), .A2(n_971), .B(n_972), .C(n_973), .Y(n_970) );
NOR2xp33_ASAP7_75t_L g1185 ( .A(n_453), .B(n_1186), .Y(n_1185) );
INVx5_ASAP7_75t_L g1295 ( .A(n_453), .Y(n_1295) );
OAI21xp33_ASAP7_75t_L g1485 ( .A1(n_454), .A2(n_1073), .B(n_1486), .Y(n_1485) );
OAI31xp33_ASAP7_75t_L g1031 ( .A1(n_455), .A2(n_1032), .A3(n_1039), .B(n_1041), .Y(n_1031) );
INVx1_ASAP7_75t_SL g1817 ( .A(n_455), .Y(n_1817) );
AND2x4_ASAP7_75t_L g455 ( .A(n_456), .B(n_458), .Y(n_455) );
AND2x4_ASAP7_75t_L g968 ( .A(n_456), .B(n_458), .Y(n_968) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g494 ( .A(n_457), .B(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g910 ( .A(n_458), .Y(n_910) );
BUFx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g465 ( .A(n_459), .Y(n_465) );
OR2x6_ASAP7_75t_L g497 ( .A(n_459), .B(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_496), .Y(n_460) );
OAI33xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_466), .A3(n_475), .B1(n_483), .B2(n_487), .B3(n_492), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_462), .A2(n_867), .B1(n_874), .B2(n_876), .Y(n_866) );
OAI33xp33_ASAP7_75t_L g918 ( .A1(n_462), .A2(n_492), .A3(n_919), .B1(n_923), .B2(n_926), .B3(n_929), .Y(n_918) );
OAI33xp33_ASAP7_75t_L g1084 ( .A1(n_462), .A2(n_492), .A3(n_1085), .B1(n_1090), .B2(n_1095), .B3(n_1098), .Y(n_1084) );
OAI33xp33_ASAP7_75t_L g1133 ( .A1(n_462), .A2(n_492), .A3(n_1134), .B1(n_1137), .B2(n_1140), .B3(n_1143), .Y(n_1133) );
INVx1_ASAP7_75t_SL g1241 ( .A(n_462), .Y(n_1241) );
OR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_465), .Y(n_462) );
OR2x6_ASAP7_75t_L g606 ( .A(n_463), .B(n_465), .Y(n_606) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g840 ( .A(n_464), .Y(n_840) );
INVx1_ASAP7_75t_L g1404 ( .A(n_464), .Y(n_1404) );
INVx2_ASAP7_75t_L g593 ( .A(n_465), .Y(n_593) );
BUFx2_ASAP7_75t_L g733 ( .A(n_465), .Y(n_733) );
OAI31xp33_ASAP7_75t_L g747 ( .A1(n_465), .A2(n_748), .A3(n_749), .B(n_768), .Y(n_747) );
OR2x2_ASAP7_75t_L g839 ( .A(n_465), .B(n_840), .Y(n_839) );
AND2x4_ASAP7_75t_L g1005 ( .A(n_465), .B(n_711), .Y(n_1005) );
AND2x4_ASAP7_75t_L g1052 ( .A(n_465), .B(n_711), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B1(n_471), .B2(n_472), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_467), .A2(n_471), .B1(n_505), .B2(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_470), .A2(n_611), .B1(n_612), .B2(n_614), .Y(n_610) );
INVx1_ASAP7_75t_L g1467 ( .A(n_470), .Y(n_1467) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g613 ( .A(n_474), .Y(n_613) );
OR2x2_ASAP7_75t_L g1412 ( .A(n_474), .B(n_638), .Y(n_1412) );
OAI22xp33_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_477), .B1(n_479), .B2(n_480), .Y(n_475) );
OAI22xp33_ASAP7_75t_L g499 ( .A1(n_476), .A2(n_479), .B1(n_500), .B2(n_501), .Y(n_499) );
OAI22xp33_ASAP7_75t_L g923 ( .A1(n_477), .A2(n_677), .B1(n_924), .B2(n_925), .Y(n_923) );
OAI22xp33_ASAP7_75t_L g926 ( .A1(n_477), .A2(n_870), .B1(n_927), .B2(n_928), .Y(n_926) );
OAI22xp33_ASAP7_75t_L g1140 ( .A1(n_477), .A2(n_484), .B1(n_1141), .B2(n_1142), .Y(n_1140) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g675 ( .A(n_478), .Y(n_675) );
INVx1_ASAP7_75t_L g739 ( .A(n_478), .Y(n_739) );
OAI221xp5_ASAP7_75t_L g876 ( .A1(n_480), .A2(n_868), .B1(n_877), .B2(n_878), .C(n_879), .Y(n_876) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g678 ( .A(n_481), .Y(n_678) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g485 ( .A(n_482), .Y(n_485) );
BUFx4f_ASAP7_75t_L g667 ( .A(n_482), .Y(n_667) );
INVx1_ASAP7_75t_L g1093 ( .A(n_482), .Y(n_1093) );
OAI22xp33_ASAP7_75t_L g1137 ( .A1(n_484), .A2(n_868), .B1(n_1138), .B2(n_1139), .Y(n_1137) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR2x6_ASAP7_75t_L g649 ( .A(n_485), .B(n_637), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g1095 ( .A1(n_485), .A2(n_661), .B1(n_1096), .B2(n_1097), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_487) );
INVx2_ASAP7_75t_L g641 ( .A(n_489), .Y(n_641) );
INVx1_ASAP7_75t_L g1010 ( .A(n_489), .Y(n_1010) );
OAI22xp5_ASAP7_75t_SL g658 ( .A1(n_492), .A2(n_606), .B1(n_659), .B2(n_674), .Y(n_658) );
INVx4_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_493), .A2(n_595), .B1(n_605), .B2(n_607), .C(n_615), .Y(n_594) );
BUFx4f_ASAP7_75t_L g875 ( .A(n_493), .Y(n_875) );
AOI33xp33_ASAP7_75t_L g1061 ( .A1(n_493), .A2(n_1062), .A3(n_1063), .B1(n_1066), .B2(n_1069), .B3(n_1074), .Y(n_1061) );
BUFx4f_ASAP7_75t_L g1330 ( .A(n_493), .Y(n_1330) );
INVx2_ASAP7_75t_SL g1385 ( .A(n_494), .Y(n_1385) );
AND2x4_ASAP7_75t_L g621 ( .A(n_495), .B(n_622), .Y(n_621) );
OAI33xp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_499), .A3(n_504), .B1(n_510), .B2(n_519), .B3(n_526), .Y(n_496) );
OAI33xp33_ASAP7_75t_L g1358 ( .A1(n_497), .A2(n_1359), .A3(n_1364), .B1(n_1367), .B2(n_1373), .B3(n_1376), .Y(n_1358) );
OAI22xp33_ASAP7_75t_L g519 ( .A1(n_500), .A2(n_520), .B1(n_521), .B2(n_525), .Y(n_519) );
BUFx2_ASAP7_75t_L g708 ( .A(n_500), .Y(n_708) );
INVx1_ASAP7_75t_L g754 ( .A(n_500), .Y(n_754) );
INVx1_ASAP7_75t_L g778 ( .A(n_500), .Y(n_778) );
OAI221xp5_ASAP7_75t_L g1116 ( .A1(n_500), .A2(n_523), .B1(n_709), .B2(n_1091), .C(n_1094), .Y(n_1116) );
OAI221xp5_ASAP7_75t_L g775 ( .A1(n_501), .A2(n_709), .B1(n_776), .B2(n_777), .C(n_779), .Y(n_775) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_503), .B(n_566), .Y(n_565) );
OR2x6_ASAP7_75t_L g712 ( .A(n_503), .B(n_572), .Y(n_712) );
OR2x2_ASAP7_75t_L g949 ( .A(n_503), .B(n_572), .Y(n_949) );
HB1xp67_ASAP7_75t_L g1363 ( .A(n_503), .Y(n_1363) );
OAI221xp5_ASAP7_75t_L g1118 ( .A1(n_505), .A2(n_1119), .B1(n_1120), .B2(n_1122), .C(n_1123), .Y(n_1118) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g1001 ( .A(n_507), .Y(n_1001) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g583 ( .A(n_508), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g720 ( .A(n_509), .Y(n_720) );
INVx2_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g889 ( .A(n_512), .Y(n_889) );
INVx2_ASAP7_75t_L g900 ( .A(n_512), .Y(n_900) );
INVx2_ASAP7_75t_L g952 ( .A(n_512), .Y(n_952) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g701 ( .A(n_513), .Y(n_701) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g773 ( .A(n_516), .Y(n_773) );
INVx2_ASAP7_75t_L g892 ( .A(n_516), .Y(n_892) );
INVx2_ASAP7_75t_L g1121 ( .A(n_516), .Y(n_1121) );
INVx2_ASAP7_75t_L g1371 ( .A(n_516), .Y(n_1371) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx3_ASAP7_75t_L g544 ( .A(n_517), .Y(n_544) );
INVx3_ASAP7_75t_L g1222 ( .A(n_517), .Y(n_1222) );
OAI221xp5_ASAP7_75t_L g1160 ( .A1(n_521), .A2(n_756), .B1(n_1161), .B2(n_1162), .C(n_1164), .Y(n_1160) );
OAI22xp33_ASAP7_75t_L g1373 ( .A1(n_521), .A2(n_1361), .B1(n_1374), .B2(n_1375), .Y(n_1373) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g751 ( .A(n_522), .Y(n_751) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx3_ASAP7_75t_L g895 ( .A(n_523), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_523), .B(n_1271), .Y(n_1270) );
BUFx3_ASAP7_75t_L g1437 ( .A(n_523), .Y(n_1437) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AOI33xp33_ASAP7_75t_L g1051 ( .A1(n_527), .A2(n_1052), .A3(n_1053), .B1(n_1056), .B2(n_1058), .B3(n_1059), .Y(n_1051) );
AOI33xp33_ASAP7_75t_L g1308 ( .A1(n_527), .A2(n_1309), .A3(n_1310), .B1(n_1311), .B2(n_1313), .B3(n_1318), .Y(n_1308) );
AOI33xp33_ASAP7_75t_L g1792 ( .A1(n_527), .A2(n_1052), .A3(n_1793), .B1(n_1794), .B2(n_1796), .B3(n_1798), .Y(n_1792) );
INVx6_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx5_ASAP7_75t_L g997 ( .A(n_528), .Y(n_997) );
OR2x6_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
NAND2x1p5_ASAP7_75t_L g620 ( .A(n_529), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g637 ( .A(n_530), .B(n_638), .Y(n_637) );
AND2x4_ASAP7_75t_L g1340 ( .A(n_530), .B(n_578), .Y(n_1340) );
BUFx2_ASAP7_75t_L g561 ( .A(n_531), .Y(n_561) );
INVx2_ASAP7_75t_L g758 ( .A(n_531), .Y(n_758) );
NAND4xp25_ASAP7_75t_L g536 ( .A(n_537), .B(n_594), .C(n_632), .D(n_644), .Y(n_536) );
OAI31xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_575), .A3(n_586), .B(n_592), .Y(n_537) );
OAI221xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_546), .B1(n_552), .B2(n_556), .C(n_562), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_542), .B1(n_543), .B2(n_545), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_540), .A2(n_553), .B1(n_554), .B2(n_555), .Y(n_552) );
BUFx2_ASAP7_75t_L g760 ( .A(n_540), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g1265 ( .A1(n_540), .A2(n_554), .B1(n_1266), .B2(n_1267), .Y(n_1265) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g1112 ( .A(n_541), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_542), .A2(n_545), .B1(n_602), .B2(n_604), .Y(n_601) );
INVx2_ASAP7_75t_SL g1169 ( .A(n_543), .Y(n_1169) );
INVx2_ASAP7_75t_L g1797 ( .A(n_543), .Y(n_1797) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g554 ( .A(n_544), .Y(n_554) );
INVx1_ASAP7_75t_L g705 ( .A(n_544), .Y(n_705) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_544), .Y(n_816) );
INVx2_ASAP7_75t_L g1115 ( .A(n_544), .Y(n_1115) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B(n_549), .Y(n_546) );
OAI221xp5_ASAP7_75t_L g945 ( .A1(n_548), .A2(n_709), .B1(n_924), .B2(n_925), .C(n_946), .Y(n_945) );
OAI221xp5_ASAP7_75t_L g1156 ( .A1(n_548), .A2(n_709), .B1(n_1138), .B2(n_1139), .C(n_1157), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_550), .B(n_692), .Y(n_691) );
BUFx2_ASAP7_75t_L g723 ( .A(n_550), .Y(n_723) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g560 ( .A(n_551), .Y(n_560) );
INVx2_ASAP7_75t_SL g897 ( .A(n_551), .Y(n_897) );
AOI222xp33_ASAP7_75t_L g632 ( .A1(n_553), .A2(n_563), .B1(n_633), .B2(n_639), .C1(n_640), .C2(n_642), .Y(n_632) );
INVx1_ASAP7_75t_L g944 ( .A(n_554), .Y(n_944) );
INVx2_ASAP7_75t_L g995 ( .A(n_554), .Y(n_995) );
INVx1_ASAP7_75t_L g1795 ( .A(n_554), .Y(n_1795) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_555), .A2(n_557), .B1(n_645), .B2(n_648), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_559), .Y(n_556) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_558), .A2(n_663), .B1(n_664), .B2(n_708), .C(n_709), .Y(n_707) );
OAI21xp5_ASAP7_75t_SL g1448 ( .A1(n_558), .A2(n_1449), .B(n_1450), .Y(n_1448) );
BUFx3_ASAP7_75t_L g1060 ( .A(n_560), .Y(n_1060) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B(n_565), .C(n_571), .Y(n_562) );
INVx1_ASAP7_75t_L g1320 ( .A(n_564), .Y(n_1320) );
NAND2x1p5_ASAP7_75t_L g1355 ( .A(n_569), .B(n_1352), .Y(n_1355) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x6_ASAP7_75t_L g732 ( .A(n_570), .B(n_572), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g1268 ( .A1(n_571), .A2(n_1216), .B(n_1269), .C(n_1270), .Y(n_1268) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g692 ( .A(n_572), .Y(n_692) );
INVx1_ASAP7_75t_L g826 ( .A(n_572), .Y(n_826) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx3_ASAP7_75t_L g695 ( .A(n_577), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_577), .A2(n_583), .B1(n_828), .B2(n_829), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_577), .A2(n_583), .B1(n_1256), .B2(n_1257), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_577), .A2(n_583), .B1(n_1431), .B2(n_1432), .Y(n_1430) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx2_ASAP7_75t_L g585 ( .A(n_578), .Y(n_585) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_579), .Y(n_815) );
INVx1_ASAP7_75t_L g994 ( .A(n_579), .Y(n_994) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_579), .Y(n_1000) );
BUFx2_ASAP7_75t_L g1057 ( .A(n_579), .Y(n_1057) );
BUFx6f_ASAP7_75t_L g1260 ( .A(n_579), .Y(n_1260) );
BUFx6f_ASAP7_75t_L g1316 ( .A(n_579), .Y(n_1316) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g696 ( .A(n_583), .Y(n_696) );
AND2x4_ASAP7_75t_L g590 ( .A(n_584), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
CKINVDCx6p67_ASAP7_75t_R g587 ( .A(n_588), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_588), .A2(n_831), .B1(n_832), .B2(n_833), .C(n_834), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g1258 ( .A1(n_588), .A2(n_1259), .B1(n_1261), .B2(n_1262), .Y(n_1258) );
AOI222xp33_ASAP7_75t_L g1425 ( .A1(n_588), .A2(n_590), .B1(n_1426), .B2(n_1427), .C1(n_1428), .C2(n_1429), .Y(n_1425) );
INVx8_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI221xp5_ASAP7_75t_SL g813 ( .A1(n_590), .A2(n_814), .B1(n_817), .B2(n_821), .C(n_822), .Y(n_813) );
INVx1_ASAP7_75t_L g820 ( .A(n_591), .Y(n_820) );
INVx1_ASAP7_75t_L g835 ( .A(n_592), .Y(n_835) );
OAI31xp33_ASAP7_75t_L g1107 ( .A1(n_592), .A2(n_1108), .A3(n_1109), .B(n_1117), .Y(n_1107) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NOR2xp67_ASAP7_75t_L g690 ( .A(n_593), .B(n_691), .Y(n_690) );
INVx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g845 ( .A(n_597), .Y(n_845) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_600), .Y(n_609) );
INVx2_ASAP7_75t_L g794 ( .A(n_600), .Y(n_794) );
INVx2_ASAP7_75t_L g980 ( .A(n_600), .Y(n_980) );
INVx2_ASAP7_75t_L g1071 ( .A(n_600), .Y(n_1071) );
INVx1_ASAP7_75t_L g1231 ( .A(n_600), .Y(n_1231) );
INVx2_ASAP7_75t_SL g1248 ( .A(n_600), .Y(n_1248) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_602), .A2(n_930), .B1(n_931), .B2(n_932), .Y(n_929) );
INVx1_ASAP7_75t_L g1064 ( .A(n_602), .Y(n_1064) );
INVx1_ASAP7_75t_L g1402 ( .A(n_602), .Y(n_1402) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g1388 ( .A(n_603), .Y(n_1388) );
AND2x4_ASAP7_75t_L g1390 ( .A(n_603), .B(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1065 ( .A(n_604), .Y(n_1065) );
INVx1_ASAP7_75t_L g1075 ( .A(n_604), .Y(n_1075) );
INVx1_ASAP7_75t_L g1102 ( .A(n_604), .Y(n_1102) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_606), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g1062 ( .A(n_606), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1462 ( .A1(n_606), .A2(n_874), .B1(n_1463), .B2(n_1469), .Y(n_1462) );
INVx4_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g1008 ( .A(n_609), .Y(n_1008) );
INVx2_ASAP7_75t_SL g791 ( .A(n_612), .Y(n_791) );
INVx1_ASAP7_75t_L g990 ( .A(n_612), .Y(n_990) );
INVx1_ASAP7_75t_L g1011 ( .A(n_612), .Y(n_1011) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx2_ASAP7_75t_L g1389 ( .A(n_613), .Y(n_1389) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_616), .Y(n_686) );
INVx1_ASAP7_75t_L g785 ( .A(n_616), .Y(n_785) );
INVx2_ASAP7_75t_L g856 ( .A(n_616), .Y(n_856) );
NAND2x1p5_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g1395 ( .A(n_618), .Y(n_1395) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
OR2x6_ASAP7_75t_L g625 ( .A(n_620), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g631 ( .A(n_620), .Y(n_631) );
OR2x2_ASAP7_75t_L g884 ( .A(n_620), .B(n_626), .Y(n_884) );
AND2x4_ASAP7_75t_L g1394 ( .A(n_621), .B(n_1395), .Y(n_1394) );
INVx1_ASAP7_75t_L g1397 ( .A(n_621), .Y(n_1397) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g786 ( .A(n_625), .Y(n_786) );
OR2x2_ASAP7_75t_L g1396 ( .A(n_626), .B(n_1397), .Y(n_1396) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g804 ( .A(n_628), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
BUFx2_ASAP7_75t_SL g1403 ( .A(n_629), .Y(n_1403) );
HB1xp67_ASAP7_75t_L g1468 ( .A(n_629), .Y(n_1468) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_SL g796 ( .A(n_630), .Y(n_796) );
BUFx3_ASAP7_75t_L g1068 ( .A(n_630), .Y(n_1068) );
BUFx4f_ASAP7_75t_L g1244 ( .A(n_630), .Y(n_1244) );
AND2x4_ASAP7_75t_L g1400 ( .A(n_630), .B(n_1391), .Y(n_1400) );
INVx1_ASAP7_75t_L g1459 ( .A(n_630), .Y(n_1459) );
INVx1_ASAP7_75t_L g1805 ( .A(n_630), .Y(n_1805) );
AND2x2_ASAP7_75t_L g655 ( .A(n_631), .B(n_656), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_633), .A2(n_640), .B1(n_755), .B2(n_761), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g851 ( .A1(n_633), .A2(n_640), .B1(n_852), .B2(n_853), .Y(n_851) );
AOI222xp33_ASAP7_75t_L g1272 ( .A1(n_633), .A2(n_642), .B1(n_645), .B2(n_1266), .C1(n_1269), .C2(n_1273), .Y(n_1272) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx2_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g1067 ( .A(n_635), .Y(n_1067) );
AND2x2_ASAP7_75t_L g640 ( .A(n_636), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OR2x6_ASAP7_75t_L g646 ( .A(n_637), .B(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g736 ( .A(n_637), .B(n_647), .Y(n_736) );
OR2x2_ASAP7_75t_L g738 ( .A(n_637), .B(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g740 ( .A(n_637), .B(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g1391 ( .A(n_638), .Y(n_1391) );
AOI22xp5_ASAP7_75t_L g1274 ( .A1(n_640), .A2(n_648), .B1(n_1267), .B2(n_1275), .Y(n_1274) );
OR2x6_ASAP7_75t_L g689 ( .A(n_642), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g1417 ( .A(n_642), .Y(n_1417) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_645), .A2(n_648), .B1(n_752), .B2(n_764), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_645), .A2(n_648), .B1(n_849), .B2(n_850), .Y(n_848) );
CKINVDCx6p67_ASAP7_75t_R g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g842 ( .A(n_647), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g1143 ( .A1(n_647), .A2(n_1086), .B1(n_1144), .B2(n_1145), .Y(n_1143) );
CKINVDCx6p67_ASAP7_75t_R g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND4x1_ASAP7_75t_L g652 ( .A(n_653), .B(n_687), .C(n_693), .D(n_734), .Y(n_652) );
NOR3xp33_ASAP7_75t_SL g653 ( .A(n_654), .B(n_658), .C(n_685), .Y(n_653) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g854 ( .A1(n_655), .A2(n_786), .B1(n_855), .B2(n_856), .C(n_857), .Y(n_854) );
NOR3xp33_ASAP7_75t_SL g865 ( .A(n_655), .B(n_866), .C(n_882), .Y(n_865) );
NOR3xp33_ASAP7_75t_SL g917 ( .A(n_655), .B(n_918), .C(n_933), .Y(n_917) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_655), .Y(n_1083) );
AOI221xp5_ASAP7_75t_L g1250 ( .A1(n_655), .A2(n_786), .B1(n_856), .B2(n_1251), .C(n_1252), .Y(n_1250) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B1(n_664), .B2(n_665), .C(n_668), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g1463 ( .A1(n_660), .A2(n_1442), .B1(n_1464), .B2(n_1465), .C(n_1466), .Y(n_1463) );
BUFx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g1469 ( .A1(n_661), .A2(n_677), .B1(n_1428), .B2(n_1429), .C(n_1470), .Y(n_1469) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g870 ( .A(n_667), .Y(n_870) );
BUFx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g741 ( .A(n_670), .Y(n_741) );
BUFx4f_ASAP7_75t_L g790 ( .A(n_670), .Y(n_790) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI22xp33_ASAP7_75t_L g1134 ( .A1(n_672), .A2(n_682), .B1(n_1135), .B2(n_1136), .Y(n_1134) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_673), .Y(n_684) );
INVx1_ASAP7_75t_L g921 ( .A(n_673), .Y(n_921) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_677), .B2(n_679), .C(n_680), .Y(n_674) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g919 ( .A1(n_682), .A2(n_920), .B1(n_921), .B2(n_922), .Y(n_919) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g1099 ( .A(n_683), .Y(n_1099) );
BUFx3_ASAP7_75t_L g1323 ( .A(n_683), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_689), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g811 ( .A(n_689), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_689), .B(n_864), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_689), .B(n_938), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_689), .B(n_1106), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_689), .B(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1427 ( .A(n_691), .Y(n_1427) );
AND2x2_ASAP7_75t_L g728 ( .A(n_692), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g958 ( .A(n_692), .B(n_729), .Y(n_958) );
OAI31xp33_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_697), .A3(n_713), .B(n_733), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_702), .B1(n_703), .B2(n_706), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g715 ( .A(n_700), .Y(n_715) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx2_ASAP7_75t_L g770 ( .A(n_701), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g1364 ( .A1(n_703), .A2(n_952), .B1(n_1365), .B2(n_1366), .Y(n_1364) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g834 ( .A(n_712), .Y(n_834) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_717), .B2(n_721), .C(n_722), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_SL g1016 ( .A(n_725), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_730), .B2(n_731), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_728), .A2(n_731), .B1(n_766), .B2(n_767), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_728), .A2(n_731), .B1(n_907), .B2(n_908), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_728), .A2(n_731), .B1(n_1125), .B2(n_1126), .Y(n_1124) );
AOI22xp5_ASAP7_75t_L g1443 ( .A1(n_728), .A2(n_731), .B1(n_1444), .B2(n_1445), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_731), .A2(n_957), .B1(n_958), .B2(n_959), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_731), .A2(n_958), .B1(n_1171), .B2(n_1172), .Y(n_1170) );
CKINVDCx11_ASAP7_75t_R g731 ( .A(n_732), .Y(n_731) );
CKINVDCx8_ASAP7_75t_R g961 ( .A(n_733), .Y(n_961) );
AOI221x1_ASAP7_75t_SL g1423 ( .A1(n_733), .A2(n_1198), .B1(n_1424), .B2(n_1451), .C(n_1462), .Y(n_1423) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_737), .Y(n_734) );
XNOR2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_860), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B1(n_808), .B2(n_859), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NAND3xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_780), .C(n_782), .Y(n_746) );
OAI221xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_752), .B1(n_753), .B2(n_755), .C(n_756), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_762), .B2(n_764), .Y(n_759) );
INVx2_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVx4_ASAP7_75t_L g902 ( .A(n_763), .Y(n_902) );
BUFx3_ASAP7_75t_L g1317 ( .A(n_763), .Y(n_1317) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_766), .A2(n_767), .B1(n_785), .B2(n_786), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B1(n_772), .B2(n_774), .Y(n_769) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NOR2xp33_ASAP7_75t_SL g782 ( .A(n_783), .B(n_805), .Y(n_782) );
NAND3xp33_ASAP7_75t_SL g783 ( .A(n_784), .B(n_787), .C(n_803), .Y(n_783) );
AOI33xp33_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_789), .A3(n_792), .B1(n_797), .B2(n_798), .B3(n_800), .Y(n_787) );
INVx1_ASAP7_75t_L g1088 ( .A(n_791), .Y(n_1088) );
BUFx6f_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g1035 ( .A(n_796), .Y(n_1035) );
NAND3xp33_ASAP7_75t_L g1229 ( .A(n_800), .B(n_1230), .C(n_1232), .Y(n_1229) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
AOI33xp33_ASAP7_75t_L g837 ( .A1(n_802), .A2(n_838), .A3(n_841), .B1(n_843), .B2(n_846), .B3(n_847), .Y(n_837) );
NAND3xp33_ASAP7_75t_L g1006 ( .A(n_802), .B(n_1007), .C(n_1009), .Y(n_1006) );
AOI33xp33_ASAP7_75t_L g1240 ( .A1(n_802), .A2(n_1241), .A3(n_1242), .B1(n_1243), .B2(n_1245), .B3(n_1249), .Y(n_1240) );
NAND3xp33_ASAP7_75t_L g1510 ( .A(n_802), .B(n_1511), .C(n_1512), .Y(n_1510) );
AOI33xp33_ASAP7_75t_L g1800 ( .A1(n_802), .A2(n_1241), .A3(n_1801), .B1(n_1802), .B2(n_1803), .B3(n_1806), .Y(n_1800) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx2_ASAP7_75t_L g859 ( .A(n_808), .Y(n_859) );
XOR2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_858), .Y(n_808) );
NOR3xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_812), .C(n_836), .Y(n_809) );
AOI31xp33_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_827), .A3(n_830), .B(n_835), .Y(n_812) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g1224 ( .A(n_820), .Y(n_1224) );
NAND2x1p5_ASAP7_75t_L g823 ( .A(n_824), .B(n_826), .Y(n_823) );
NAND2x1_ASAP7_75t_SL g1351 ( .A(n_824), .B(n_1352), .Y(n_1351) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
NOR3xp33_ASAP7_75t_L g1433 ( .A(n_834), .B(n_1434), .C(n_1446), .Y(n_1433) );
AOI22xp33_ASAP7_75t_L g1377 ( .A1(n_835), .A2(n_1378), .B1(n_1413), .B2(n_1414), .Y(n_1377) );
NAND4xp25_ASAP7_75t_L g836 ( .A(n_837), .B(n_848), .C(n_851), .D(n_854), .Y(n_836) );
NAND3xp33_ASAP7_75t_L g987 ( .A(n_838), .B(n_988), .C(n_989), .Y(n_987) );
NAND3xp33_ASAP7_75t_L g1225 ( .A(n_838), .B(n_1226), .C(n_1227), .Y(n_1225) );
NAND3xp33_ASAP7_75t_L g1507 ( .A(n_838), .B(n_1508), .C(n_1509), .Y(n_1507) );
INVx3_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g883 ( .A(n_856), .Y(n_883) );
AO22x2_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_914), .B1(n_915), .B2(n_962), .Y(n_860) );
INVx1_ASAP7_75t_L g962 ( .A(n_861), .Y(n_962) );
AND4x1_ASAP7_75t_L g862 ( .A(n_863), .B(n_865), .C(n_885), .D(n_911), .Y(n_862) );
OAI221xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_869), .B1(n_870), .B2(n_871), .C(n_872), .Y(n_867) );
OAI22xp33_ASAP7_75t_L g1090 ( .A1(n_868), .A2(n_1091), .B1(n_1092), .B2(n_1094), .Y(n_1090) );
OAI21xp33_ASAP7_75t_L g894 ( .A1(n_871), .A2(n_895), .B(n_896), .Y(n_894) );
INVx2_ASAP7_75t_SL g931 ( .A(n_873), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_875), .Y(n_874) );
INVx2_ASAP7_75t_SL g1086 ( .A(n_880), .Y(n_1086) );
OAI31xp33_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_887), .A3(n_898), .B(n_909), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_890), .B1(n_891), .B2(n_893), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_889), .A2(n_920), .B1(n_922), .B2(n_943), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g1152 ( .A1(n_889), .A2(n_1135), .B1(n_1136), .B2(n_1153), .Y(n_1152) );
OAI22xp5_ASAP7_75t_SL g1165 ( .A1(n_889), .A2(n_1166), .B1(n_1167), .B2(n_1168), .Y(n_1165) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
AND2x4_ASAP7_75t_L g1345 ( .A(n_897), .B(n_1340), .Y(n_1345) );
OAI221xp5_ASAP7_75t_L g899 ( .A1(n_900), .A2(n_901), .B1(n_902), .B2(n_903), .C(n_904), .Y(n_899) );
OAI221xp5_ASAP7_75t_L g951 ( .A1(n_902), .A2(n_952), .B1(n_953), .B2(n_954), .C(n_955), .Y(n_951) );
INVx2_ASAP7_75t_SL g1312 ( .A(n_902), .Y(n_1312) );
INVx2_ASAP7_75t_L g1447 ( .A(n_902), .Y(n_1447) );
AND2x6_ASAP7_75t_L g1342 ( .A(n_905), .B(n_1340), .Y(n_1342) );
NAND2x1p5_ASAP7_75t_L g1357 ( .A(n_905), .B(n_1352), .Y(n_1357) );
OAI21xp5_ASAP7_75t_L g1253 ( .A1(n_909), .A2(n_1254), .B(n_1263), .Y(n_1253) );
BUFx8_ASAP7_75t_SL g909 ( .A(n_910), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .Y(n_911) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
AND4x1_ASAP7_75t_L g916 ( .A(n_917), .B(n_934), .C(n_937), .D(n_939), .Y(n_916) );
NOR2xp33_ASAP7_75t_L g934 ( .A(n_935), .B(n_936), .Y(n_934) );
OAI31xp33_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_941), .A3(n_950), .B(n_960), .Y(n_939) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx2_ASAP7_75t_SL g946 ( .A(n_947), .Y(n_946) );
INVx2_ASAP7_75t_SL g947 ( .A(n_948), .Y(n_947) );
OAI31xp33_ASAP7_75t_L g1149 ( .A1(n_960), .A2(n_1150), .A3(n_1151), .B(n_1159), .Y(n_1149) );
INVx2_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
XNOR2x1_ASAP7_75t_L g963 ( .A(n_964), .B(n_1177), .Y(n_963) );
XNOR2xp5_ASAP7_75t_L g964 ( .A(n_965), .B(n_1078), .Y(n_964) );
XNOR2x1_ASAP7_75t_L g965 ( .A(n_966), .B(n_1029), .Y(n_965) );
AO211x2_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_969), .B(n_986), .C(n_1012), .Y(n_967) );
BUFx6f_ASAP7_75t_L g1198 ( .A(n_968), .Y(n_1198) );
NAND3xp33_ASAP7_75t_L g969 ( .A(n_970), .B(n_977), .C(n_982), .Y(n_969) );
INVx1_ASAP7_75t_L g1293 ( .A(n_974), .Y(n_1293) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
BUFx4f_ASAP7_75t_L g1460 ( .A(n_975), .Y(n_1460) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_979), .A2(n_984), .B1(n_1285), .B2(n_1286), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1452 ( .A1(n_979), .A2(n_984), .B1(n_1453), .B2(n_1454), .Y(n_1452) );
CKINVDCx6p67_ASAP7_75t_R g1040 ( .A(n_984), .Y(n_1040) );
NAND4xp25_ASAP7_75t_L g986 ( .A(n_987), .B(n_991), .C(n_998), .D(n_1006), .Y(n_986) );
NAND3xp33_ASAP7_75t_L g991 ( .A(n_992), .B(n_996), .C(n_997), .Y(n_991) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
NAND3xp33_ASAP7_75t_L g1214 ( .A(n_997), .B(n_1215), .C(n_1217), .Y(n_1214) );
CKINVDCx8_ASAP7_75t_R g1376 ( .A(n_997), .Y(n_1376) );
NAND3xp33_ASAP7_75t_L g1504 ( .A(n_997), .B(n_1505), .C(n_1506), .Y(n_1504) );
NAND3xp33_ASAP7_75t_L g998 ( .A(n_999), .B(n_1002), .C(n_1005), .Y(n_998) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
INVx2_ASAP7_75t_SL g1055 ( .A(n_1004), .Y(n_1055) );
BUFx2_ASAP7_75t_L g1799 ( .A(n_1004), .Y(n_1799) );
BUFx3_ASAP7_75t_L g1309 ( .A(n_1005), .Y(n_1309) );
AOI31xp33_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1020), .A3(n_1024), .B(n_1028), .Y(n_1012) );
INVx2_ASAP7_75t_SL g1015 ( .A(n_1016), .Y(n_1015) );
INVx2_ASAP7_75t_L g1206 ( .A(n_1016), .Y(n_1206) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1018), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_1021), .A2(n_1201), .B1(n_1202), .B2(n_1203), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_1021), .A2(n_1203), .B1(n_1302), .B2(n_1303), .Y(n_1301) );
AOI22xp33_ASAP7_75t_L g1488 ( .A1(n_1021), .A2(n_1203), .B1(n_1489), .B2(n_1490), .Y(n_1488) );
AOI22xp5_ASAP7_75t_L g1781 ( .A1(n_1021), .A2(n_1203), .B1(n_1782), .B2(n_1783), .Y(n_1781) );
INVx5_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx4_ASAP7_75t_L g1306 ( .A(n_1027), .Y(n_1306) );
AO21x1_ASAP7_75t_SL g1042 ( .A1(n_1028), .A2(n_1043), .B(n_1048), .Y(n_1042) );
CKINVDCx16_ASAP7_75t_R g1212 ( .A(n_1028), .Y(n_1212) );
AOI31xp33_ASAP7_75t_L g1296 ( .A1(n_1028), .A2(n_1297), .A3(n_1301), .B(n_1304), .Y(n_1296) );
AND4x1_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1042), .C(n_1051), .D(n_1061), .Y(n_1030) );
NAND4xp25_ASAP7_75t_L g1077 ( .A(n_1031), .B(n_1042), .C(n_1051), .D(n_1061), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1035), .Y(n_1033) );
NAND3xp33_ASAP7_75t_L g1218 ( .A(n_1052), .B(n_1219), .C(n_1223), .Y(n_1218) );
NAND3xp33_ASAP7_75t_L g1501 ( .A(n_1052), .B(n_1502), .C(n_1503), .Y(n_1501) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
AOI33xp33_ASAP7_75t_L g1321 ( .A1(n_1062), .A2(n_1322), .A3(n_1326), .B1(n_1328), .B2(n_1329), .B3(n_1330), .Y(n_1321) );
HB1xp67_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
BUFx3_ASAP7_75t_L g1327 ( .A(n_1071), .Y(n_1327) );
BUFx6f_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1073), .Y(n_1382) );
AND2x4_ASAP7_75t_L g1406 ( .A(n_1073), .B(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1075), .Y(n_1465) );
AOI22xp5_ASAP7_75t_L g1078 ( .A1(n_1079), .A2(n_1080), .B1(n_1130), .B2(n_1176), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
AND4x1_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1105), .C(n_1107), .D(n_1127), .Y(n_1081) );
NOR3xp33_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1084), .C(n_1104), .Y(n_1082) );
NOR3xp33_ASAP7_75t_SL g1132 ( .A(n_1083), .B(n_1133), .C(n_1146), .Y(n_1132) );
OAI22xp33_ASAP7_75t_L g1085 ( .A1(n_1086), .A2(n_1087), .B1(n_1088), .B2(n_1089), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_1087), .A2(n_1089), .B1(n_1111), .B2(n_1113), .Y(n_1110) );
HB1xp67_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1093), .Y(n_1191) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_1099), .A2(n_1100), .B1(n_1101), .B2(n_1103), .Y(n_1098) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1129), .Y(n_1127) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1130), .Y(n_1176) );
AND4x1_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1147), .C(n_1149), .D(n_1173), .Y(n_1131) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
BUFx2_ASAP7_75t_L g1361 ( .A(n_1157), .Y(n_1361) );
INVx2_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
NOR2xp33_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1175), .Y(n_1173) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
OAI22x1_ASAP7_75t_L g1179 ( .A1(n_1180), .A2(n_1181), .B1(n_1235), .B2(n_1236), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1183), .Y(n_1234) );
AOI221x1_ASAP7_75t_L g1183 ( .A1(n_1184), .A2(n_1198), .B1(n_1199), .B2(n_1212), .C(n_1213), .Y(n_1183) );
NAND3xp33_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1192), .C(n_1195), .Y(n_1184) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1188), .Y(n_1484) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
AOI211x1_ASAP7_75t_L g1282 ( .A1(n_1198), .A2(n_1283), .B(n_1296), .C(n_1307), .Y(n_1282) );
AOI221x1_ASAP7_75t_L g1475 ( .A1(n_1198), .A2(n_1212), .B1(n_1476), .B2(n_1487), .C(n_1500), .Y(n_1475) );
AOI211xp5_ASAP7_75t_L g1779 ( .A1(n_1212), .A2(n_1780), .B(n_1791), .C(n_1807), .Y(n_1779) );
NAND4xp25_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1218), .C(n_1225), .D(n_1229), .Y(n_1213) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
INVx2_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
AND2x4_ASAP7_75t_L g1339 ( .A(n_1222), .B(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1222), .Y(n_1441) );
INVx2_ASAP7_75t_SL g1235 ( .A(n_1236), .Y(n_1235) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
NAND4xp75_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1253), .C(n_1272), .D(n_1274), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1250), .Y(n_1239) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1258), .Y(n_1254) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
XOR2xp5_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1419), .Y(n_1278) );
AOI22xp5_ASAP7_75t_L g1279 ( .A1(n_1280), .A2(n_1281), .B1(n_1331), .B2(n_1418), .Y(n_1279) );
INVx2_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
NAND4xp25_ASAP7_75t_SL g1283 ( .A(n_1284), .B(n_1287), .C(n_1290), .D(n_1295), .Y(n_1283) );
BUFx2_ASAP7_75t_L g1461 ( .A(n_1295), .Y(n_1461) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1321), .Y(n_1307) );
INVx3_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx2_ASAP7_75t_SL g1315 ( .A(n_1316), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1316), .B(n_1340), .Y(n_1347) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1331), .Y(n_1418) );
HB1xp67_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1377), .Y(n_1333) );
NOR3xp33_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1348), .C(n_1358), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1343), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_1337), .A2(n_1338), .B1(n_1341), .B2(n_1342), .Y(n_1336) );
BUFx2_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g1343 ( .A1(n_1344), .A2(n_1345), .B1(n_1346), .B2(n_1347), .Y(n_1343) );
INVx2_ASAP7_75t_SL g1349 ( .A(n_1350), .Y(n_1349) );
INVx2_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx3_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
BUFx4f_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
BUFx2_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
OAI22xp33_ASAP7_75t_L g1359 ( .A1(n_1360), .A2(n_1361), .B1(n_1362), .B2(n_1363), .Y(n_1359) );
OAI22xp5_ASAP7_75t_L g1367 ( .A1(n_1368), .A2(n_1369), .B1(n_1370), .B2(n_1372), .Y(n_1367) );
OAI22xp5_ASAP7_75t_L g1439 ( .A1(n_1368), .A2(n_1440), .B1(n_1441), .B2(n_1442), .Y(n_1439) );
AOI221xp5_ASAP7_75t_L g1379 ( .A1(n_1369), .A2(n_1380), .B1(n_1386), .B2(n_1390), .C(n_1392), .Y(n_1379) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_1372), .A2(n_1374), .B1(n_1409), .B2(n_1411), .Y(n_1408) );
AOI221xp5_ASAP7_75t_L g1398 ( .A1(n_1375), .A2(n_1399), .B1(n_1401), .B2(n_1405), .C(n_1406), .Y(n_1398) );
NAND3xp33_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1398), .C(n_1408), .Y(n_1378) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
INVx2_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_SL g1407 ( .A(n_1397), .Y(n_1407) );
BUFx6f_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
INVx6_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
INVx4_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
INVx5_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
AND2x4_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1417), .Y(n_1415) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
AOI22xp5_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1422), .B1(n_1473), .B2(n_1515), .Y(n_1420) );
INVx2_ASAP7_75t_SL g1421 ( .A(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1423), .Y(n_1472) );
NAND3xp33_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1430), .C(n_1433), .Y(n_1424) );
OAI21xp5_ASAP7_75t_SL g1434 ( .A1(n_1435), .A2(n_1439), .B(n_1443), .Y(n_1434) );
OAI21xp5_ASAP7_75t_L g1435 ( .A1(n_1436), .A2(n_1437), .B(n_1438), .Y(n_1435) );
NAND4xp25_ASAP7_75t_SL g1451 ( .A(n_1452), .B(n_1455), .C(n_1457), .D(n_1461), .Y(n_1451) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
HB1xp67_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1474), .Y(n_1515) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1475), .Y(n_1514) );
NAND2xp5_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1480), .Y(n_1476) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
NAND4xp25_ASAP7_75t_L g1500 ( .A(n_1501), .B(n_1504), .C(n_1507), .D(n_1510), .Y(n_1500) );
OAI221xp5_ASAP7_75t_SL g1517 ( .A1(n_1518), .A2(n_1772), .B1(n_1775), .B2(n_1818), .C(n_1823), .Y(n_1517) );
NOR3xp33_ASAP7_75t_L g1518 ( .A(n_1519), .B(n_1683), .C(n_1729), .Y(n_1518) );
AOI21xp5_ASAP7_75t_L g1519 ( .A1(n_1520), .A2(n_1634), .B(n_1673), .Y(n_1519) );
AOI221xp5_ASAP7_75t_L g1520 ( .A1(n_1521), .A2(n_1567), .B1(n_1583), .B2(n_1589), .C(n_1597), .Y(n_1520) );
INVxp67_ASAP7_75t_SL g1521 ( .A(n_1522), .Y(n_1521) );
NAND2xp5_ASAP7_75t_L g1522 ( .A(n_1523), .B(n_1542), .Y(n_1522) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1523), .Y(n_1655) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1523), .Y(n_1691) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_1523), .B(n_1686), .Y(n_1702) );
HB1xp67_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
INVx2_ASAP7_75t_SL g1587 ( .A(n_1524), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1524), .B(n_1580), .Y(n_1632) );
OR2x2_ASAP7_75t_L g1639 ( .A(n_1524), .B(n_1580), .Y(n_1639) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1525), .Y(n_1577) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1525), .Y(n_1676) );
BUFx3_ASAP7_75t_L g1774 ( .A(n_1525), .Y(n_1774) );
AND2x4_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1529), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1526), .B(n_1529), .Y(n_1553) );
HB1xp67_ASAP7_75t_L g1837 ( .A(n_1526), .Y(n_1837) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
AND2x4_ASAP7_75t_L g1531 ( .A(n_1527), .B(n_1529), .Y(n_1531) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
NAND2xp5_ASAP7_75t_L g1537 ( .A(n_1528), .B(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1530), .Y(n_1538) );
INVx1_ASAP7_75t_SL g1562 ( .A(n_1531), .Y(n_1562) );
INVx2_ASAP7_75t_L g1595 ( .A(n_1531), .Y(n_1595) );
OAI22xp33_ASAP7_75t_L g1532 ( .A1(n_1533), .A2(n_1534), .B1(n_1539), .B2(n_1540), .Y(n_1532) );
OAI22xp5_ASAP7_75t_L g1564 ( .A1(n_1534), .A2(n_1540), .B1(n_1565), .B2(n_1566), .Y(n_1564) );
OAI22xp33_ASAP7_75t_L g1570 ( .A1(n_1534), .A2(n_1571), .B1(n_1572), .B2(n_1573), .Y(n_1570) );
BUFx3_ASAP7_75t_L g1680 ( .A(n_1534), .Y(n_1680) );
BUFx6f_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
OAI22xp5_ASAP7_75t_L g1555 ( .A1(n_1535), .A2(n_1540), .B1(n_1556), .B2(n_1557), .Y(n_1555) );
OR2x2_ASAP7_75t_L g1535 ( .A(n_1536), .B(n_1537), .Y(n_1535) );
OR2x2_ASAP7_75t_L g1540 ( .A(n_1536), .B(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1536), .Y(n_1549) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1537), .Y(n_1548) );
HB1xp67_ASAP7_75t_L g1836 ( .A(n_1538), .Y(n_1836) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1540), .Y(n_1574) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1541), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1558), .Y(n_1542) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_1543), .B(n_1590), .Y(n_1657) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1543), .B(n_1624), .Y(n_1669) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
NOR2xp33_ASAP7_75t_L g1616 ( .A(n_1544), .B(n_1601), .Y(n_1616) );
OR2x2_ASAP7_75t_L g1705 ( .A(n_1544), .B(n_1558), .Y(n_1705) );
OR2x2_ASAP7_75t_L g1754 ( .A(n_1544), .B(n_1591), .Y(n_1754) );
OR2x2_ASAP7_75t_L g1544 ( .A(n_1545), .B(n_1554), .Y(n_1544) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1545), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1545), .B(n_1558), .Y(n_1609) );
AND2x2_ASAP7_75t_L g1621 ( .A(n_1545), .B(n_1622), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1662 ( .A(n_1545), .B(n_1554), .Y(n_1662) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1546), .B(n_1552), .Y(n_1545) );
AND2x4_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1549), .Y(n_1547) );
AND2x4_ASAP7_75t_L g1550 ( .A(n_1549), .B(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1553), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1554), .B(n_1590), .Y(n_1589) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1554), .B(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1554), .Y(n_1622) );
NOR2xp33_ASAP7_75t_L g1735 ( .A(n_1554), .B(n_1596), .Y(n_1735) );
CKINVDCx6p67_ASAP7_75t_R g1596 ( .A(n_1558), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1615 ( .A(n_1558), .B(n_1616), .Y(n_1615) );
OAI331xp33_ASAP7_75t_L g1635 ( .A1(n_1558), .A2(n_1622), .A3(n_1636), .B1(n_1640), .B2(n_1643), .B3(n_1645), .C1(n_1647), .Y(n_1635) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_1558), .B(n_1621), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1558), .B(n_1603), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1718 ( .A(n_1558), .B(n_1604), .Y(n_1718) );
OR2x2_ASAP7_75t_L g1725 ( .A(n_1558), .B(n_1604), .Y(n_1725) );
OR2x6_ASAP7_75t_SL g1558 ( .A(n_1559), .B(n_1564), .Y(n_1558) );
OAI22xp5_ASAP7_75t_L g1559 ( .A1(n_1560), .A2(n_1561), .B1(n_1562), .B2(n_1563), .Y(n_1559) );
XNOR2xp5_ASAP7_75t_L g1778 ( .A(n_1561), .B(n_1779), .Y(n_1778) );
OAI22xp5_ASAP7_75t_L g1575 ( .A1(n_1562), .A2(n_1576), .B1(n_1577), .B2(n_1578), .Y(n_1575) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1567), .Y(n_1658) );
A2O1A1Ixp33_ASAP7_75t_SL g1761 ( .A1(n_1567), .A2(n_1744), .B(n_1762), .C(n_1763), .Y(n_1761) );
AND2x2_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1579), .Y(n_1567) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1568), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1568), .B(n_1611), .Y(n_1626) );
OR2x2_ASAP7_75t_L g1649 ( .A(n_1568), .B(n_1580), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1653 ( .A(n_1568), .B(n_1580), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1665 ( .A(n_1568), .B(n_1632), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1568), .B(n_1587), .Y(n_1685) );
NAND2xp5_ASAP7_75t_L g1720 ( .A(n_1568), .B(n_1673), .Y(n_1720) );
INVx3_ASAP7_75t_L g1749 ( .A(n_1568), .Y(n_1749) );
INVx3_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1569), .B(n_1580), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1646 ( .A(n_1569), .B(n_1591), .Y(n_1646) );
OR2x2_ASAP7_75t_L g1770 ( .A(n_1569), .B(n_1639), .Y(n_1770) );
OR2x2_ASAP7_75t_L g1569 ( .A(n_1570), .B(n_1575), .Y(n_1569) );
HB1xp67_ASAP7_75t_L g1682 ( .A(n_1573), .Y(n_1682) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
OAI211xp5_ASAP7_75t_SL g1597 ( .A1(n_1579), .A2(n_1598), .B(n_1605), .C(n_1627), .Y(n_1597) );
AOI22xp33_ASAP7_75t_SL g1738 ( .A1(n_1579), .A2(n_1704), .B1(n_1739), .B2(n_1743), .Y(n_1738) );
O2A1O1Ixp33_ASAP7_75t_L g1743 ( .A1(n_1579), .A2(n_1601), .B(n_1632), .C(n_1688), .Y(n_1743) );
INVx2_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
OR2x2_ASAP7_75t_L g1586 ( .A(n_1580), .B(n_1587), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1580), .B(n_1587), .Y(n_1644) );
OAI22xp5_ASAP7_75t_L g1689 ( .A1(n_1580), .A2(n_1625), .B1(n_1690), .B2(n_1692), .Y(n_1689) );
AND2x4_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1582), .Y(n_1580) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1584), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1584 ( .A(n_1585), .B(n_1588), .Y(n_1584) );
NAND2xp5_ASAP7_75t_L g1760 ( .A(n_1585), .B(n_1687), .Y(n_1760) );
INVx2_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
OR2x2_ASAP7_75t_L g1751 ( .A(n_1586), .B(n_1687), .Y(n_1751) );
INVx2_ASAP7_75t_SL g1611 ( .A(n_1587), .Y(n_1611) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1588), .B(n_1629), .Y(n_1628) );
NAND2xp5_ASAP7_75t_L g1618 ( .A(n_1590), .B(n_1603), .Y(n_1618) );
NAND2xp5_ASAP7_75t_L g1713 ( .A(n_1590), .B(n_1662), .Y(n_1713) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1596), .Y(n_1590) );
INVx4_ASAP7_75t_L g1601 ( .A(n_1591), .Y(n_1601) );
INVx2_ASAP7_75t_L g1608 ( .A(n_1591), .Y(n_1608) );
NOR2xp33_ASAP7_75t_L g1624 ( .A(n_1591), .B(n_1596), .Y(n_1624) );
NAND2xp5_ASAP7_75t_L g1694 ( .A(n_1591), .B(n_1662), .Y(n_1694) );
OR2x2_ASAP7_75t_L g1704 ( .A(n_1591), .B(n_1705), .Y(n_1704) );
AOI322xp5_ASAP7_75t_L g1708 ( .A1(n_1591), .A2(n_1632), .A3(n_1638), .B1(n_1644), .B2(n_1709), .C1(n_1712), .C2(n_1714), .Y(n_1708) );
AND2x2_ASAP7_75t_L g1737 ( .A(n_1591), .B(n_1644), .Y(n_1737) );
AND2x6_ASAP7_75t_L g1591 ( .A(n_1592), .B(n_1593), .Y(n_1591) );
INVx2_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
OAI22xp5_ASAP7_75t_L g1674 ( .A1(n_1595), .A2(n_1675), .B1(n_1676), .B2(n_1677), .Y(n_1674) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1596), .B(n_1603), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1633 ( .A(n_1596), .B(n_1621), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1596), .B(n_1661), .Y(n_1660) );
NOR2xp33_ASAP7_75t_L g1693 ( .A(n_1596), .B(n_1694), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1596), .B(n_1622), .Y(n_1740) );
OR2x2_ASAP7_75t_L g1765 ( .A(n_1596), .B(n_1622), .Y(n_1765) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1601), .B(n_1602), .Y(n_1600) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1601), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1637 ( .A(n_1601), .B(n_1638), .Y(n_1637) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1601), .B(n_1633), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1661 ( .A(n_1601), .B(n_1662), .Y(n_1661) );
NOR2xp33_ASAP7_75t_L g1741 ( .A(n_1601), .B(n_1742), .Y(n_1741) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1602), .B(n_1629), .Y(n_1707) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1603), .Y(n_1642) );
OAI22xp5_ASAP7_75t_SL g1756 ( .A1(n_1604), .A2(n_1757), .B1(n_1758), .B2(n_1760), .Y(n_1756) );
AOI211xp5_ASAP7_75t_L g1605 ( .A1(n_1606), .A2(n_1610), .B(n_1613), .C(n_1617), .Y(n_1605) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
NAND2xp5_ASAP7_75t_L g1607 ( .A(n_1608), .B(n_1609), .Y(n_1607) );
INVx2_ASAP7_75t_L g1687 ( .A(n_1608), .Y(n_1687) );
NAND2xp5_ASAP7_75t_L g1727 ( .A(n_1608), .B(n_1728), .Y(n_1727) );
OAI32xp33_ASAP7_75t_L g1739 ( .A1(n_1608), .A2(n_1632), .A3(n_1688), .B1(n_1740), .B2(n_1741), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1611), .B(n_1612), .Y(n_1610) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1611), .Y(n_1614) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1611), .Y(n_1629) );
NOR2xp33_ASAP7_75t_L g1716 ( .A(n_1611), .B(n_1717), .Y(n_1716) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1611), .Y(n_1728) );
OAI22xp5_ASAP7_75t_L g1752 ( .A1(n_1611), .A2(n_1688), .B1(n_1753), .B2(n_1755), .Y(n_1752) );
NAND2xp5_ASAP7_75t_L g1753 ( .A(n_1611), .B(n_1754), .Y(n_1753) );
OAI21xp33_ASAP7_75t_L g1700 ( .A1(n_1612), .A2(n_1701), .B(n_1703), .Y(n_1700) );
NOR2xp33_ASAP7_75t_L g1613 ( .A(n_1614), .B(n_1615), .Y(n_1613) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1615), .Y(n_1697) );
AOI21xp33_ASAP7_75t_SL g1617 ( .A1(n_1618), .A2(n_1619), .B(n_1625), .Y(n_1617) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1618), .Y(n_1755) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1619), .Y(n_1721) );
OR2x2_ASAP7_75t_L g1619 ( .A(n_1620), .B(n_1623), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1641 ( .A(n_1620), .B(n_1642), .Y(n_1641) );
NOR2xp33_ASAP7_75t_L g1663 ( .A(n_1620), .B(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1621), .Y(n_1620) );
NOR3xp33_ASAP7_75t_L g1767 ( .A(n_1622), .B(n_1687), .C(n_1768), .Y(n_1767) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1626), .Y(n_1625) );
OAI21xp5_ASAP7_75t_L g1627 ( .A1(n_1628), .A2(n_1630), .B(n_1633), .Y(n_1627) );
AOI221xp5_ASAP7_75t_SL g1715 ( .A1(n_1628), .A2(n_1716), .B1(n_1719), .B2(n_1721), .C(n_1722), .Y(n_1715) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1631), .B(n_1632), .Y(n_1630) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1633), .Y(n_1711) );
NOR5xp2_ASAP7_75t_L g1634 ( .A(n_1635), .B(n_1651), .C(n_1663), .D(n_1666), .E(n_1670), .Y(n_1634) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
A2O1A1Ixp33_ASAP7_75t_L g1771 ( .A1(n_1637), .A2(n_1670), .B(n_1735), .C(n_1749), .Y(n_1771) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
NOR2xp33_ASAP7_75t_L g1670 ( .A(n_1639), .B(n_1671), .Y(n_1670) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
NOR2x1_ASAP7_75t_R g1699 ( .A(n_1642), .B(n_1687), .Y(n_1699) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
NAND2xp5_ASAP7_75t_L g1667 ( .A(n_1644), .B(n_1668), .Y(n_1667) );
NAND2xp5_ASAP7_75t_L g1732 ( .A(n_1644), .B(n_1672), .Y(n_1732) );
INVxp67_ASAP7_75t_L g1645 ( .A(n_1646), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1648), .B(n_1650), .Y(n_1647) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
OAI22xp5_ASAP7_75t_SL g1651 ( .A1(n_1652), .A2(n_1654), .B1(n_1658), .B2(n_1659), .Y(n_1651) );
AOI21xp33_ASAP7_75t_L g1722 ( .A1(n_1652), .A2(n_1720), .B(n_1723), .Y(n_1722) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
AND2x2_ASAP7_75t_L g1763 ( .A(n_1653), .B(n_1764), .Y(n_1763) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1655), .B(n_1656), .Y(n_1654) );
AND2x2_ASAP7_75t_L g1757 ( .A(n_1655), .B(n_1713), .Y(n_1757) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
OR2x2_ASAP7_75t_L g1690 ( .A(n_1657), .B(n_1691), .Y(n_1690) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
AOI21xp33_ASAP7_75t_L g1695 ( .A1(n_1664), .A2(n_1696), .B(n_1698), .Y(n_1695) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1673), .Y(n_1745) );
NAND2xp5_ASAP7_75t_L g1748 ( .A(n_1673), .B(n_1749), .Y(n_1748) );
CKINVDCx5p33_ASAP7_75t_R g1768 ( .A(n_1673), .Y(n_1768) );
OR2x6_ASAP7_75t_SL g1673 ( .A(n_1674), .B(n_1678), .Y(n_1673) );
OAI22xp5_ASAP7_75t_L g1678 ( .A1(n_1679), .A2(n_1680), .B1(n_1681), .B2(n_1682), .Y(n_1678) );
NAND4xp25_ASAP7_75t_L g1683 ( .A(n_1684), .B(n_1700), .C(n_1708), .D(n_1715), .Y(n_1683) );
AOI211xp5_ASAP7_75t_SL g1684 ( .A1(n_1685), .A2(n_1686), .B(n_1689), .C(n_1695), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1687), .B(n_1688), .Y(n_1686) );
NAND2xp5_ASAP7_75t_L g1717 ( .A(n_1687), .B(n_1718), .Y(n_1717) );
NOR2x1_ASAP7_75t_L g1764 ( .A(n_1687), .B(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1688), .Y(n_1710) );
OAI31xp33_ASAP7_75t_L g1766 ( .A1(n_1688), .A2(n_1714), .A3(n_1767), .B(n_1769), .Y(n_1766) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1694), .Y(n_1762) );
INVxp67_ASAP7_75t_SL g1696 ( .A(n_1697), .Y(n_1696) );
INVxp33_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
NAND2xp33_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1706), .Y(n_1703) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1704), .Y(n_1714) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1705), .Y(n_1759) );
INVxp33_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
NAND2xp5_ASAP7_75t_L g1709 ( .A(n_1710), .B(n_1711), .Y(n_1709) );
NOR2xp33_ASAP7_75t_L g1758 ( .A(n_1712), .B(n_1759), .Y(n_1758) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
AOI22xp5_ASAP7_75t_L g1746 ( .A1(n_1719), .A2(n_1747), .B1(n_1750), .B2(n_1756), .Y(n_1746) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
NAND2xp5_ASAP7_75t_L g1723 ( .A(n_1724), .B(n_1726), .Y(n_1723) );
OAI21xp5_ASAP7_75t_SL g1750 ( .A1(n_1724), .A2(n_1751), .B(n_1752), .Y(n_1750) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
NAND5xp2_ASAP7_75t_L g1729 ( .A(n_1730), .B(n_1746), .C(n_1761), .D(n_1766), .E(n_1771), .Y(n_1729) );
OAI31xp33_ASAP7_75t_SL g1730 ( .A1(n_1731), .A2(n_1733), .A3(n_1738), .B(n_1744), .Y(n_1730) );
INVxp67_ASAP7_75t_SL g1731 ( .A(n_1732), .Y(n_1731) );
NOR2xp33_ASAP7_75t_L g1733 ( .A(n_1734), .B(n_1736), .Y(n_1733) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1735), .Y(n_1734) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1740), .Y(n_1742) );
CKINVDCx14_ASAP7_75t_R g1744 ( .A(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
INVx1_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
HB1xp67_ASAP7_75t_L g1772 ( .A(n_1773), .Y(n_1772) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
INVxp67_ASAP7_75t_SL g1775 ( .A(n_1776), .Y(n_1775) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
INVx1_ASAP7_75t_L g1777 ( .A(n_1778), .Y(n_1777) );
HB1xp67_ASAP7_75t_L g1830 ( .A(n_1779), .Y(n_1830) );
NAND2xp5_ASAP7_75t_SL g1791 ( .A(n_1792), .B(n_1800), .Y(n_1791) );
INVx1_ASAP7_75t_L g1804 ( .A(n_1805), .Y(n_1804) );
AOI31xp33_ASAP7_75t_SL g1807 ( .A1(n_1808), .A2(n_1811), .A3(n_1814), .B(n_1817), .Y(n_1807) );
CKINVDCx14_ASAP7_75t_R g1818 ( .A(n_1819), .Y(n_1818) );
BUFx2_ASAP7_75t_L g1819 ( .A(n_1820), .Y(n_1819) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1821), .Y(n_1820) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
INVx1_ASAP7_75t_L g1824 ( .A(n_1825), .Y(n_1824) );
CKINVDCx5p33_ASAP7_75t_R g1825 ( .A(n_1826), .Y(n_1825) );
A2O1A1Ixp33_ASAP7_75t_L g1834 ( .A1(n_1827), .A2(n_1835), .B(n_1837), .C(n_1838), .Y(n_1834) );
INVxp33_ASAP7_75t_SL g1828 ( .A(n_1829), .Y(n_1828) );
INVx1_ASAP7_75t_L g1832 ( .A(n_1830), .Y(n_1832) );
HB1xp67_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1836), .Y(n_1835) );
endmodule