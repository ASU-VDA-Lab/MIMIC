module fake_netlist_1_7236_n_717 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_717);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_717;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_47), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_77), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_7), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_71), .Y(n_83) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_76), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_72), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_20), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_35), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_56), .Y(n_88) );
INVxp33_ASAP7_75t_L g89 ( .A(n_79), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_41), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_69), .Y(n_92) );
HB1xp67_ASAP7_75t_L g93 ( .A(n_43), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_2), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_2), .Y(n_95) );
CKINVDCx11_ASAP7_75t_R g96 ( .A(n_58), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_63), .Y(n_97) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_40), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_74), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_26), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_66), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_7), .Y(n_102) );
BUFx2_ASAP7_75t_L g103 ( .A(n_57), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_1), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_39), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_55), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_73), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_16), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_21), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_53), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_5), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_24), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_30), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_48), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_13), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_25), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_37), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_54), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_62), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_38), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_17), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_36), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_34), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_27), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_67), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_65), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_10), .Y(n_127) );
CKINVDCx14_ASAP7_75t_R g128 ( .A(n_51), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_93), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_103), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_104), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_103), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_96), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g134 ( .A1(n_122), .A2(n_0), .B1(n_3), .B2(n_4), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_104), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_80), .B(n_4), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_84), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_82), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_89), .B(n_5), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_87), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_94), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_82), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_95), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_96), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_128), .B(n_6), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_122), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_95), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_102), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_126), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_84), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_111), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_126), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_84), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_90), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_81), .B(n_6), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_125), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_83), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_90), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_83), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g165 ( .A1(n_115), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_85), .B(n_8), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_101), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_101), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_124), .B(n_125), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_91), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_91), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_92), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_133), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_131), .B(n_117), .Y(n_174) );
INVx4_ASAP7_75t_L g175 ( .A(n_169), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_130), .B(n_129), .Y(n_177) );
NOR3xp33_ASAP7_75t_L g178 ( .A(n_165), .B(n_92), .C(n_123), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
BUFx4f_ASAP7_75t_L g180 ( .A(n_169), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_169), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
INVx5_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_151), .B(n_123), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_168), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
INVxp33_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_162), .B(n_109), .Y(n_188) );
INVxp67_ASAP7_75t_SL g189 ( .A(n_148), .Y(n_189) );
INVx1_ASAP7_75t_SL g190 ( .A(n_162), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_146), .B(n_117), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_141), .B(n_124), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_164), .B(n_108), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_164), .B(n_107), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_133), .B(n_9), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
INVx1_ASAP7_75t_SL g198 ( .A(n_167), .Y(n_198) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_141), .B(n_110), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_167), .B(n_106), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_159), .B(n_112), .Y(n_203) );
INVx4_ASAP7_75t_SL g204 ( .A(n_139), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_161), .B(n_105), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_147), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_152), .B(n_113), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_138), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_139), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_155), .B(n_121), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_149), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_170), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_149), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_170), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_149), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_171), .Y(n_218) );
OR2x2_ASAP7_75t_L g219 ( .A(n_147), .B(n_11), .Y(n_219) );
INVx1_ASAP7_75t_SL g220 ( .A(n_150), .Y(n_220) );
INVx2_ASAP7_75t_SL g221 ( .A(n_171), .Y(n_221) );
INVxp67_ASAP7_75t_SL g222 ( .A(n_172), .Y(n_222) );
NOR2x1p5_ASAP7_75t_L g223 ( .A(n_150), .B(n_99), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_157), .B(n_120), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_172), .B(n_119), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_137), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_137), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_140), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_154), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_142), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_142), .B(n_118), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_153), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_140), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_136), .A2(n_116), .B1(n_114), .B2(n_100), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_144), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_153), .B(n_97), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_193), .B(n_166), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_221), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_218), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_175), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_175), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_185), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_221), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_175), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_230), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_230), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_218), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_218), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_178), .A2(n_156), .B1(n_160), .B2(n_86), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_193), .B(n_156), .Y(n_250) );
NAND2x1p5_ASAP7_75t_L g251 ( .A(n_185), .B(n_132), .Y(n_251) );
NOR2xp33_ASAP7_75t_R g252 ( .A(n_173), .B(n_144), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_192), .B(n_134), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_199), .A2(n_88), .B1(n_98), .B2(n_154), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_189), .B(n_98), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_181), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_174), .B(n_98), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_226), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_180), .B(n_98), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_181), .B(n_98), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_226), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_211), .B(n_158), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_180), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_211), .B(n_158), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_226), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_173), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_181), .B(n_158), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_200), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_222), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_179), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_232), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_184), .B(n_158), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_180), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_184), .B(n_11), .Y(n_274) );
NOR2x1p5_ASAP7_75t_L g275 ( .A(n_206), .B(n_12), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_227), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_210), .Y(n_277) );
CKINVDCx11_ASAP7_75t_R g278 ( .A(n_220), .Y(n_278) );
NAND3xp33_ASAP7_75t_L g279 ( .A(n_177), .B(n_154), .C(n_139), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_199), .B(n_154), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_206), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_184), .B(n_12), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_227), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_192), .B(n_13), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_195), .B(n_45), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_214), .Y(n_286) );
OAI22xp33_ASAP7_75t_L g287 ( .A1(n_187), .A2(n_14), .B1(n_15), .B2(n_18), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_223), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_182), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_216), .Y(n_290) );
OR2x6_ASAP7_75t_L g291 ( .A(n_196), .B(n_14), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_197), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_176), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_224), .B(n_15), .Y(n_294) );
INVx4_ASAP7_75t_L g295 ( .A(n_224), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_190), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_176), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_188), .B(n_22), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_187), .B(n_23), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_231), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_236), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_203), .A2(n_28), .B(n_29), .Y(n_302) );
BUFx12f_ASAP7_75t_L g303 ( .A(n_233), .Y(n_303) );
INVx4_ASAP7_75t_L g304 ( .A(n_196), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_304), .B(n_198), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_295), .B(n_194), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_296), .Y(n_307) );
INVx2_ASAP7_75t_SL g308 ( .A(n_296), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_300), .B(n_202), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_237), .A2(n_205), .B(n_207), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_242), .Y(n_311) );
A2O1A1Ixp33_ASAP7_75t_L g312 ( .A1(n_292), .A2(n_225), .B(n_234), .C(n_219), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_301), .B(n_219), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_274), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_247), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_274), .A2(n_235), .B1(n_233), .B2(n_228), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_289), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_247), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_282), .A2(n_235), .B1(n_183), .B2(n_217), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_247), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_250), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_282), .A2(n_229), .B1(n_217), .B2(n_215), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_257), .A2(n_229), .B(n_215), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_247), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_280), .A2(n_213), .B(n_212), .C(n_208), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_267), .A2(n_213), .B(n_212), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_286), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_295), .B(n_204), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_255), .A2(n_208), .B(n_201), .Y(n_330) );
INVx5_ASAP7_75t_L g331 ( .A(n_273), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_304), .B(n_31), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_286), .Y(n_333) );
AOI22x1_ASAP7_75t_L g334 ( .A1(n_302), .A2(n_238), .B1(n_243), .B2(n_245), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_278), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_240), .Y(n_336) );
INVxp67_ASAP7_75t_L g337 ( .A(n_291), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_270), .B(n_204), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_241), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_278), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_280), .A2(n_201), .B(n_186), .C(n_204), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_245), .B(n_204), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_288), .B(n_32), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_286), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_273), .Y(n_345) );
CKINVDCx11_ASAP7_75t_R g346 ( .A(n_303), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_252), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_294), .A2(n_284), .B(n_287), .C(n_254), .Y(n_348) );
NOR2xp33_ASAP7_75t_SL g349 ( .A(n_291), .B(n_183), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_244), .Y(n_350) );
INVx4_ASAP7_75t_L g351 ( .A(n_273), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_286), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_253), .A2(n_186), .B1(n_183), .B2(n_191), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_266), .B(n_183), .C(n_209), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_252), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_281), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_291), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_313), .B(n_249), .Y(n_359) );
AO21x2_ASAP7_75t_L g360 ( .A1(n_348), .A2(n_298), .B(n_287), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_336), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_313), .B(n_249), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_337), .B(n_316), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_307), .B(n_251), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_309), .B(n_246), .Y(n_365) );
BUFx2_ASAP7_75t_R g366 ( .A(n_340), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_309), .B(n_251), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g368 ( .A(n_331), .B(n_273), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_310), .A2(n_298), .B(n_246), .Y(n_369) );
OAI21x1_ASAP7_75t_L g370 ( .A1(n_334), .A2(n_259), .B(n_299), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_333), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_341), .A2(n_259), .B(n_279), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_308), .A2(n_263), .B1(n_269), .B2(n_256), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_306), .B(n_268), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_333), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_326), .A2(n_272), .B(n_264), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_312), .B(n_268), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_333), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_306), .B(n_271), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_263), .B1(n_290), .B2(n_277), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_346), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_324), .A2(n_330), .B(n_327), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_339), .B(n_248), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_350), .B(n_248), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_344), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_328), .A2(n_262), .B(n_238), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_357), .A2(n_275), .B1(n_239), .B2(n_285), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_317), .A2(n_285), .B(n_243), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_344), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_305), .B(n_265), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_375), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_365), .B(n_332), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_365), .B(n_314), .Y(n_393) );
BUFx12f_ASAP7_75t_SL g394 ( .A(n_374), .Y(n_394) );
AOI222xp33_ASAP7_75t_L g395 ( .A1(n_363), .A2(n_335), .B1(n_355), .B2(n_349), .C1(n_319), .C2(n_347), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_358), .Y(n_396) );
BUFx10_ASAP7_75t_L g397 ( .A(n_381), .Y(n_397) );
AOI21xp33_ASAP7_75t_L g398 ( .A1(n_360), .A2(n_319), .B(n_332), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_358), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_367), .A2(n_335), .B1(n_321), .B2(n_356), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_361), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_367), .A2(n_323), .B1(n_311), .B2(n_344), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_361), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_364), .A2(n_331), .B1(n_351), .B2(n_345), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_359), .A2(n_353), .B1(n_331), .B2(n_276), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_383), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_370), .A2(n_352), .B(n_338), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
AOI22xp33_ASAP7_75t_SL g409 ( .A1(n_364), .A2(n_331), .B1(n_343), .B2(n_320), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_384), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_384), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_375), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_374), .B(n_320), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_362), .B(n_315), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_387), .A2(n_351), .B1(n_345), .B2(n_283), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_379), .B(n_318), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_377), .A2(n_260), .B1(n_258), .B2(n_329), .C(n_261), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_375), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_406), .B(n_360), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_406), .B(n_360), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_412), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_396), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_419), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_419), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_408), .B(n_390), .Y(n_427) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_408), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_410), .B(n_369), .Y(n_429) );
BUFx3_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_401), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_410), .B(n_386), .Y(n_432) );
INVx2_ASAP7_75t_R g433 ( .A(n_411), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_411), .B(n_386), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_392), .B(n_378), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_392), .A2(n_373), .B1(n_390), .B2(n_380), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_391), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_415), .Y(n_439) );
NOR2xp33_ASAP7_75t_R g440 ( .A(n_394), .B(n_366), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_399), .B(n_368), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_414), .B(n_369), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_417), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_412), .Y(n_444) );
OAI21x1_ASAP7_75t_L g445 ( .A1(n_413), .A2(n_370), .B(n_382), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_394), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_413), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_393), .B(n_368), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_391), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_391), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_414), .Y(n_451) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_398), .A2(n_382), .B(n_388), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_407), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_391), .B(n_389), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_391), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_428), .B(n_402), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_442), .B(n_407), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_422), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_442), .B(n_407), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_442), .B(n_400), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_453), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_422), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_446), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_424), .Y(n_464) );
OAI321xp33_ASAP7_75t_L g465 ( .A1(n_446), .A2(n_416), .A3(n_404), .B1(n_405), .B2(n_388), .C(n_418), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_428), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_430), .A2(n_395), .B1(n_409), .B2(n_260), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_424), .B(n_368), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_420), .B(n_389), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_438), .Y(n_470) );
INVx4_ASAP7_75t_L g471 ( .A(n_430), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_432), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_430), .A2(n_354), .B1(n_376), .B2(n_397), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_432), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_432), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_451), .A2(n_376), .B1(n_397), .B2(n_276), .Y(n_476) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_453), .A2(n_372), .B(n_389), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_420), .B(n_378), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_449), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_420), .B(n_378), .Y(n_480) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_445), .A2(n_452), .B(n_429), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_434), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_434), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_434), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_449), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_445), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_441), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_440), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_421), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_441), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_421), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_439), .B(n_371), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_443), .A2(n_397), .B1(n_325), .B2(n_385), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_439), .B(n_371), .Y(n_494) );
INVx4_ASAP7_75t_L g495 ( .A(n_438), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_431), .B(n_371), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_451), .B(n_385), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_449), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_431), .B(n_371), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_445), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_436), .B(n_375), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_436), .B(n_375), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_444), .B(n_372), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_444), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_447), .B(n_265), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_443), .B(n_265), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_460), .B(n_448), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_472), .B(n_452), .Y(n_508) );
INVx3_ASAP7_75t_L g509 ( .A(n_495), .Y(n_509) );
NOR2x1p5_ASAP7_75t_L g510 ( .A(n_463), .B(n_448), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_461), .Y(n_511) );
OAI31xp33_ASAP7_75t_SL g512 ( .A1(n_460), .A2(n_435), .A3(n_454), .B(n_447), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_487), .B(n_427), .Y(n_514) );
NAND4xp25_ASAP7_75t_L g515 ( .A(n_467), .B(n_437), .C(n_427), .D(n_429), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_458), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_490), .B(n_423), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_472), .B(n_452), .Y(n_518) );
NOR3xp33_ASAP7_75t_SL g519 ( .A(n_488), .B(n_465), .C(n_492), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_463), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_466), .B(n_423), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_462), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_474), .B(n_423), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_462), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_464), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_497), .B(n_435), .Y(n_526) );
NOR3xp33_ASAP7_75t_SL g527 ( .A(n_488), .B(n_329), .C(n_338), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_464), .Y(n_528) );
OAI221xp5_ASAP7_75t_L g529 ( .A1(n_493), .A2(n_426), .B1(n_425), .B2(n_455), .C(n_438), .Y(n_529) );
OAI211xp5_ASAP7_75t_L g530 ( .A1(n_493), .A2(n_454), .B(n_455), .C(n_438), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_504), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_463), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_474), .B(n_452), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_475), .B(n_433), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_475), .B(n_433), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_466), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_482), .B(n_425), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_461), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_482), .B(n_433), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_504), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_461), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_468), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_468), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_489), .B(n_435), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_489), .B(n_426), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_491), .B(n_426), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_483), .B(n_425), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_483), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_497), .B(n_435), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_484), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_484), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_496), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_499), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_491), .B(n_454), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_486), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_473), .B(n_450), .C(n_455), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_457), .B(n_450), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_499), .B(n_450), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_456), .B(n_455), .Y(n_559) );
NOR2xp67_ASAP7_75t_L g560 ( .A(n_471), .B(n_449), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_457), .B(n_449), .Y(n_561) );
OAI31xp33_ASAP7_75t_L g562 ( .A1(n_456), .A2(n_342), .A3(n_42), .B(n_44), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_496), .Y(n_563) );
OAI211xp5_ASAP7_75t_L g564 ( .A1(n_471), .A2(n_449), .B(n_265), .C(n_261), .Y(n_564) );
AOI31xp33_ASAP7_75t_L g565 ( .A1(n_476), .A2(n_342), .A3(n_46), .B(n_49), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_511), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_511), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_507), .B(n_459), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_543), .B(n_459), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_548), .B(n_469), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_541), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_550), .B(n_469), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_513), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_554), .B(n_478), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_516), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_522), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g577 ( .A1(n_515), .A2(n_494), .B1(n_492), .B2(n_465), .C(n_501), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_557), .B(n_480), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_524), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_557), .B(n_480), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_551), .B(n_514), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_552), .B(n_478), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_563), .B(n_503), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_526), .B(n_471), .Y(n_584) );
OR2x6_ASAP7_75t_L g585 ( .A(n_510), .B(n_471), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_553), .B(n_494), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_525), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_541), .Y(n_588) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_538), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_536), .B(n_502), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_528), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_542), .B(n_503), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_519), .A2(n_506), .B1(n_495), .B2(n_470), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_561), .B(n_481), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_531), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_544), .B(n_501), .Y(n_596) );
BUFx3_ASAP7_75t_L g597 ( .A(n_509), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_544), .B(n_502), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_561), .B(n_481), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_540), .B(n_506), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_519), .A2(n_470), .B1(n_495), .B2(n_505), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_517), .B(n_470), .Y(n_602) );
AND2x4_ASAP7_75t_L g603 ( .A(n_509), .B(n_495), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_508), .B(n_481), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_508), .B(n_481), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_549), .B(n_485), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_521), .B(n_477), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_518), .B(n_477), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_545), .B(n_477), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_547), .B(n_477), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_547), .B(n_505), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_518), .B(n_500), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_538), .Y(n_613) );
NOR2xp33_ASAP7_75t_SL g614 ( .A(n_520), .B(n_479), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_546), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_559), .B(n_498), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_533), .B(n_500), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_512), .B(n_500), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_573), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_575), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_581), .A2(n_533), .B1(n_529), .B2(n_530), .C(n_534), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_597), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_585), .B(n_509), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_618), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_597), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_568), .B(n_558), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_578), .B(n_532), .Y(n_627) );
AOI21xp33_ASAP7_75t_SL g628 ( .A1(n_585), .A2(n_565), .B(n_532), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_578), .B(n_534), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_576), .Y(n_630) );
INVxp67_ASAP7_75t_L g631 ( .A(n_602), .Y(n_631) );
OAI32xp33_ASAP7_75t_L g632 ( .A1(n_593), .A2(n_556), .A3(n_523), .B1(n_537), .B2(n_535), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_589), .Y(n_633) );
INVx2_ASAP7_75t_SL g634 ( .A(n_584), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_585), .A2(n_564), .B(n_560), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_604), .B(n_539), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_569), .B(n_539), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_577), .A2(n_562), .B1(n_535), .B2(n_479), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_579), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_587), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_589), .Y(n_641) );
AOI32xp33_ASAP7_75t_L g642 ( .A1(n_603), .A2(n_527), .A3(n_498), .B1(n_485), .B2(n_479), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_604), .B(n_555), .Y(n_643) );
AOI32xp33_ASAP7_75t_L g644 ( .A1(n_603), .A2(n_527), .A3(n_498), .B1(n_485), .B2(n_479), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_591), .A2(n_555), .B(n_486), .C(n_498), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_580), .B(n_486), .Y(n_646) );
NOR2xp33_ASAP7_75t_SL g647 ( .A(n_603), .B(n_485), .Y(n_647) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_601), .B(n_449), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_595), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_615), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_605), .B(n_33), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_566), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_586), .A2(n_261), .B1(n_276), .B2(n_209), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_580), .B(n_50), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g655 ( .A1(n_586), .A2(n_261), .B(n_276), .C(n_209), .Y(n_655) );
INVx2_ASAP7_75t_SL g656 ( .A(n_606), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_628), .A2(n_614), .B1(n_596), .B2(n_598), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_619), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_629), .B(n_599), .Y(n_659) );
AOI22x1_ASAP7_75t_L g660 ( .A1(n_635), .A2(n_609), .B1(n_607), .B2(n_613), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_624), .B(n_590), .Y(n_661) );
A2O1A1Ixp33_ASAP7_75t_SL g662 ( .A1(n_651), .A2(n_605), .B(n_608), .C(n_610), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_620), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_633), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_630), .Y(n_665) );
NAND4xp25_ASAP7_75t_L g666 ( .A(n_638), .B(n_608), .C(n_592), .D(n_582), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_639), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_640), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_649), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_650), .Y(n_670) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_632), .A2(n_599), .B(n_594), .C(n_583), .Y(n_671) );
AOI21xp33_ASAP7_75t_L g672 ( .A1(n_642), .A2(n_600), .B(n_616), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_621), .B(n_594), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_646), .Y(n_674) );
INVx3_ASAP7_75t_SL g675 ( .A(n_623), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_643), .B(n_617), .Y(n_676) );
NAND2xp33_ASAP7_75t_L g677 ( .A(n_644), .B(n_574), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_631), .A2(n_617), .B1(n_612), .B2(n_572), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_641), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g680 ( .A1(n_671), .A2(n_622), .B1(n_625), .B2(n_648), .C(n_655), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g681 ( .A1(n_677), .A2(n_623), .B(n_634), .C(n_655), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_657), .A2(n_625), .B(n_622), .C(n_654), .Y(n_682) );
OAI21xp5_ASAP7_75t_SL g683 ( .A1(n_657), .A2(n_648), .B(n_653), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_666), .A2(n_647), .B(n_645), .C(n_627), .Y(n_684) );
INVx1_ASAP7_75t_SL g685 ( .A(n_675), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_673), .A2(n_643), .B1(n_636), .B2(n_656), .C(n_626), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_660), .A2(n_647), .B(n_637), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_661), .A2(n_612), .B1(n_570), .B2(n_611), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_675), .B(n_652), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g690 ( .A(n_661), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_658), .Y(n_691) );
AOI321xp33_ASAP7_75t_L g692 ( .A1(n_672), .A2(n_588), .A3(n_571), .B1(n_567), .B2(n_566), .C(n_64), .Y(n_692) );
OAI21xp5_ASAP7_75t_L g693 ( .A1(n_662), .A2(n_588), .B(n_571), .Y(n_693) );
OAI21xp5_ASAP7_75t_L g694 ( .A1(n_682), .A2(n_662), .B(n_678), .Y(n_694) );
O2A1O1Ixp33_ASAP7_75t_L g695 ( .A1(n_684), .A2(n_670), .B(n_663), .C(n_665), .Y(n_695) );
OAI222xp33_ASAP7_75t_L g696 ( .A1(n_685), .A2(n_674), .B1(n_676), .B2(n_667), .C1(n_669), .C2(n_668), .Y(n_696) );
OAI211xp5_ASAP7_75t_L g697 ( .A1(n_683), .A2(n_681), .B(n_684), .C(n_680), .Y(n_697) );
OAI221xp5_ASAP7_75t_SL g698 ( .A1(n_686), .A2(n_659), .B1(n_664), .B2(n_679), .C(n_567), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_690), .A2(n_209), .B1(n_191), .B2(n_183), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_689), .A2(n_209), .B1(n_191), .B2(n_297), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_687), .B(n_297), .C(n_293), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_697), .Y(n_702) );
NOR3xp33_ASAP7_75t_SL g703 ( .A(n_694), .B(n_693), .C(n_692), .Y(n_703) );
NOR2x1_ASAP7_75t_L g704 ( .A(n_696), .B(n_691), .Y(n_704) );
XNOR2x1_ASAP7_75t_L g705 ( .A(n_700), .B(n_688), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_698), .B(n_52), .Y(n_706) );
XOR2xp5_ASAP7_75t_L g707 ( .A(n_702), .B(n_699), .Y(n_707) );
NOR3xp33_ASAP7_75t_L g708 ( .A(n_706), .B(n_695), .C(n_701), .Y(n_708) );
AOI31xp33_ASAP7_75t_L g709 ( .A1(n_704), .A2(n_59), .A3(n_60), .B(n_61), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_707), .Y(n_710) );
INVxp33_ASAP7_75t_SL g711 ( .A(n_708), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_710), .Y(n_712) );
OAI211xp5_ASAP7_75t_L g713 ( .A1(n_710), .A2(n_703), .B(n_709), .C(n_705), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_712), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_711), .B(n_713), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_710), .B1(n_191), .B2(n_293), .Y(n_716) );
OAI222xp33_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_68), .B1(n_70), .B2(n_75), .C1(n_78), .C2(n_191), .Y(n_717) );
endmodule