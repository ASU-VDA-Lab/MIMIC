module real_aes_8906_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g269 ( .A1(n_0), .A2(n_270), .B(n_271), .C(n_274), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_1), .B(n_211), .Y(n_275) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_3), .B(n_181), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_4), .A2(n_151), .B(n_154), .C(n_474), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_5), .A2(n_171), .B(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_6), .A2(n_171), .B(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_7), .B(n_211), .Y(n_520) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_8), .A2(n_138), .B(n_191), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_9), .A2(n_454), .B1(n_457), .B2(n_458), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_9), .Y(n_458) );
AND2x6_ASAP7_75t_L g151 ( .A(n_10), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_11), .A2(n_151), .B(n_154), .C(n_157), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_12), .A2(n_48), .B1(n_455), .B2(n_456), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_12), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_13), .B(n_43), .Y(n_115) );
INVx1_ASAP7_75t_L g490 ( .A(n_14), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_15), .B(n_161), .Y(n_476) );
INVx1_ASAP7_75t_L g143 ( .A(n_16), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_17), .B(n_181), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_18), .A2(n_159), .B(n_498), .C(n_500), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_19), .B(n_211), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_20), .B(n_235), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_21), .A2(n_154), .B(n_198), .C(n_231), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_22), .A2(n_163), .B(n_273), .C(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_23), .B(n_161), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_24), .B(n_161), .Y(n_541) );
CKINVDCx16_ASAP7_75t_R g548 ( .A(n_25), .Y(n_548) );
INVx1_ASAP7_75t_L g540 ( .A(n_26), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_27), .A2(n_154), .B(n_194), .C(n_198), .Y(n_193) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_28), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_29), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_30), .A2(n_104), .B1(n_116), .B2(n_742), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_31), .B(n_449), .Y(n_450) );
INVx1_ASAP7_75t_L g531 ( .A(n_32), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_33), .A2(n_171), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g149 ( .A(n_34), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_35), .A2(n_173), .B(n_184), .C(n_219), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_36), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_37), .A2(n_273), .B(n_517), .C(n_519), .Y(n_516) );
INVxp67_ASAP7_75t_L g532 ( .A(n_38), .Y(n_532) );
OAI321xp33_ASAP7_75t_L g122 ( .A1(n_39), .A2(n_123), .A3(n_445), .B1(n_446), .B2(n_447), .C(n_450), .Y(n_122) );
INVx1_ASAP7_75t_L g446 ( .A(n_39), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_40), .B(n_196), .Y(n_195) );
CKINVDCx14_ASAP7_75t_R g515 ( .A(n_41), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_42), .A2(n_154), .B(n_198), .C(n_539), .Y(n_538) );
AOI222xp33_ASAP7_75t_SL g452 ( .A1(n_44), .A2(n_453), .B1(n_459), .B2(n_733), .C1(n_734), .C2(n_738), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_45), .A2(n_274), .B(n_488), .C(n_489), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_46), .B(n_229), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_47), .Y(n_166) );
INVx1_ASAP7_75t_L g456 ( .A(n_48), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_49), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_50), .B(n_171), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_51), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_52), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_53), .A2(n_173), .B(n_175), .C(n_184), .Y(n_172) );
INVx1_ASAP7_75t_L g272 ( .A(n_54), .Y(n_272) );
INVx1_ASAP7_75t_L g176 ( .A(n_55), .Y(n_176) );
INVx1_ASAP7_75t_L g505 ( .A(n_56), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_57), .B(n_171), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_58), .A2(n_61), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_58), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_59), .Y(n_238) );
CKINVDCx14_ASAP7_75t_R g486 ( .A(n_60), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_61), .Y(n_126) );
INVx1_ASAP7_75t_L g152 ( .A(n_62), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_63), .B(n_171), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_64), .B(n_211), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_65), .A2(n_205), .B(n_207), .C(n_209), .Y(n_204) );
INVx1_ASAP7_75t_L g142 ( .A(n_66), .Y(n_142) );
INVx1_ASAP7_75t_SL g518 ( .A(n_67), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_68), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_69), .B(n_181), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_70), .B(n_211), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_71), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g551 ( .A(n_72), .Y(n_551) );
CKINVDCx16_ASAP7_75t_R g268 ( .A(n_73), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_74), .B(n_178), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_75), .A2(n_154), .B(n_184), .C(n_245), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g203 ( .A(n_76), .Y(n_203) );
INVx1_ASAP7_75t_L g109 ( .A(n_77), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_78), .A2(n_171), .B(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_79), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_80), .A2(n_171), .B(n_495), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_81), .A2(n_229), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g496 ( .A(n_82), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_83), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_84), .B(n_177), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_85), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_86), .A2(n_171), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g499 ( .A(n_87), .Y(n_499) );
INVx2_ASAP7_75t_L g140 ( .A(n_88), .Y(n_140) );
INVx1_ASAP7_75t_L g475 ( .A(n_89), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_90), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_91), .B(n_161), .Y(n_160) );
OR2x2_ASAP7_75t_L g111 ( .A(n_92), .B(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g462 ( .A(n_92), .B(n_113), .Y(n_462) );
INVx2_ASAP7_75t_L g732 ( .A(n_92), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_93), .A2(n_154), .B(n_184), .C(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_94), .B(n_171), .Y(n_217) );
INVx1_ASAP7_75t_L g220 ( .A(n_95), .Y(n_220) );
INVxp67_ASAP7_75t_L g208 ( .A(n_96), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_97), .B(n_138), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_98), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g145 ( .A(n_99), .Y(n_145) );
INVx1_ASAP7_75t_L g246 ( .A(n_100), .Y(n_246) );
INVx2_ASAP7_75t_L g508 ( .A(n_101), .Y(n_508) );
AND2x2_ASAP7_75t_L g187 ( .A(n_102), .B(n_186), .Y(n_187) );
BUFx4f_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
CKINVDCx6p67_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g743 ( .A(n_106), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_SL g445 ( .A(n_111), .Y(n_445) );
INVx1_ASAP7_75t_SL g449 ( .A(n_111), .Y(n_449) );
NOR2x2_ASAP7_75t_L g740 ( .A(n_112), .B(n_732), .Y(n_740) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g731 ( .A(n_113), .B(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_451), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g741 ( .A(n_121), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_123), .B(n_448), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_128), .B2(n_129), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22x1_ASAP7_75t_SL g734 ( .A1(n_128), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_734) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g459 ( .A1(n_129), .A2(n_460), .B1(n_463), .B2(n_729), .Y(n_459) );
OR3x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_343), .C(n_408), .Y(n_129) );
NAND4xp25_ASAP7_75t_SL g130 ( .A(n_131), .B(n_284), .C(n_310), .D(n_333), .Y(n_130) );
AOI221xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_212), .B1(n_253), .B2(n_260), .C(n_276), .Y(n_131) );
CKINVDCx14_ASAP7_75t_R g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_133), .A2(n_277), .B1(n_301), .B2(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_188), .Y(n_133) );
INVx1_ASAP7_75t_SL g337 ( .A(n_134), .Y(n_337) );
OR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_168), .Y(n_134) );
OR2x2_ASAP7_75t_L g258 ( .A(n_135), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g279 ( .A(n_135), .B(n_189), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_135), .B(n_199), .Y(n_292) );
AND2x2_ASAP7_75t_L g309 ( .A(n_135), .B(n_168), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_135), .B(n_256), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_135), .B(n_308), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_135), .B(n_188), .Y(n_430) );
AOI211xp5_ASAP7_75t_SL g441 ( .A1(n_135), .A2(n_347), .B(n_442), .C(n_443), .Y(n_441) );
INVx5_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_136), .B(n_189), .Y(n_313) );
AND2x2_ASAP7_75t_L g316 ( .A(n_136), .B(n_190), .Y(n_316) );
OR2x2_ASAP7_75t_L g361 ( .A(n_136), .B(n_189), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_136), .B(n_199), .Y(n_370) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_144), .B(n_165), .Y(n_136) );
INVx3_ASAP7_75t_L g211 ( .A(n_137), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_137), .B(n_223), .Y(n_222) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_137), .A2(n_243), .B(n_251), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_137), .B(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_137), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_137), .B(n_543), .Y(n_542) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_137), .A2(n_547), .B(n_553), .Y(n_546) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_138), .A2(n_192), .B(n_193), .Y(n_191) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_138), .Y(n_200) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g186 ( .A(n_140), .B(n_141), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_153), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_146), .A2(n_472), .B(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_146), .A2(n_186), .B(n_537), .C(n_538), .Y(n_536) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_146), .A2(n_548), .B(n_549), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
AND2x4_ASAP7_75t_L g171 ( .A(n_147), .B(n_151), .Y(n_171) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
INVx1_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
INVx1_ASAP7_75t_L g164 ( .A(n_149), .Y(n_164) );
INVx1_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx3_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
INVx1_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
INVx4_ASAP7_75t_SL g185 ( .A(n_151), .Y(n_185) );
BUFx3_ASAP7_75t_L g198 ( .A(n_151), .Y(n_198) );
INVx5_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx3_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_155), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_160), .B(n_162), .Y(n_157) );
INVx5_ASAP7_75t_L g181 ( .A(n_159), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_159), .B(n_490), .Y(n_489) );
INVx4_ASAP7_75t_L g273 ( .A(n_161), .Y(n_273) );
INVx2_ASAP7_75t_L g488 ( .A(n_161), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_162), .A2(n_195), .B(n_197), .Y(n_194) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVx2_ASAP7_75t_L g525 ( .A(n_167), .Y(n_525) );
INVx5_ASAP7_75t_SL g259 ( .A(n_168), .Y(n_259) );
AND2x2_ASAP7_75t_L g278 ( .A(n_168), .B(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_168), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g364 ( .A(n_168), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g396 ( .A(n_168), .B(n_199), .Y(n_396) );
OR2x2_ASAP7_75t_L g402 ( .A(n_168), .B(n_292), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_168), .B(n_352), .Y(n_411) );
OR2x6_ASAP7_75t_L g168 ( .A(n_169), .B(n_187), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_172), .B(n_186), .Y(n_169) );
BUFx2_ASAP7_75t_L g229 ( .A(n_171), .Y(n_229) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_174), .A2(n_185), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_SL g267 ( .A1(n_174), .A2(n_185), .B(n_268), .C(n_269), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_SL g485 ( .A1(n_174), .A2(n_185), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_174), .A2(n_185), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_174), .A2(n_185), .B(n_505), .C(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_174), .A2(n_185), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_SL g527 ( .A1(n_174), .A2(n_185), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_180), .C(n_182), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_177), .A2(n_182), .B(n_220), .C(n_221), .Y(n_219) );
O2A1O1Ixp5_ASAP7_75t_L g474 ( .A1(n_177), .A2(n_475), .B(n_476), .C(n_477), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_177), .A2(n_477), .B(n_551), .C(n_552), .Y(n_550) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx4_ASAP7_75t_L g206 ( .A(n_179), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_181), .B(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g270 ( .A(n_181), .Y(n_270) );
OAI22xp33_ASAP7_75t_L g530 ( .A1(n_181), .A2(n_206), .B1(n_531), .B2(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_181), .A2(n_234), .B(n_540), .C(n_541), .Y(n_539) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g274 ( .A(n_183), .Y(n_274) );
INVx1_ASAP7_75t_L g500 ( .A(n_183), .Y(n_500) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_186), .A2(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g236 ( .A(n_186), .Y(n_236) );
INVx1_ASAP7_75t_L g239 ( .A(n_186), .Y(n_239) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_186), .A2(n_484), .B(n_491), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_199), .Y(n_188) );
AND2x2_ASAP7_75t_L g293 ( .A(n_189), .B(n_259), .Y(n_293) );
INVx1_ASAP7_75t_SL g306 ( .A(n_189), .Y(n_306) );
OR2x2_ASAP7_75t_L g341 ( .A(n_189), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g347 ( .A(n_189), .B(n_199), .Y(n_347) );
AND2x2_ASAP7_75t_L g405 ( .A(n_189), .B(n_256), .Y(n_405) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_190), .B(n_259), .Y(n_332) );
INVx3_ASAP7_75t_L g256 ( .A(n_199), .Y(n_256) );
OR2x2_ASAP7_75t_L g298 ( .A(n_199), .B(n_259), .Y(n_298) );
AND2x2_ASAP7_75t_L g308 ( .A(n_199), .B(n_306), .Y(n_308) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_199), .Y(n_356) );
AND2x2_ASAP7_75t_L g365 ( .A(n_199), .B(n_279), .Y(n_365) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_210), .Y(n_199) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_200), .A2(n_494), .B(n_501), .Y(n_493) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_200), .A2(n_503), .B(n_509), .Y(n_502) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_200), .A2(n_513), .B(n_520), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_205), .A2(n_246), .B(n_247), .C(n_248), .Y(n_245) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_206), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_206), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g234 ( .A(n_209), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_209), .B(n_530), .Y(n_529) );
OA21x2_ASAP7_75t_L g265 ( .A1(n_211), .A2(n_266), .B(n_275), .Y(n_265) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_212), .A2(n_382), .B1(n_384), .B2(n_386), .C(n_389), .Y(n_381) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
AND2x2_ASAP7_75t_L g355 ( .A(n_214), .B(n_336), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_214), .B(n_414), .Y(n_418) );
OR2x2_ASAP7_75t_L g439 ( .A(n_214), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_214), .B(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx5_ASAP7_75t_L g286 ( .A(n_215), .Y(n_286) );
AND2x2_ASAP7_75t_L g363 ( .A(n_215), .B(n_226), .Y(n_363) );
AND2x2_ASAP7_75t_L g424 ( .A(n_215), .B(n_303), .Y(n_424) );
AND2x2_ASAP7_75t_L g437 ( .A(n_215), .B(n_256), .Y(n_437) );
OR2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_222), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_240), .Y(n_224) );
AND2x4_ASAP7_75t_L g263 ( .A(n_225), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g282 ( .A(n_225), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g289 ( .A(n_225), .Y(n_289) );
AND2x2_ASAP7_75t_L g358 ( .A(n_225), .B(n_336), .Y(n_358) );
AND2x2_ASAP7_75t_L g368 ( .A(n_225), .B(n_286), .Y(n_368) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_225), .Y(n_376) );
AND2x2_ASAP7_75t_L g388 ( .A(n_225), .B(n_265), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_225), .B(n_320), .Y(n_392) );
AND2x2_ASAP7_75t_L g429 ( .A(n_225), .B(n_424), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_225), .B(n_303), .Y(n_440) );
OR2x2_ASAP7_75t_L g442 ( .A(n_225), .B(n_378), .Y(n_442) );
INVx5_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g328 ( .A(n_226), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g338 ( .A(n_226), .B(n_283), .Y(n_338) );
AND2x2_ASAP7_75t_L g350 ( .A(n_226), .B(n_265), .Y(n_350) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_226), .Y(n_380) );
AND2x4_ASAP7_75t_L g414 ( .A(n_226), .B(n_264), .Y(n_414) );
OR2x6_ASAP7_75t_L g226 ( .A(n_227), .B(n_237), .Y(n_226) );
AOI21xp5_ASAP7_75t_SL g227 ( .A1(n_228), .A2(n_230), .B(n_235), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_236), .B(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AO21x2_ASAP7_75t_L g470 ( .A1(n_239), .A2(n_471), .B(n_478), .Y(n_470) );
BUFx2_ASAP7_75t_L g262 ( .A(n_240), .Y(n_262) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g303 ( .A(n_241), .Y(n_303) );
AND2x2_ASAP7_75t_L g336 ( .A(n_241), .B(n_265), .Y(n_336) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g283 ( .A(n_242), .B(n_265), .Y(n_283) );
BUFx2_ASAP7_75t_L g329 ( .A(n_242), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_250), .Y(n_243) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx3_ASAP7_75t_L g519 ( .A(n_249), .Y(n_519) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_255), .B(n_337), .Y(n_416) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_256), .B(n_279), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_256), .B(n_259), .Y(n_318) );
AND2x2_ASAP7_75t_L g373 ( .A(n_256), .B(n_309), .Y(n_373) );
AOI221xp5_ASAP7_75t_SL g310 ( .A1(n_257), .A2(n_311), .B1(n_319), .B2(n_321), .C(n_325), .Y(n_310) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g305 ( .A(n_258), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g346 ( .A(n_258), .B(n_347), .Y(n_346) );
OAI321xp33_ASAP7_75t_L g353 ( .A1(n_258), .A2(n_312), .A3(n_354), .B1(n_356), .B2(n_357), .C(n_359), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_259), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_262), .B(n_414), .Y(n_432) );
AND2x2_ASAP7_75t_L g319 ( .A(n_263), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_263), .B(n_323), .Y(n_322) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_264), .Y(n_295) );
AND2x2_ASAP7_75t_L g302 ( .A(n_264), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_264), .B(n_377), .Y(n_407) );
INVx1_ASAP7_75t_L g444 ( .A(n_264), .Y(n_444) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_273), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g477 ( .A(n_274), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B(n_281), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_278), .A2(n_388), .B(n_437), .C(n_438), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_279), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_279), .B(n_317), .Y(n_383) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g326 ( .A(n_283), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_283), .B(n_286), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_283), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_283), .B(n_368), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_287), .B1(n_299), .B2(n_304), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g300 ( .A(n_286), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g323 ( .A(n_286), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g335 ( .A(n_286), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_286), .B(n_329), .Y(n_371) );
OR2x2_ASAP7_75t_L g378 ( .A(n_286), .B(n_303), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_286), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g428 ( .A(n_286), .B(n_414), .Y(n_428) );
OAI22xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .B1(n_294), .B2(n_296), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g334 ( .A(n_289), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_292), .A2(n_307), .B1(n_375), .B2(n_379), .Y(n_374) );
INVx1_ASAP7_75t_L g422 ( .A(n_293), .Y(n_422) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g333 ( .A1(n_297), .A2(n_334), .B1(n_337), .B2(n_338), .C(n_339), .Y(n_333) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g312 ( .A(n_298), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_302), .B(n_368), .Y(n_400) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_303), .Y(n_320) );
INVx1_ASAP7_75t_L g324 ( .A(n_303), .Y(n_324) );
NAND2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g342 ( .A(n_309), .Y(n_342) );
AND2x2_ASAP7_75t_L g351 ( .A(n_309), .B(n_352), .Y(n_351) );
NAND2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx2_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g395 ( .A(n_316), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_319), .A2(n_345), .B1(n_348), .B2(n_351), .C(n_353), .Y(n_344) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_323), .B(n_380), .Y(n_379) );
AOI21xp33_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_327), .B(n_330), .Y(n_325) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
CKINVDCx16_ASAP7_75t_R g427 ( .A(n_330), .Y(n_427) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
OR2x2_ASAP7_75t_L g369 ( .A(n_332), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g390 ( .A(n_335), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_335), .B(n_395), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_338), .B(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND4xp25_ASAP7_75t_L g343 ( .A(n_344), .B(n_362), .C(n_381), .D(n_394), .Y(n_343) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g352 ( .A(n_347), .Y(n_352) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g385 ( .A(n_356), .B(n_361), .Y(n_385) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI211xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B(n_366), .C(n_374), .Y(n_362) );
AOI211xp5_ASAP7_75t_L g433 ( .A1(n_364), .A2(n_406), .B(n_434), .C(n_441), .Y(n_433) );
INVx1_ASAP7_75t_SL g393 ( .A(n_365), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B1(n_371), .B2(n_372), .Y(n_366) );
INVx1_ASAP7_75t_L g397 ( .A(n_371), .Y(n_397) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_377), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_377), .B(n_388), .Y(n_421) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g398 ( .A(n_388), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B(n_393), .Y(n_389) );
INVxp33_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI322xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .A3(n_398), .B1(n_399), .B2(n_401), .C1(n_403), .C2(n_406), .Y(n_394) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND3xp33_ASAP7_75t_SL g408 ( .A(n_409), .B(n_426), .C(n_433), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B1(n_415), .B2(n_417), .C(n_419), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g425 ( .A(n_414), .Y(n_425) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_429), .B2(n_430), .C(n_431), .Y(n_426) );
NAND2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVxp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_450), .B(n_452), .C(n_741), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_453), .Y(n_733) );
INVx1_ASAP7_75t_L g457 ( .A(n_454), .Y(n_457) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g735 ( .A(n_461), .Y(n_735) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g736 ( .A(n_463), .Y(n_736) );
OR2x2_ASAP7_75t_SL g463 ( .A(n_464), .B(n_684), .Y(n_463) );
NAND5xp2_ASAP7_75t_L g464 ( .A(n_465), .B(n_596), .C(n_634), .D(n_655), .E(n_672), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_568), .C(n_589), .Y(n_465) );
OAI221xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_510), .B1(n_534), .B2(n_555), .C(n_559), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_480), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_469), .B(n_557), .Y(n_576) );
OR2x2_ASAP7_75t_L g603 ( .A(n_469), .B(n_493), .Y(n_603) );
AND2x2_ASAP7_75t_L g617 ( .A(n_469), .B(n_493), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_469), .B(n_483), .Y(n_631) );
AND2x2_ASAP7_75t_L g669 ( .A(n_469), .B(n_633), .Y(n_669) );
AND2x2_ASAP7_75t_L g698 ( .A(n_469), .B(n_608), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_469), .B(n_580), .Y(n_715) );
INVx4_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g595 ( .A(n_470), .B(n_492), .Y(n_595) );
BUFx3_ASAP7_75t_L g620 ( .A(n_470), .Y(n_620) );
AND2x2_ASAP7_75t_L g649 ( .A(n_470), .B(n_493), .Y(n_649) );
AND3x2_ASAP7_75t_L g662 ( .A(n_470), .B(n_663), .C(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g585 ( .A(n_480), .Y(n_585) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_492), .Y(n_480) );
AOI32xp33_ASAP7_75t_L g640 ( .A1(n_481), .A2(n_592), .A3(n_641), .B1(n_644), .B2(n_645), .Y(n_640) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g567 ( .A(n_482), .B(n_492), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_482), .B(n_595), .Y(n_638) );
AND2x2_ASAP7_75t_L g645 ( .A(n_482), .B(n_617), .Y(n_645) );
OR2x2_ASAP7_75t_L g651 ( .A(n_482), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_482), .B(n_606), .Y(n_676) );
OR2x2_ASAP7_75t_L g694 ( .A(n_482), .B(n_522), .Y(n_694) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g558 ( .A(n_483), .B(n_502), .Y(n_558) );
INVx2_ASAP7_75t_L g580 ( .A(n_483), .Y(n_580) );
OR2x2_ASAP7_75t_L g602 ( .A(n_483), .B(n_502), .Y(n_602) );
AND2x2_ASAP7_75t_L g607 ( .A(n_483), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_483), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g663 ( .A(n_483), .B(n_557), .Y(n_663) );
INVx1_ASAP7_75t_SL g714 ( .A(n_492), .Y(n_714) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .Y(n_492) );
INVx1_ASAP7_75t_SL g557 ( .A(n_493), .Y(n_557) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_493), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_493), .B(n_643), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_493), .B(n_580), .C(n_698), .Y(n_709) );
INVx2_ASAP7_75t_L g608 ( .A(n_502), .Y(n_608) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_502), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_521), .Y(n_510) );
INVx1_ASAP7_75t_L g644 ( .A(n_511), .Y(n_644) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g562 ( .A(n_512), .B(n_545), .Y(n_562) );
INVx2_ASAP7_75t_L g579 ( .A(n_512), .Y(n_579) );
AND2x2_ASAP7_75t_L g584 ( .A(n_512), .B(n_546), .Y(n_584) );
AND2x2_ASAP7_75t_L g599 ( .A(n_512), .B(n_535), .Y(n_599) );
AND2x2_ASAP7_75t_L g611 ( .A(n_512), .B(n_583), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_521), .B(n_627), .Y(n_626) );
NAND2x1p5_ASAP7_75t_L g683 ( .A(n_521), .B(n_584), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_521), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_521), .B(n_578), .Y(n_706) );
BUFx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g544 ( .A(n_522), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_522), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g588 ( .A(n_522), .B(n_535), .Y(n_588) );
AND2x2_ASAP7_75t_L g614 ( .A(n_522), .B(n_545), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_522), .B(n_654), .Y(n_653) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_526), .B(n_533), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AO21x2_ASAP7_75t_L g572 ( .A1(n_524), .A2(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g573 ( .A(n_526), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_533), .Y(n_574) );
OR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_544), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_535), .B(n_565), .Y(n_564) );
AND2x4_ASAP7_75t_L g578 ( .A(n_535), .B(n_579), .Y(n_578) );
INVx3_ASAP7_75t_SL g583 ( .A(n_535), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_535), .B(n_570), .Y(n_636) );
OR2x2_ASAP7_75t_L g646 ( .A(n_535), .B(n_572), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_535), .B(n_614), .Y(n_674) );
OR2x2_ASAP7_75t_L g704 ( .A(n_535), .B(n_545), .Y(n_704) );
AND2x2_ASAP7_75t_L g708 ( .A(n_535), .B(n_546), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_535), .B(n_584), .Y(n_721) );
AND2x2_ASAP7_75t_L g728 ( .A(n_535), .B(n_610), .Y(n_728) );
OR2x6_ASAP7_75t_L g535 ( .A(n_536), .B(n_542), .Y(n_535) );
INVx1_ASAP7_75t_SL g671 ( .A(n_544), .Y(n_671) );
AND2x2_ASAP7_75t_L g610 ( .A(n_545), .B(n_572), .Y(n_610) );
AND2x2_ASAP7_75t_L g624 ( .A(n_545), .B(n_579), .Y(n_624) );
AND2x2_ASAP7_75t_L g627 ( .A(n_545), .B(n_583), .Y(n_627) );
INVx1_ASAP7_75t_L g654 ( .A(n_545), .Y(n_654) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
BUFx2_ASAP7_75t_L g566 ( .A(n_546), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g725 ( .A1(n_556), .A2(n_602), .B(n_726), .C(n_727), .Y(n_725) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g632 ( .A(n_557), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_558), .B(n_575), .Y(n_590) );
AND2x2_ASAP7_75t_L g616 ( .A(n_558), .B(n_617), .Y(n_616) );
OAI21xp5_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_563), .B(n_567), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_561), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g587 ( .A(n_562), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_562), .B(n_583), .Y(n_628) );
AND2x2_ASAP7_75t_L g719 ( .A(n_562), .B(n_570), .Y(n_719) );
INVxp67_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g592 ( .A(n_566), .B(n_579), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_566), .B(n_577), .Y(n_593) );
OAI322xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_576), .A3(n_577), .B1(n_580), .B2(n_581), .C1(n_585), .C2(n_586), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_575), .Y(n_569) );
AND2x2_ASAP7_75t_L g680 ( .A(n_570), .B(n_592), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_570), .B(n_644), .Y(n_726) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g623 ( .A(n_572), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g689 ( .A(n_576), .B(n_602), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_577), .B(n_671), .Y(n_670) );
INVx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_578), .B(n_610), .Y(n_667) );
AND2x2_ASAP7_75t_L g613 ( .A(n_579), .B(n_583), .Y(n_613) );
AND2x2_ASAP7_75t_L g621 ( .A(n_580), .B(n_622), .Y(n_621) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_580), .A2(n_659), .B(n_719), .C(n_720), .Y(n_718) );
AOI21xp33_ASAP7_75t_L g691 ( .A1(n_581), .A2(n_594), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_583), .B(n_610), .Y(n_650) );
AND2x2_ASAP7_75t_L g656 ( .A(n_583), .B(n_624), .Y(n_656) );
AND2x2_ASAP7_75t_L g690 ( .A(n_583), .B(n_592), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_584), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_SL g700 ( .A(n_584), .Y(n_700) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_588), .A2(n_616), .B1(n_618), .B2(n_623), .Y(n_615) );
OAI22xp5_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_591), .B1(n_593), .B2(n_594), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_590), .A2(n_626), .B1(n_628), .B2(n_629), .Y(n_625) );
INVxp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_595), .A2(n_697), .B1(n_699), .B2(n_701), .C(n_705), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_600), .B(n_604), .C(n_625), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
OR2x2_ASAP7_75t_L g666 ( .A(n_602), .B(n_619), .Y(n_666) );
INVx1_ASAP7_75t_L g717 ( .A(n_602), .Y(n_717) );
OAI221xp5_ASAP7_75t_L g604 ( .A1(n_603), .A2(n_605), .B1(n_609), .B2(n_612), .C(n_615), .Y(n_604) );
INVx2_ASAP7_75t_SL g659 ( .A(n_603), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g724 ( .A(n_606), .Y(n_724) );
AND2x2_ASAP7_75t_L g648 ( .A(n_607), .B(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g633 ( .A(n_608), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g695 ( .A(n_611), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_619), .B(n_721), .Y(n_720) );
CKINVDCx16_ASAP7_75t_R g619 ( .A(n_620), .Y(n_619) );
INVxp67_ASAP7_75t_L g664 ( .A(n_622), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_623), .A2(n_635), .B(n_637), .C(n_639), .Y(n_634) );
INVx1_ASAP7_75t_L g712 ( .A(n_626), .Y(n_712) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_630), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx2_ASAP7_75t_L g643 ( .A(n_633), .Y(n_643) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI222xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_646), .B1(n_647), .B2(n_650), .C1(n_651), .C2(n_653), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g679 ( .A(n_643), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_646), .B(n_700), .Y(n_699) );
NAND2xp33_ASAP7_75t_SL g677 ( .A(n_647), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g652 ( .A(n_649), .Y(n_652) );
AND2x2_ASAP7_75t_L g716 ( .A(n_649), .B(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g682 ( .A(n_652), .B(n_679), .Y(n_682) );
INVx1_ASAP7_75t_L g711 ( .A(n_653), .Y(n_711) );
AOI211xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B(n_660), .C(n_665), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_659), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AOI322xp5_ASAP7_75t_L g710 ( .A1(n_662), .A2(n_690), .A3(n_695), .B1(n_711), .B2(n_712), .C1(n_713), .C2(n_716), .Y(n_710) );
AND2x2_ASAP7_75t_L g697 ( .A(n_663), .B(n_698), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_668), .B2(n_670), .Y(n_665) );
INVxp33_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B1(n_677), .B2(n_680), .C(n_681), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NAND5xp2_ASAP7_75t_L g684 ( .A(n_685), .B(n_696), .C(n_710), .D(n_718), .E(n_722), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_690), .B(n_691), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVxp33_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g722 ( .A1(n_698), .A2(n_723), .B(n_724), .C(n_725), .Y(n_722) );
AOI31xp33_ASAP7_75t_L g705 ( .A1(n_700), .A2(n_706), .A3(n_707), .B(n_709), .Y(n_705) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g723 ( .A(n_721), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g737 ( .A(n_730), .Y(n_737) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
endmodule