module real_jpeg_29925_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_0),
.A2(n_26),
.B1(n_33),
.B2(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_0),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_1),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_88)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_2),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_3),
.A2(n_26),
.B1(n_33),
.B2(n_49),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_49),
.B1(n_62),
.B2(n_63),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_4),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_4),
.A2(n_61),
.B(n_62),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_100),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_4),
.B(n_39),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_39),
.B(n_43),
.C(n_181),
.D(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_4),
.B(n_71),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_4),
.A2(n_25),
.B(n_194),
.Y(n_212)
);

A2O1A1O1Ixp25_ASAP7_75t_L g224 ( 
.A1(n_4),
.A2(n_63),
.B(n_74),
.C(n_113),
.D(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_4),
.B(n_63),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_5),
.A2(n_26),
.B1(n_33),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_5),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_8),
.A2(n_56),
.B1(n_57),
.B2(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_8),
.A2(n_26),
.B1(n_33),
.B2(n_66),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_66),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_10),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_80),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_80),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_10),
.A2(n_26),
.B1(n_33),
.B2(n_80),
.Y(n_196)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_11),
.B(n_39),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_45),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_11),
.B(n_26),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_12),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_12),
.A2(n_39),
.B1(n_40),
.B2(n_55),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_55),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_13),
.A2(n_41),
.B1(n_62),
.B2(n_63),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_41),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_135),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_114),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_21),
.B(n_114),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.C(n_89),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_22),
.B(n_81),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_53),
.C(n_67),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_24),
.B(n_37),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_25),
.A2(n_35),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_25),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_25),
.A2(n_83),
.B(n_85),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_25),
.A2(n_83),
.B1(n_106),
.B2(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_25),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_25),
.B(n_196),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_31),
.A2(n_84),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

AOI32xp33_ASAP7_75t_L g180 ( 
.A1(n_33),
.A2(n_40),
.A3(n_45),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_33),
.B(n_214),
.Y(n_213)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_38),
.A2(n_50),
.B(n_147),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_44),
.B(n_46),
.C(n_47),
.Y(n_43)
);

AOI32xp33_ASAP7_75t_L g232 ( 
.A1(n_39),
.A2(n_62),
.A3(n_225),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_40),
.B(n_76),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_48),
.B1(n_50),
.B2(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_42),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_43),
.A2(n_47),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_43),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_43),
.A2(n_47),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_50),
.B(n_149),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_50),
.A2(n_147),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_50),
.B(n_100),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_67),
.B2(n_68),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B1(n_59),
.B2(n_65),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_56),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_60),
.B(n_100),
.C(n_101),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_58),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_59),
.B(n_96),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_63),
.B1(n_72),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_65),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B(n_73),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_69),
.A2(n_70),
.B1(n_109),
.B2(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_79),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_70),
.A2(n_73),
.B(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_71),
.A2(n_74),
.B1(n_111),
.B2(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_76),
.Y(n_233)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_87),
.Y(n_124)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_83),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_83),
.A2(n_201),
.B(n_209),
.Y(n_208)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_84),
.B(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_84),
.A2(n_210),
.B(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_88),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_89),
.A2(n_90),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.C(n_107),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_91),
.A2(n_92),
.B1(n_107),
.B2(n_108),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B(n_95),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_94),
.B(n_100),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_100),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_104),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B(n_112),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_134),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_123),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_133),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B(n_130),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_173),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_159),
.B(n_172),
.Y(n_138)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_139),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_156),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_140),
.B(n_156),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.C(n_144),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_144),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.C(n_153),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_146),
.B1(n_153),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_150),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_160),
.B(n_162),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.C(n_167),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_163),
.B(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_166),
.B(n_167),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.C(n_171),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_168),
.B(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_169),
.B(n_171),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_170),
.Y(n_231)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_252),
.C(n_253),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_247),
.B(n_251),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_236),
.B(n_246),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_220),
.B(n_235),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_197),
.B(n_219),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_179),
.B(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_183),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_193),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_205),
.B(n_218),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_199),
.B(n_204),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_211),
.B(n_217),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_207),
.B(n_208),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_221),
.B(n_222),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_226),
.C(n_229),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_232),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_238),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_249),
.Y(n_251)
);


endmodule