module real_aes_7630_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_503;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g233 ( .A(n_0), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_1), .A2(n_28), .B1(n_223), .B2(n_270), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_2), .B(n_242), .Y(n_250) );
INVx1_ASAP7_75t_L g196 ( .A(n_3), .Y(n_196) );
AND2x6_ASAP7_75t_L g238 ( .A(n_3), .B(n_194), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_3), .B(n_530), .Y(n_529) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_4), .A2(n_23), .B1(n_91), .B2(n_92), .Y(n_90) );
INVx1_ASAP7_75t_L g214 ( .A(n_5), .Y(n_214) );
INVx1_ASAP7_75t_L g217 ( .A(n_6), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_7), .A2(n_37), .B1(n_155), .B2(n_159), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_8), .B(n_219), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_9), .B(n_210), .Y(n_316) );
AO32x2_ASAP7_75t_L g286 ( .A1(n_10), .A2(n_209), .A3(n_242), .B1(n_261), .B2(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_11), .B(n_223), .Y(n_283) );
OAI22xp5_ASAP7_75t_SL g175 ( .A1(n_12), .A2(n_29), .B1(n_176), .B2(n_177), .Y(n_175) );
INVx1_ASAP7_75t_L g177 ( .A(n_12), .Y(n_177) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_13), .A2(n_26), .B1(n_91), .B2(n_95), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_14), .B(n_210), .Y(n_239) );
INVx1_ASAP7_75t_L g85 ( .A(n_15), .Y(n_85) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_16), .A2(n_172), .B1(n_179), .B2(n_180), .Y(n_171) );
INVx1_ASAP7_75t_L g179 ( .A(n_16), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_16), .A2(n_36), .B1(n_223), .B2(n_270), .Y(n_289) );
AOI22xp33_ASAP7_75t_SL g272 ( .A1(n_17), .A2(n_61), .B1(n_219), .B2(n_223), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_18), .B(n_223), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_18), .A2(n_81), .B1(n_169), .B2(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_18), .Y(n_528) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_19), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_20), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_21), .B(n_263), .Y(n_304) );
INVx2_ASAP7_75t_L g221 ( .A(n_22), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_24), .B(n_223), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_25), .B(n_263), .Y(n_285) );
OAI221xp5_ASAP7_75t_L g187 ( .A1(n_26), .A2(n_42), .B1(n_56), .B2(n_188), .C(n_189), .Y(n_187) );
INVxp67_ASAP7_75t_L g190 ( .A(n_26), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_27), .A2(n_81), .B1(n_168), .B2(n_169), .Y(n_80) );
INVx1_ASAP7_75t_L g168 ( .A(n_27), .Y(n_168) );
INVx1_ASAP7_75t_L g176 ( .A(n_29), .Y(n_176) );
AOI22xp33_ASAP7_75t_SL g136 ( .A1(n_30), .A2(n_74), .B1(n_137), .B2(n_141), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_31), .B(n_223), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_32), .A2(n_68), .B1(n_270), .B2(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_33), .B(n_223), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_34), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_35), .B(n_231), .Y(n_249) );
AOI22xp33_ASAP7_75t_SL g314 ( .A1(n_38), .A2(n_45), .B1(n_219), .B2(n_223), .Y(n_314) );
INVx1_ASAP7_75t_L g125 ( .A(n_39), .Y(n_125) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_40), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_40), .B(n_223), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_41), .B(n_223), .Y(n_278) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_42), .A2(n_64), .B1(n_91), .B2(n_95), .Y(n_100) );
INVxp67_ASAP7_75t_L g191 ( .A(n_42), .Y(n_191) );
INVx1_ASAP7_75t_L g131 ( .A(n_43), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_44), .A2(n_59), .B1(n_182), .B2(n_183), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_44), .Y(n_182) );
INVx1_ASAP7_75t_L g194 ( .A(n_46), .Y(n_194) );
AOI22xp33_ASAP7_75t_SL g162 ( .A1(n_47), .A2(n_75), .B1(n_163), .B2(n_165), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_48), .B(n_223), .Y(n_234) );
INVx1_ASAP7_75t_L g213 ( .A(n_49), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_50), .Y(n_188) );
AO32x2_ASAP7_75t_L g267 ( .A1(n_51), .A2(n_242), .A3(n_261), .B1(n_268), .B2(n_273), .Y(n_267) );
INVx1_ASAP7_75t_L g257 ( .A(n_52), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_53), .A2(n_60), .B1(n_147), .B2(n_149), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g114 ( .A1(n_54), .A2(n_58), .B1(n_115), .B2(n_120), .Y(n_114) );
INVx1_ASAP7_75t_L g299 ( .A(n_55), .Y(n_299) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_56), .A2(n_71), .B1(n_91), .B2(n_92), .Y(n_98) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_57), .B(n_219), .Y(n_300) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_59), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_62), .B(n_270), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_63), .B(n_219), .Y(n_303) );
INVx1_ASAP7_75t_L g536 ( .A(n_63), .Y(n_536) );
INVx1_ASAP7_75t_L g107 ( .A(n_65), .Y(n_107) );
INVx2_ASAP7_75t_L g211 ( .A(n_66), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_67), .B(n_219), .Y(n_246) );
INVx1_ASAP7_75t_L g101 ( .A(n_69), .Y(n_101) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_70), .A2(n_77), .B1(n_219), .B2(n_220), .Y(n_313) );
INVx1_ASAP7_75t_L g91 ( .A(n_72), .Y(n_91) );
INVx1_ASAP7_75t_L g93 ( .A(n_72), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_73), .B(n_219), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_76), .A2(n_81), .B1(n_169), .B2(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_76), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_184), .B1(n_197), .B2(n_518), .C(n_526), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_170), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_81), .Y(n_169) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
AND2x2_ASAP7_75t_L g82 ( .A(n_83), .B(n_134), .Y(n_82) );
NOR3xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_106), .C(n_124), .Y(n_83) );
OAI22xp5_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_86), .B1(n_101), .B2(n_102), .Y(n_84) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
OR2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_96), .Y(n_87) );
INVx2_ASAP7_75t_L g140 ( .A(n_88), .Y(n_140) );
OR2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
AND2x2_ASAP7_75t_L g105 ( .A(n_89), .B(n_94), .Y(n_105) );
AND2x2_ASAP7_75t_L g145 ( .A(n_89), .B(n_130), .Y(n_145) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g111 ( .A(n_90), .B(n_94), .Y(n_111) );
AND2x2_ASAP7_75t_L g119 ( .A(n_90), .B(n_100), .Y(n_119) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g95 ( .A(n_93), .Y(n_95) );
INVx2_ASAP7_75t_L g130 ( .A(n_94), .Y(n_130) );
INVx1_ASAP7_75t_L g167 ( .A(n_94), .Y(n_167) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
NAND2x1p5_ASAP7_75t_L g104 ( .A(n_97), .B(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g164 ( .A(n_97), .B(n_145), .Y(n_164) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_99), .Y(n_97) );
INVx1_ASAP7_75t_L g113 ( .A(n_98), .Y(n_113) );
INVx1_ASAP7_75t_L g118 ( .A(n_98), .Y(n_118) );
INVx1_ASAP7_75t_L g123 ( .A(n_98), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_98), .B(n_100), .Y(n_152) );
AND2x2_ASAP7_75t_L g112 ( .A(n_99), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g144 ( .A(n_100), .B(n_123), .Y(n_144) );
BUFx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx3_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g158 ( .A(n_105), .B(n_112), .Y(n_158) );
AND2x2_ASAP7_75t_L g161 ( .A(n_105), .B(n_144), .Y(n_161) );
OAI21xp33_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_108), .B(n_114), .Y(n_106) );
INVx2_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x6_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x4_ASAP7_75t_L g121 ( .A(n_111), .B(n_122), .Y(n_121) );
AND2x6_ASAP7_75t_L g139 ( .A(n_112), .B(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g148 ( .A(n_112), .B(n_145), .Y(n_148) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g129 ( .A(n_118), .B(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g128 ( .A(n_119), .B(n_129), .Y(n_128) );
NAND2x1p5_ASAP7_75t_L g132 ( .A(n_119), .B(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_131), .B2(n_132), .Y(n_124) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g133 ( .A(n_130), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_153), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_146), .Y(n_135) );
INVx5_ASAP7_75t_SL g137 ( .A(n_138), .Y(n_137) );
INVx11_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx4f_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x4_ASAP7_75t_L g150 ( .A(n_145), .B(n_151), .Y(n_150) );
BUFx2_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
BUFx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OR2x6_ASAP7_75t_L g166 ( .A(n_152), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_162), .Y(n_153) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx8_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
XNOR2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_181), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_172), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B1(n_175), .B2(n_178), .Y(n_172) );
INVx1_ASAP7_75t_L g178 ( .A(n_173), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
AND3x1_ASAP7_75t_SL g186 ( .A(n_187), .B(n_192), .C(n_195), .Y(n_186) );
INVxp67_ASAP7_75t_L g530 ( .A(n_187), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_192), .A2(n_533), .B(n_535), .Y(n_532) );
INVx1_ASAP7_75t_L g540 ( .A(n_192), .Y(n_540) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OAI322xp33_ASAP7_75t_L g526 ( .A1(n_193), .A2(n_527), .A3(n_529), .B1(n_531), .B2(n_536), .C1(n_537), .C2(n_539), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_193), .B(n_196), .Y(n_535) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OR2x2_ASAP7_75t_SL g539 ( .A(n_195), .B(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_199), .B(n_484), .Y(n_198) );
NOR3xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_388), .C(n_472), .Y(n_199) );
NAND4xp25_ASAP7_75t_L g200 ( .A(n_201), .B(n_331), .C(n_353), .D(n_369), .Y(n_200) );
AOI221xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_264), .B1(n_290), .B2(n_309), .C(n_317), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_240), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_204), .B(n_309), .Y(n_343) );
NAND4xp25_ASAP7_75t_L g383 ( .A(n_204), .B(n_371), .C(n_384), .D(n_386), .Y(n_383) );
INVxp67_ASAP7_75t_L g500 ( .A(n_204), .Y(n_500) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_L g382 ( .A(n_205), .B(n_320), .Y(n_382) );
AND2x2_ASAP7_75t_L g406 ( .A(n_205), .B(n_240), .Y(n_406) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g373 ( .A(n_206), .B(n_308), .Y(n_373) );
AND2x2_ASAP7_75t_L g413 ( .A(n_206), .B(n_394), .Y(n_413) );
AND2x2_ASAP7_75t_L g430 ( .A(n_206), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_206), .B(n_241), .Y(n_454) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g307 ( .A(n_207), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g325 ( .A(n_207), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g337 ( .A(n_207), .B(n_241), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_207), .B(n_251), .Y(n_359) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_215), .B(n_239), .Y(n_207) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_208), .A2(n_252), .B(n_262), .Y(n_251) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_210), .Y(n_242) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
AND2x2_ASAP7_75t_SL g263 ( .A(n_211), .B(n_212), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_229), .B(n_238), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_222), .C(n_225), .Y(n_216) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g224 ( .A(n_221), .Y(n_224) );
INVx1_ASAP7_75t_L g232 ( .A(n_221), .Y(n_232) );
INVx3_ASAP7_75t_L g298 ( .A(n_223), .Y(n_298) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g270 ( .A(n_224), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_224), .Y(n_271) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_226), .A2(n_302), .B(n_303), .Y(n_301) );
INVx4_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g523 ( .A(n_227), .Y(n_523) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g237 ( .A(n_228), .Y(n_237) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_228), .Y(n_260) );
INVx1_ASAP7_75t_L g281 ( .A(n_228), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_233), .B(n_234), .C(n_235), .Y(n_229) );
O2A1O1Ixp5_ASAP7_75t_L g256 ( .A1(n_230), .A2(n_257), .B(n_258), .C(n_259), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_230), .B(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_230), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_235), .A2(n_248), .B(n_249), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_235), .A2(n_260), .B1(n_288), .B2(n_289), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_235), .A2(n_260), .B1(n_313), .B2(n_314), .Y(n_312) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_236), .A2(n_245), .B(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_236), .A2(n_254), .B(n_255), .Y(n_253) );
O2A1O1Ixp5_ASAP7_75t_SL g297 ( .A1(n_236), .A2(n_298), .B(n_299), .C(n_300), .Y(n_297) );
INVx5_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OAI22xp5_ASAP7_75t_SL g268 ( .A1(n_237), .A2(n_260), .B1(n_269), .B2(n_272), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_238), .A2(n_244), .B(n_247), .Y(n_243) );
BUFx3_ASAP7_75t_L g261 ( .A(n_238), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g276 ( .A1(n_238), .A2(n_277), .B(n_282), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_238), .A2(n_297), .B(n_301), .Y(n_296) );
INVx4_ASAP7_75t_SL g525 ( .A(n_238), .Y(n_525) );
AND2x2_ASAP7_75t_L g340 ( .A(n_240), .B(n_341), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_240), .A2(n_390), .B1(n_393), .B2(n_395), .C(n_399), .Y(n_389) );
AND2x2_ASAP7_75t_L g448 ( .A(n_240), .B(n_413), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_240), .B(n_430), .Y(n_482) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_251), .Y(n_240) );
INVx3_ASAP7_75t_L g308 ( .A(n_241), .Y(n_308) );
AND2x2_ASAP7_75t_L g357 ( .A(n_241), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g411 ( .A(n_241), .B(n_326), .Y(n_411) );
AND2x2_ASAP7_75t_L g469 ( .A(n_241), .B(n_470), .Y(n_469) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_250), .Y(n_241) );
INVx4_ASAP7_75t_L g311 ( .A(n_242), .Y(n_311) );
AND2x2_ASAP7_75t_L g309 ( .A(n_251), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g326 ( .A(n_251), .Y(n_326) );
INVx1_ASAP7_75t_L g381 ( .A(n_251), .Y(n_381) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_251), .Y(n_387) );
AND2x2_ASAP7_75t_L g432 ( .A(n_251), .B(n_308), .Y(n_432) );
OR2x2_ASAP7_75t_L g471 ( .A(n_251), .B(n_310), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_256), .B(n_261), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_259), .A2(n_283), .B(n_284), .Y(n_282) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND3xp33_ASAP7_75t_L g330 ( .A(n_261), .B(n_311), .C(n_312), .Y(n_330) );
INVx2_ASAP7_75t_L g273 ( .A(n_263), .Y(n_273) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_263), .A2(n_276), .B(n_285), .Y(n_275) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_263), .A2(n_296), .B(n_304), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_264), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_274), .Y(n_264) );
AND2x2_ASAP7_75t_L g467 ( .A(n_265), .B(n_464), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_265), .B(n_449), .Y(n_499) );
BUFx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g398 ( .A(n_266), .B(n_322), .Y(n_398) );
AND2x2_ASAP7_75t_L g447 ( .A(n_266), .B(n_293), .Y(n_447) );
INVx1_ASAP7_75t_L g493 ( .A(n_266), .Y(n_493) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_267), .Y(n_306) );
AND2x2_ASAP7_75t_L g348 ( .A(n_267), .B(n_322), .Y(n_348) );
INVx1_ASAP7_75t_L g365 ( .A(n_267), .Y(n_365) );
AND2x2_ASAP7_75t_L g371 ( .A(n_267), .B(n_286), .Y(n_371) );
AND2x2_ASAP7_75t_L g439 ( .A(n_274), .B(n_347), .Y(n_439) );
INVx2_ASAP7_75t_L g504 ( .A(n_274), .Y(n_504) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_286), .Y(n_274) );
AND2x2_ASAP7_75t_L g321 ( .A(n_275), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g334 ( .A(n_275), .B(n_294), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_275), .B(n_293), .Y(n_362) );
INVx1_ASAP7_75t_L g368 ( .A(n_275), .Y(n_368) );
INVx1_ASAP7_75t_L g385 ( .A(n_275), .Y(n_385) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_275), .Y(n_397) );
INVx2_ASAP7_75t_L g465 ( .A(n_275), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_279), .B(n_280), .Y(n_277) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g322 ( .A(n_286), .Y(n_322) );
BUFx2_ASAP7_75t_L g419 ( .A(n_286), .Y(n_419) );
AND2x2_ASAP7_75t_L g464 ( .A(n_286), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_305), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_292), .B(n_401), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_292), .A2(n_463), .B(n_477), .Y(n_487) );
AND2x2_ASAP7_75t_L g512 ( .A(n_292), .B(n_398), .Y(n_512) );
BUFx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g434 ( .A(n_294), .Y(n_434) );
AND2x2_ASAP7_75t_L g463 ( .A(n_294), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_295), .Y(n_347) );
INVx2_ASAP7_75t_L g366 ( .A(n_295), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_295), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx2_ASAP7_75t_L g320 ( .A(n_306), .Y(n_320) );
OR2x2_ASAP7_75t_L g333 ( .A(n_306), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g401 ( .A(n_306), .B(n_397), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_306), .B(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g502 ( .A(n_306), .B(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_306), .B(n_439), .Y(n_514) );
AND2x2_ASAP7_75t_L g393 ( .A(n_307), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g416 ( .A(n_307), .B(n_309), .Y(n_416) );
INVx2_ASAP7_75t_L g328 ( .A(n_308), .Y(n_328) );
AND2x2_ASAP7_75t_L g356 ( .A(n_308), .B(n_329), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_308), .B(n_381), .Y(n_437) );
AND2x2_ASAP7_75t_L g351 ( .A(n_309), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g498 ( .A(n_309), .Y(n_498) );
AND2x2_ASAP7_75t_L g510 ( .A(n_309), .B(n_373), .Y(n_510) );
AND2x2_ASAP7_75t_L g336 ( .A(n_310), .B(n_326), .Y(n_336) );
INVx1_ASAP7_75t_L g431 ( .A(n_310), .Y(n_431) );
AO21x1_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B(n_315), .Y(n_310) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g329 ( .A(n_316), .B(n_330), .Y(n_329) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_323), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_320), .B(n_367), .Y(n_376) );
OR2x2_ASAP7_75t_L g508 ( .A(n_320), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g425 ( .A(n_321), .B(n_366), .Y(n_425) );
AND2x2_ASAP7_75t_L g433 ( .A(n_321), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g492 ( .A(n_321), .B(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g516 ( .A(n_321), .B(n_363), .Y(n_516) );
NOR2xp67_ASAP7_75t_L g474 ( .A(n_322), .B(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g503 ( .A(n_322), .B(n_366), .Y(n_503) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2x1p5_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
AND2x2_ASAP7_75t_L g355 ( .A(n_325), .B(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g517 ( .A(n_325), .Y(n_517) );
NOR2x1_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g352 ( .A(n_328), .Y(n_352) );
AND2x2_ASAP7_75t_L g403 ( .A(n_328), .B(n_336), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_328), .B(n_471), .Y(n_497) );
INVx2_ASAP7_75t_L g342 ( .A(n_329), .Y(n_342) );
INVx3_ASAP7_75t_L g394 ( .A(n_329), .Y(n_394) );
OR2x2_ASAP7_75t_L g422 ( .A(n_329), .B(n_423), .Y(n_422) );
AOI311xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .A3(n_337), .B(n_338), .C(n_349), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g369 ( .A1(n_332), .A2(n_370), .B(n_372), .C(n_374), .Y(n_369) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_SL g354 ( .A(n_334), .Y(n_354) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g372 ( .A(n_336), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_336), .B(n_352), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_336), .B(n_337), .Y(n_505) );
AND2x2_ASAP7_75t_L g427 ( .A(n_337), .B(n_341), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_343), .B(n_344), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g485 ( .A(n_341), .B(n_373), .Y(n_485) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_342), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g379 ( .A(n_342), .Y(n_379) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
AND2x2_ASAP7_75t_L g370 ( .A(n_346), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g415 ( .A(n_348), .Y(n_415) );
AND2x4_ASAP7_75t_L g477 ( .A(n_348), .B(n_446), .Y(n_477) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI222xp33_ASAP7_75t_L g428 ( .A1(n_351), .A2(n_417), .B1(n_429), .B2(n_433), .C1(n_435), .C2(n_439), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B(n_357), .C(n_360), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_354), .B(n_398), .Y(n_421) );
INVx1_ASAP7_75t_L g443 ( .A(n_356), .Y(n_443) );
INVx1_ASAP7_75t_L g377 ( .A(n_358), .Y(n_377) );
OR2x2_ASAP7_75t_L g442 ( .A(n_359), .B(n_443), .Y(n_442) );
OAI21xp33_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_363), .B(n_367), .Y(n_360) );
NAND3xp33_ASAP7_75t_L g378 ( .A(n_361), .B(n_379), .C(n_380), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_361), .A2(n_398), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_365), .Y(n_418) );
AND2x2_ASAP7_75t_SL g384 ( .A(n_366), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g475 ( .A(n_366), .Y(n_475) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_366), .Y(n_491) );
INVx2_ASAP7_75t_L g449 ( .A(n_367), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_371), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g423 ( .A(n_373), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B1(n_378), .B2(n_382), .C(n_383), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_377), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_SL g511 ( .A(n_377), .Y(n_511) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g392 ( .A(n_384), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_384), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g450 ( .A(n_384), .B(n_398), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_384), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g483 ( .A(n_384), .B(n_418), .Y(n_483) );
BUFx3_ASAP7_75t_L g446 ( .A(n_385), .Y(n_446) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND5xp2_ASAP7_75t_L g388 ( .A(n_389), .B(n_407), .C(n_428), .D(n_440), .E(n_455), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI32xp33_ASAP7_75t_L g480 ( .A1(n_392), .A2(n_419), .A3(n_435), .B1(n_481), .B2(n_483), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_394), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g404 ( .A(n_398), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_402), .B1(n_404), .B2(n_405), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_414), .B1(n_416), .B2(n_417), .C(n_420), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g479 ( .A(n_411), .B(n_430), .Y(n_479) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_416), .A2(n_477), .B1(n_495), .B2(n_500), .C(n_501), .Y(n_494) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx2_ASAP7_75t_L g460 ( .A(n_419), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B1(n_424), .B2(n_426), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g438 ( .A(n_430), .Y(n_438) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_444), .B1(n_448), .B2(n_449), .C1(n_450), .C2(n_451), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_449), .A2(n_496), .B1(n_498), .B2(n_499), .Y(n_495) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_458), .B(n_461), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI21xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_466), .B(n_468), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g509 ( .A(n_464), .Y(n_509) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_476), .B(n_478), .C(n_480), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AOI211xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_488), .C(n_513), .Y(n_484) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_485), .Y(n_489) );
INVxp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI211xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_494), .C(n_506), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AOI21xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_504), .B(n_505), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_510), .B1(n_511), .B2(n_512), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AOI21xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_517), .Y(n_513) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_524), .Y(n_520) );
INVx1_ASAP7_75t_L g534 ( .A(n_521), .Y(n_534) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
endmodule