module fake_jpeg_4360_n_77 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_8),
.B(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_1),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_53),
.B1(n_38),
.B2(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_2),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_55),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_45),
.B1(n_36),
.B2(n_43),
.Y(n_64)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_57),
.B1(n_60),
.B2(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_64),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_62),
.C(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_35),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_66),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_70),
.B(n_64),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_71),
.A2(n_59),
.B(n_15),
.C(n_18),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_13),
.B(n_21),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_25),
.B(n_27),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_33),
.Y(n_77)
);


endmodule