module fake_netlist_1_1108_n_1395 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1395);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1395;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_533;
wire n_1010;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_659;
wire n_432;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1390;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g343 ( .A(n_74), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_98), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_237), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_325), .Y(n_346) );
INVxp33_ASAP7_75t_SL g347 ( .A(n_48), .Y(n_347) );
INVxp67_ASAP7_75t_SL g348 ( .A(n_44), .Y(n_348) );
INVxp67_ASAP7_75t_SL g349 ( .A(n_224), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_137), .Y(n_350) );
CKINVDCx16_ASAP7_75t_R g351 ( .A(n_88), .Y(n_351) );
INVxp67_ASAP7_75t_SL g352 ( .A(n_226), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_232), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_229), .Y(n_354) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_220), .Y(n_355) );
INVxp33_ASAP7_75t_L g356 ( .A(n_333), .Y(n_356) );
NOR2xp67_ASAP7_75t_L g357 ( .A(n_276), .B(n_102), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_277), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_216), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_42), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_194), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_40), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_298), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_263), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_107), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_234), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_288), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_70), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_179), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_66), .Y(n_370) );
CKINVDCx16_ASAP7_75t_R g371 ( .A(n_19), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_144), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_160), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_329), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_38), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_334), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_135), .Y(n_377) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_341), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_173), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_73), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_174), .Y(n_381) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_311), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_46), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_191), .Y(n_384) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_183), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_327), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_7), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_134), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_274), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_176), .Y(n_390) );
BUFx2_ASAP7_75t_SL g391 ( .A(n_72), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_293), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_273), .Y(n_393) );
BUFx3_ASAP7_75t_L g394 ( .A(n_31), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_193), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_147), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_19), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_188), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_342), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_331), .Y(n_400) );
INVxp33_ASAP7_75t_L g401 ( .A(n_38), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_324), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_233), .B(n_121), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_150), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_119), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_225), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_256), .Y(n_407) );
INVxp33_ASAP7_75t_L g408 ( .A(n_209), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_279), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_4), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_94), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_207), .B(n_208), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_236), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_62), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_51), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_257), .Y(n_416) );
INVxp33_ASAP7_75t_L g417 ( .A(n_243), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_81), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_154), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_162), .Y(n_420) );
CKINVDCx16_ASAP7_75t_R g421 ( .A(n_300), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_20), .Y(n_422) );
CKINVDCx16_ASAP7_75t_R g423 ( .A(n_286), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_275), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_303), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_5), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_6), .Y(n_427) );
CKINVDCx16_ASAP7_75t_R g428 ( .A(n_136), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_142), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_56), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_248), .Y(n_431) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_211), .Y(n_432) );
CKINVDCx16_ASAP7_75t_R g433 ( .A(n_250), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_41), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_187), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_45), .Y(n_436) );
CKINVDCx16_ASAP7_75t_R g437 ( .A(n_3), .Y(n_437) );
INVxp67_ASAP7_75t_SL g438 ( .A(n_164), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_269), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_109), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_210), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_172), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_88), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_18), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_111), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_238), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_266), .Y(n_447) );
BUFx5_ASAP7_75t_L g448 ( .A(n_181), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_301), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_34), .Y(n_450) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_13), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_204), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_268), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_136), .Y(n_454) );
NOR2xp67_ASAP7_75t_L g455 ( .A(n_282), .B(n_240), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_56), .B(n_152), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_337), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_156), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_170), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_21), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_217), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_143), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_206), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_51), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_114), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_221), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_27), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_184), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_192), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_104), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_280), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_171), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_205), .Y(n_473) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_45), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_272), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_93), .Y(n_476) );
INVxp33_ASAP7_75t_L g477 ( .A(n_69), .Y(n_477) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_163), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_72), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_95), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_200), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_259), .Y(n_482) );
INVxp33_ASAP7_75t_SL g483 ( .A(n_134), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_319), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_147), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_267), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_261), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_131), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_228), .Y(n_489) );
INVxp67_ASAP7_75t_SL g490 ( .A(n_219), .Y(n_490) );
INVxp33_ASAP7_75t_L g491 ( .A(n_107), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_58), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_44), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_306), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_96), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_201), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_161), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_52), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_53), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_190), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_10), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_339), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_93), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_145), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_58), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_28), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_84), .Y(n_507) );
INVxp67_ASAP7_75t_SL g508 ( .A(n_336), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_242), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_43), .Y(n_510) );
INVxp33_ASAP7_75t_SL g511 ( .A(n_29), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_335), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_223), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_130), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_199), .Y(n_515) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_81), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_10), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_264), .Y(n_518) );
INVxp67_ASAP7_75t_L g519 ( .A(n_37), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_12), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_32), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_245), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_299), .Y(n_523) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_457), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_386), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_351), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_526) );
NOR2xp33_ASAP7_75t_SL g527 ( .A(n_355), .B(n_148), .Y(n_527) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_386), .A2(n_0), .B(n_1), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_457), .Y(n_529) );
BUFx3_ASAP7_75t_L g530 ( .A(n_400), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_389), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_457), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_401), .B(n_2), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_389), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_401), .B(n_3), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_390), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_469), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_457), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_390), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_421), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_517), .B(n_4), .Y(n_541) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_457), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_356), .B(n_5), .Y(n_543) );
INVxp67_ASAP7_75t_L g544 ( .A(n_523), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_477), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_489), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_522), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_522), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_418), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_489), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_477), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_489), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_418), .Y(n_553) );
OA21x2_ASAP7_75t_L g554 ( .A1(n_407), .A2(n_6), .B(n_7), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_506), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_506), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_489), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_489), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_394), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_356), .B(n_8), .Y(n_560) );
INVx6_ASAP7_75t_L g561 ( .A(n_448), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_448), .Y(n_562) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_400), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_410), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_545), .B(n_408), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_562), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_545), .B(n_408), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_524), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_551), .B(n_417), .Y(n_569) );
INVx3_ASAP7_75t_L g570 ( .A(n_561), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_551), .Y(n_571) );
OAI21xp33_ASAP7_75t_L g572 ( .A1(n_525), .A2(n_417), .B(n_491), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_524), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_537), .B(n_491), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_537), .B(n_393), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_527), .A2(n_483), .B1(n_511), .B2(n_347), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_562), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_562), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_562), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_525), .B(n_345), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_524), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_533), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_561), .Y(n_583) );
INVx4_ASAP7_75t_L g584 ( .A(n_561), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_524), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_561), .Y(n_586) );
BUFx2_ASAP7_75t_L g587 ( .A(n_533), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_525), .B(n_407), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_561), .Y(n_589) );
INVx4_ASAP7_75t_L g590 ( .A(n_561), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_524), .Y(n_591) );
BUFx8_ASAP7_75t_SL g592 ( .A(n_540), .Y(n_592) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_524), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_544), .B(n_423), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_534), .B(n_346), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_534), .B(n_517), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_534), .B(n_394), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_531), .B(n_459), .Y(n_598) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_524), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_533), .B(n_371), .Y(n_600) );
BUFx3_ASAP7_75t_L g601 ( .A(n_530), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_524), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_544), .B(n_433), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_554), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_531), .B(n_459), .Y(n_605) );
INVx4_ASAP7_75t_L g606 ( .A(n_554), .Y(n_606) );
INVx4_ASAP7_75t_L g607 ( .A(n_554), .Y(n_607) );
BUFx5_ASAP7_75t_L g608 ( .A(n_604), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_606), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_582), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_606), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_571), .B(n_535), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_587), .B(n_535), .Y(n_613) );
INVx5_ASAP7_75t_L g614 ( .A(n_584), .Y(n_614) );
A2O1A1Ixp33_ASAP7_75t_L g615 ( .A1(n_572), .A2(n_536), .B(n_547), .C(n_539), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_587), .B(n_535), .Y(n_616) );
BUFx4f_ASAP7_75t_L g617 ( .A(n_600), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_594), .A2(n_527), .B1(n_560), .B2(n_540), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_594), .A2(n_560), .B1(n_543), .B2(n_483), .Y(n_619) );
INVx3_ASAP7_75t_L g620 ( .A(n_596), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_575), .B(n_536), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_587), .B(n_539), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_594), .A2(n_543), .B1(n_511), .B2(n_347), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_582), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_594), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_606), .B(n_547), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_596), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_596), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_606), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_596), .Y(n_630) );
AND2x4_ASAP7_75t_L g631 ( .A(n_565), .B(n_541), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_596), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_565), .B(n_548), .Y(n_633) );
INVx5_ASAP7_75t_L g634 ( .A(n_584), .Y(n_634) );
INVx5_ASAP7_75t_L g635 ( .A(n_584), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_601), .Y(n_636) );
BUFx5_ASAP7_75t_L g637 ( .A(n_604), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_603), .A2(n_379), .B1(n_381), .B2(n_364), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_565), .B(n_548), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_574), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_565), .B(n_530), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_567), .B(n_541), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_606), .A2(n_554), .B1(n_528), .B2(n_559), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_596), .Y(n_644) );
INVx3_ASAP7_75t_L g645 ( .A(n_597), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_567), .B(n_530), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g647 ( .A(n_603), .B(n_526), .C(n_437), .Y(n_647) );
INVxp33_ASAP7_75t_L g648 ( .A(n_574), .Y(n_648) );
OR2x6_ASAP7_75t_L g649 ( .A(n_600), .B(n_526), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_606), .B(n_441), .Y(n_650) );
BUFx12f_ASAP7_75t_SL g651 ( .A(n_574), .Y(n_651) );
INVx2_ASAP7_75t_SL g652 ( .A(n_567), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_601), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_592), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_597), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_597), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_571), .Y(n_657) );
OR2x6_ASAP7_75t_L g658 ( .A(n_600), .B(n_391), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_607), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_600), .B(n_428), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_607), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_567), .B(n_530), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_603), .Y(n_663) );
NOR2xp67_ASAP7_75t_L g664 ( .A(n_576), .B(n_559), .Y(n_664) );
BUFx2_ASAP7_75t_L g665 ( .A(n_603), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g666 ( .A1(n_576), .A2(n_516), .B1(n_505), .B2(n_364), .Y(n_666) );
INVx3_ASAP7_75t_L g667 ( .A(n_597), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_569), .B(n_379), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_597), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_572), .A2(n_553), .B(n_555), .C(n_549), .Y(n_670) );
BUFx4f_ASAP7_75t_L g671 ( .A(n_569), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_597), .Y(n_672) );
BUFx3_ASAP7_75t_L g673 ( .A(n_601), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_569), .A2(n_381), .B1(n_360), .B2(n_370), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_607), .Y(n_675) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_607), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_572), .A2(n_362), .B1(n_375), .B2(n_370), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_607), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_607), .B(n_354), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_588), .Y(n_680) );
INVx1_ASAP7_75t_SL g681 ( .A(n_592), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_576), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_588), .Y(n_683) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_604), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_575), .B(n_362), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_671), .A2(n_598), .B1(n_595), .B2(n_580), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_666), .A2(n_595), .B1(n_580), .B2(n_444), .C(n_422), .Y(n_687) );
INVx2_ASAP7_75t_SL g688 ( .A(n_671), .Y(n_688) );
INVx2_ASAP7_75t_SL g689 ( .A(n_680), .Y(n_689) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_684), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_647), .A2(n_598), .B1(n_595), .B2(n_580), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_684), .Y(n_692) );
BUFx3_ASAP7_75t_L g693 ( .A(n_673), .Y(n_693) );
INVx3_ASAP7_75t_L g694 ( .A(n_645), .Y(n_694) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_684), .Y(n_695) );
AND2x4_ASAP7_75t_L g696 ( .A(n_652), .B(n_605), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_631), .B(n_605), .Y(n_697) );
INVx1_ASAP7_75t_SL g698 ( .A(n_657), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_683), .A2(n_422), .B1(n_444), .B2(n_350), .Y(n_699) );
INVx3_ASAP7_75t_L g700 ( .A(n_645), .Y(n_700) );
BUFx5_ASAP7_75t_L g701 ( .A(n_655), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_631), .A2(n_350), .B1(n_577), .B2(n_566), .Y(n_702) );
NAND2x1p5_ASAP7_75t_L g703 ( .A(n_667), .B(n_554), .Y(n_703) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_684), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_642), .B(n_566), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_642), .B(n_566), .Y(n_706) );
NOR2xp67_ASAP7_75t_L g707 ( .A(n_638), .B(n_375), .Y(n_707) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_636), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_612), .B(n_554), .Y(n_709) );
INVx4_ASAP7_75t_L g710 ( .A(n_614), .Y(n_710) );
BUFx4f_ASAP7_75t_L g711 ( .A(n_658), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_667), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_627), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_624), .A2(n_578), .B1(n_579), .B2(n_577), .Y(n_714) );
BUFx2_ASAP7_75t_L g715 ( .A(n_651), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_676), .Y(n_716) );
INVx3_ASAP7_75t_L g717 ( .A(n_673), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_676), .Y(n_718) );
BUFx3_ASAP7_75t_L g719 ( .A(n_636), .Y(n_719) );
INVx4_ASAP7_75t_L g720 ( .A(n_614), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_676), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_625), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_676), .Y(n_723) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_636), .Y(n_724) );
BUFx2_ASAP7_75t_SL g725 ( .A(n_625), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_608), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_630), .Y(n_727) );
AND2x4_ASAP7_75t_L g728 ( .A(n_658), .B(n_348), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_613), .B(n_577), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_632), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_644), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_608), .Y(n_732) );
INVx3_ASAP7_75t_L g733 ( .A(n_620), .Y(n_733) );
BUFx3_ASAP7_75t_L g734 ( .A(n_636), .Y(n_734) );
INVx3_ASAP7_75t_SL g735 ( .A(n_654), .Y(n_735) );
BUFx2_ASAP7_75t_L g736 ( .A(n_663), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_616), .B(n_578), .Y(n_737) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_614), .Y(n_738) );
AND2x4_ASAP7_75t_L g739 ( .A(n_658), .B(n_368), .Y(n_739) );
INVx3_ASAP7_75t_L g740 ( .A(n_620), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_663), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_656), .Y(n_742) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_634), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_608), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_608), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_624), .B(n_578), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_681), .Y(n_747) );
INVxp67_ASAP7_75t_SL g748 ( .A(n_668), .Y(n_748) );
NOR3xp33_ASAP7_75t_L g749 ( .A(n_666), .B(n_519), .C(n_470), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_665), .A2(n_377), .B1(n_397), .B2(n_380), .Y(n_750) );
BUFx2_ASAP7_75t_SL g751 ( .A(n_640), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_669), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_672), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_608), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_648), .B(n_377), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_617), .Y(n_756) );
INVx2_ASAP7_75t_SL g757 ( .A(n_617), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_621), .B(n_579), .Y(n_758) );
INVx4_ASAP7_75t_L g759 ( .A(n_634), .Y(n_759) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_634), .Y(n_760) );
BUFx10_ASAP7_75t_L g761 ( .A(n_610), .Y(n_761) );
AND2x4_ASAP7_75t_L g762 ( .A(n_664), .B(n_451), .Y(n_762) );
AND2x4_ASAP7_75t_L g763 ( .A(n_633), .B(n_474), .Y(n_763) );
BUFx2_ASAP7_75t_L g764 ( .A(n_608), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_647), .B(n_586), .C(n_583), .Y(n_765) );
OAI21x1_ASAP7_75t_SL g766 ( .A1(n_670), .A2(n_528), .B(n_456), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_637), .Y(n_767) );
AND2x4_ASAP7_75t_L g768 ( .A(n_639), .B(n_549), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_622), .B(n_380), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_637), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_619), .B(n_397), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_628), .B(n_553), .Y(n_772) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_634), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_649), .A2(n_528), .B1(n_391), .B2(n_344), .Y(n_774) );
INVx3_ASAP7_75t_L g775 ( .A(n_628), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_649), .A2(n_528), .B1(n_365), .B2(n_372), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_641), .Y(n_777) );
INVx2_ASAP7_75t_SL g778 ( .A(n_637), .Y(n_778) );
BUFx2_ASAP7_75t_L g779 ( .A(n_637), .Y(n_779) );
BUFx3_ASAP7_75t_L g780 ( .A(n_635), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_648), .B(n_528), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_637), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_637), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_674), .B(n_528), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_646), .Y(n_785) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_660), .Y(n_786) );
INVxp67_ASAP7_75t_L g787 ( .A(n_685), .Y(n_787) );
AOI22xp33_ASAP7_75t_SL g788 ( .A1(n_682), .A2(n_460), .B1(n_495), .B2(n_440), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_662), .Y(n_789) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_635), .Y(n_790) );
NAND2x1p5_ASAP7_75t_L g791 ( .A(n_635), .B(n_626), .Y(n_791) );
OAI21xp5_ASAP7_75t_L g792 ( .A1(n_626), .A2(n_586), .B(n_583), .Y(n_792) );
AOI21x1_ASAP7_75t_L g793 ( .A1(n_679), .A2(n_586), .B(n_583), .Y(n_793) );
AND2x4_ASAP7_75t_L g794 ( .A(n_649), .B(n_555), .Y(n_794) );
BUFx8_ASAP7_75t_L g795 ( .A(n_609), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_623), .A2(n_460), .B1(n_495), .B2(n_440), .Y(n_796) );
INVxp67_ASAP7_75t_L g797 ( .A(n_650), .Y(n_797) );
AND2x4_ASAP7_75t_L g798 ( .A(n_618), .B(n_556), .Y(n_798) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_650), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g800 ( .A1(n_679), .A2(n_590), .B(n_584), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_677), .Y(n_801) );
INVx3_ASAP7_75t_L g802 ( .A(n_635), .Y(n_802) );
INVx4_ASAP7_75t_L g803 ( .A(n_711), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_794), .A2(n_611), .B1(n_629), .B2(n_609), .Y(n_804) );
AOI221xp5_ASAP7_75t_L g805 ( .A1(n_687), .A2(n_670), .B1(n_615), .B2(n_405), .C(n_411), .Y(n_805) );
BUFx3_ASAP7_75t_L g806 ( .A(n_795), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_689), .Y(n_807) );
INVx3_ASAP7_75t_L g808 ( .A(n_710), .Y(n_808) );
BUFx6f_ASAP7_75t_L g809 ( .A(n_690), .Y(n_809) );
O2A1O1Ixp33_ASAP7_75t_SL g810 ( .A1(n_778), .A2(n_615), .B(n_359), .C(n_361), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_698), .B(n_507), .Y(n_811) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_702), .A2(n_507), .B1(n_629), .B2(n_611), .Y(n_812) );
INVx3_ASAP7_75t_L g813 ( .A(n_710), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_794), .A2(n_659), .B1(n_675), .B2(n_661), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_697), .B(n_659), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_689), .Y(n_816) );
INVx1_ASAP7_75t_SL g817 ( .A(n_725), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_697), .B(n_678), .Y(n_818) );
BUFx6f_ASAP7_75t_L g819 ( .A(n_690), .Y(n_819) );
BUFx12f_ASAP7_75t_L g820 ( .A(n_747), .Y(n_820) );
BUFx2_ASAP7_75t_L g821 ( .A(n_741), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_794), .A2(n_678), .B1(n_643), .B2(n_434), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_696), .B(n_643), .Y(n_823) );
OAI22xp5_ASAP7_75t_SL g824 ( .A1(n_741), .A2(n_373), .B1(n_413), .B2(n_384), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_772), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_690), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_690), .Y(n_827) );
AOI221xp5_ASAP7_75t_L g828 ( .A1(n_749), .A2(n_414), .B1(n_415), .B2(n_396), .C(n_343), .Y(n_828) );
INVx6_ASAP7_75t_L g829 ( .A(n_795), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_758), .A2(n_456), .B1(n_403), .B2(n_653), .Y(n_830) );
OAI222xp33_ASAP7_75t_L g831 ( .A1(n_699), .A2(n_403), .B1(n_387), .B2(n_436), .C1(n_383), .C2(n_388), .Y(n_831) );
OR2x6_ASAP7_75t_L g832 ( .A(n_757), .B(n_383), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_695), .Y(n_833) );
OR2x2_ASAP7_75t_L g834 ( .A(n_722), .B(n_556), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_772), .Y(n_835) );
NAND2x1p5_ASAP7_75t_L g836 ( .A(n_711), .B(n_584), .Y(n_836) );
NOR2xp33_ASAP7_75t_R g837 ( .A(n_756), .B(n_373), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_784), .A2(n_434), .B1(n_410), .B2(n_427), .Y(n_838) );
BUFx3_ASAP7_75t_L g839 ( .A(n_795), .Y(n_839) );
OAI22xp5_ASAP7_75t_SL g840 ( .A1(n_788), .A2(n_413), .B1(n_425), .B2(n_384), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_784), .A2(n_434), .B1(n_410), .B2(n_429), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_772), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_798), .A2(n_410), .B1(n_434), .B2(n_430), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g844 ( .A1(n_748), .A2(n_425), .B1(n_446), .B2(n_431), .Y(n_844) );
NAND3xp33_ASAP7_75t_SL g845 ( .A(n_747), .B(n_446), .C(n_431), .Y(n_845) );
BUFx10_ASAP7_75t_L g846 ( .A(n_728), .Y(n_846) );
BUFx10_ASAP7_75t_L g847 ( .A(n_728), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_787), .B(n_388), .Y(n_848) );
CKINVDCx6p67_ASAP7_75t_R g849 ( .A(n_735), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_768), .Y(n_850) );
OR2x2_ASAP7_75t_L g851 ( .A(n_722), .B(n_436), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_768), .Y(n_852) );
AOI21xp5_ASAP7_75t_SL g853 ( .A1(n_778), .A2(n_352), .B(n_349), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_801), .B(n_584), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_786), .B(n_426), .Y(n_855) );
AOI22xp33_ASAP7_75t_SL g856 ( .A1(n_736), .A2(n_494), .B1(n_458), .B2(n_445), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_695), .Y(n_857) );
INVx4_ASAP7_75t_L g858 ( .A(n_738), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_695), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_746), .A2(n_402), .B1(n_374), .B2(n_378), .Y(n_860) );
OR2x2_ASAP7_75t_L g861 ( .A(n_736), .B(n_443), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_695), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_696), .A2(n_382), .B1(n_385), .B2(n_353), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_735), .Y(n_864) );
CKINVDCx5p33_ASAP7_75t_R g865 ( .A(n_715), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_715), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_704), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_798), .A2(n_434), .B1(n_410), .B2(n_450), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_798), .A2(n_763), .B1(n_765), .B2(n_777), .Y(n_869) );
AOI21xp5_ASAP7_75t_L g870 ( .A1(n_800), .A2(n_590), .B(n_589), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_768), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_704), .Y(n_872) );
BUFx6f_ASAP7_75t_L g873 ( .A(n_704), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_756), .Y(n_874) );
AOI222xp33_ASAP7_75t_L g875 ( .A1(n_707), .A2(n_454), .B1(n_462), .B2(n_467), .C1(n_465), .C2(n_464), .Y(n_875) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_764), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g877 ( .A1(n_801), .A2(n_479), .B1(n_480), .B2(n_476), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_691), .B(n_485), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g879 ( .A1(n_755), .A2(n_493), .B1(n_498), .B2(n_492), .C(n_488), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_704), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_705), .Y(n_881) );
BUFx3_ASAP7_75t_L g882 ( .A(n_738), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_703), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_706), .A2(n_432), .B1(n_478), .B2(n_438), .Y(n_884) );
INVx3_ASAP7_75t_L g885 ( .A(n_710), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_716), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_785), .A2(n_501), .B1(n_503), .B2(n_499), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_686), .A2(n_490), .B1(n_508), .B2(n_504), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_789), .A2(n_514), .B1(n_520), .B2(n_510), .Y(n_889) );
OR2x2_ASAP7_75t_L g890 ( .A(n_750), .B(n_521), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_709), .A2(n_563), .B1(n_358), .B2(n_366), .Y(n_891) );
BUFx12f_ASAP7_75t_L g892 ( .A(n_728), .Y(n_892) );
OAI22xp33_ASAP7_75t_L g893 ( .A1(n_729), .A2(n_357), .B1(n_367), .B2(n_363), .Y(n_893) );
INVx4_ASAP7_75t_L g894 ( .A(n_738), .Y(n_894) );
OAI21xp5_ASAP7_75t_L g895 ( .A1(n_792), .A2(n_589), .B(n_570), .Y(n_895) );
OR2x6_ASAP7_75t_L g896 ( .A(n_757), .B(n_751), .Y(n_896) );
NOR4xp25_ASAP7_75t_L g897 ( .A(n_774), .B(n_564), .C(n_376), .D(n_395), .Y(n_897) );
AOI221xp5_ASAP7_75t_L g898 ( .A1(n_769), .A2(n_762), .B1(n_771), .B2(n_739), .C(n_796), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_739), .A2(n_448), .B1(n_392), .B2(n_398), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_762), .A2(n_563), .B1(n_399), .B2(n_404), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_762), .A2(n_563), .B1(n_406), .B2(n_409), .Y(n_901) );
OAI21x1_ASAP7_75t_L g902 ( .A1(n_793), .A2(n_515), .B(n_512), .Y(n_902) );
CKINVDCx11_ASAP7_75t_R g903 ( .A(n_761), .Y(n_903) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_761), .A2(n_448), .B1(n_416), .B2(n_419), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_761), .B(n_8), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_688), .B(n_590), .Y(n_906) );
AOI221xp5_ASAP7_75t_L g907 ( .A1(n_742), .A2(n_420), .B1(n_435), .B2(n_424), .C(n_369), .Y(n_907) );
AOI22xp33_ASAP7_75t_SL g908 ( .A1(n_688), .A2(n_448), .B1(n_439), .B2(n_447), .Y(n_908) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_764), .Y(n_909) );
AND2x4_ASAP7_75t_L g910 ( .A(n_720), .B(n_590), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_752), .Y(n_911) );
CKINVDCx16_ASAP7_75t_R g912 ( .A(n_780), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_716), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_737), .B(n_590), .Y(n_914) );
BUFx3_ASAP7_75t_L g915 ( .A(n_738), .Y(n_915) );
BUFx3_ASAP7_75t_L g916 ( .A(n_743), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_781), .A2(n_563), .B1(n_442), .B2(n_452), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_718), .Y(n_918) );
AOI22xp33_ASAP7_75t_SL g919 ( .A1(n_779), .A2(n_448), .B1(n_453), .B2(n_449), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_714), .B(n_590), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_713), .B(n_461), .Y(n_921) );
AOI22xp5_ASAP7_75t_SL g922 ( .A1(n_797), .A2(n_412), .B1(n_466), .B2(n_463), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_753), .A2(n_472), .B1(n_473), .B2(n_471), .C(n_468), .Y(n_923) );
OAI221xp5_ASAP7_75t_L g924 ( .A1(n_776), .A2(n_481), .B1(n_484), .B2(n_482), .C(n_475), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_779), .A2(n_486), .B1(n_496), .B2(n_487), .Y(n_925) );
INVx4_ASAP7_75t_SL g926 ( .A(n_743), .Y(n_926) );
OA21x2_ASAP7_75t_L g927 ( .A1(n_766), .A2(n_515), .B(n_512), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_718), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_781), .A2(n_563), .B1(n_497), .B2(n_502), .Y(n_929) );
OAI221xp5_ASAP7_75t_L g930 ( .A1(n_799), .A2(n_509), .B1(n_518), .B2(n_513), .C(n_500), .Y(n_930) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_694), .B(n_570), .Y(n_931) );
INVxp33_ASAP7_75t_L g932 ( .A(n_837), .Y(n_932) );
OAI22xp33_ASAP7_75t_L g933 ( .A1(n_832), .A2(n_727), .B1(n_731), .B2(n_730), .Y(n_933) );
OAI22xp33_ASAP7_75t_L g934 ( .A1(n_832), .A2(n_732), .B1(n_744), .B2(n_726), .Y(n_934) );
AOI21xp33_ASAP7_75t_L g935 ( .A1(n_830), .A2(n_802), .B(n_766), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_911), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_881), .B(n_898), .Y(n_937) );
OR2x2_ASAP7_75t_L g938 ( .A(n_912), .B(n_720), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_834), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_869), .A2(n_701), .B1(n_712), .B2(n_694), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_832), .A2(n_812), .B1(n_869), .B2(n_822), .Y(n_941) );
OAI21xp5_ASAP7_75t_L g942 ( .A1(n_822), .A2(n_793), .B(n_791), .Y(n_942) );
INVx2_ASAP7_75t_SL g943 ( .A(n_829), .Y(n_943) );
OAI22xp33_ASAP7_75t_L g944 ( .A1(n_806), .A2(n_745), .B1(n_767), .B2(n_754), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_839), .B(n_759), .Y(n_945) );
OR2x6_ASAP7_75t_L g946 ( .A(n_839), .B(n_759), .Y(n_946) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_821), .B(n_694), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_886), .Y(n_948) );
BUFx2_ASAP7_75t_L g949 ( .A(n_892), .Y(n_949) );
AOI221xp5_ASAP7_75t_L g950 ( .A1(n_828), .A2(n_700), .B1(n_740), .B2(n_775), .C(n_733), .Y(n_950) );
OAI21xp5_ASAP7_75t_L g951 ( .A1(n_897), .A2(n_791), .B(n_723), .Y(n_951) );
INVx4_ASAP7_75t_L g952 ( .A(n_903), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_875), .A2(n_701), .B1(n_700), .B2(n_733), .Y(n_953) );
AOI221xp5_ASAP7_75t_L g954 ( .A1(n_831), .A2(n_700), .B1(n_740), .B2(n_775), .C(n_733), .Y(n_954) );
OR2x6_ASAP7_75t_L g955 ( .A(n_803), .B(n_743), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_805), .A2(n_701), .B1(n_775), .B2(n_740), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_886), .Y(n_957) );
OAI222xp33_ASAP7_75t_L g958 ( .A1(n_896), .A2(n_802), .B1(n_791), .B2(n_783), .C1(n_782), .C2(n_745), .Y(n_958) );
OAI21xp33_ASAP7_75t_L g959 ( .A1(n_843), .A2(n_780), .B(n_693), .Y(n_959) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_864), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_823), .A2(n_692), .B(n_754), .Y(n_961) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_840), .A2(n_701), .B1(n_802), .B2(n_760), .Y(n_962) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_849), .Y(n_963) );
OAI21x1_ASAP7_75t_L g964 ( .A1(n_902), .A2(n_692), .B(n_767), .Y(n_964) );
OAI221xp5_ASAP7_75t_L g965 ( .A1(n_877), .A2(n_717), .B1(n_693), .B2(n_723), .C(n_721), .Y(n_965) );
AOI221xp5_ASAP7_75t_L g966 ( .A1(n_879), .A2(n_717), .B1(n_773), .B2(n_760), .C(n_743), .Y(n_966) );
AND2x2_ASAP7_75t_L g967 ( .A(n_811), .B(n_760), .Y(n_967) );
OAI211xp5_ASAP7_75t_L g968 ( .A1(n_856), .A2(n_455), .B(n_564), .C(n_532), .Y(n_968) );
BUFx6f_ASAP7_75t_L g969 ( .A(n_809), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_887), .B(n_760), .Y(n_970) );
NOR2xp33_ASAP7_75t_L g971 ( .A(n_824), .B(n_773), .Y(n_971) );
BUFx2_ASAP7_75t_L g972 ( .A(n_896), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_815), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_850), .A2(n_790), .B1(n_773), .B2(n_734), .Y(n_974) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_803), .A2(n_782), .B1(n_783), .B2(n_770), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_843), .A2(n_770), .B1(n_734), .B2(n_719), .Y(n_976) );
AOI22xp5_ASAP7_75t_L g977 ( .A1(n_854), .A2(n_790), .B1(n_719), .B2(n_724), .Y(n_977) );
OAI222xp33_ASAP7_75t_L g978 ( .A1(n_930), .A2(n_564), .B1(n_11), .B2(n_12), .C1(n_13), .C2(n_14), .Y(n_978) );
AOI222xp33_ASAP7_75t_L g979 ( .A1(n_848), .A2(n_563), .B1(n_529), .B2(n_550), .C1(n_558), .C2(n_557), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_818), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_889), .B(n_708), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_852), .A2(n_563), .B1(n_448), .B2(n_708), .Y(n_982) );
AO22x1_ASAP7_75t_L g983 ( .A1(n_905), .A2(n_724), .B1(n_708), .B2(n_15), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_871), .A2(n_563), .B1(n_724), .B2(n_708), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_851), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_921), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_868), .A2(n_532), .B1(n_538), .B2(n_529), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_878), .A2(n_532), .B1(n_538), .B2(n_529), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_855), .B(n_9), .Y(n_989) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_868), .A2(n_538), .B1(n_546), .B2(n_529), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_861), .A2(n_546), .B1(n_557), .B2(n_550), .Y(n_991) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_876), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_893), .A2(n_546), .B1(n_557), .B2(n_550), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_846), .B(n_11), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_893), .A2(n_550), .B1(n_558), .B2(n_557), .Y(n_995) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_907), .A2(n_558), .B1(n_570), .B2(n_552), .C(n_542), .Y(n_996) );
INVx4_ASAP7_75t_L g997 ( .A(n_926), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_825), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_876), .A2(n_558), .B1(n_570), .B2(n_552), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_890), .B(n_15), .Y(n_1000) );
OAI22xp5_ASAP7_75t_SL g1001 ( .A1(n_820), .A2(n_18), .B1(n_16), .B2(n_17), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_854), .A2(n_552), .B1(n_542), .B2(n_568), .Y(n_1002) );
OAI221xp5_ASAP7_75t_L g1003 ( .A1(n_817), .A2(n_570), .B1(n_542), .B2(n_552), .C(n_591), .Y(n_1003) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_909), .A2(n_552), .B1(n_542), .B2(n_20), .Y(n_1004) );
AO21x2_ASAP7_75t_L g1005 ( .A1(n_810), .A2(n_573), .B(n_568), .Y(n_1005) );
OAI22xp33_ASAP7_75t_L g1006 ( .A1(n_909), .A2(n_552), .B1(n_542), .B2(n_21), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_923), .A2(n_552), .B1(n_542), .B2(n_568), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_838), .A2(n_841), .B1(n_891), .B2(n_924), .Y(n_1008) );
OAI221xp5_ASAP7_75t_L g1009 ( .A1(n_863), .A2(n_542), .B1(n_552), .B2(n_602), .C(n_591), .Y(n_1009) );
AOI222xp33_ASAP7_75t_L g1010 ( .A1(n_884), .A2(n_542), .B1(n_17), .B2(n_22), .C1(n_23), .C2(n_24), .Y(n_1010) );
OAI33xp33_ASAP7_75t_L g1011 ( .A1(n_888), .A2(n_602), .A3(n_591), .B1(n_585), .B2(n_581), .B3(n_573), .Y(n_1011) );
AOI211xp5_ASAP7_75t_L g1012 ( .A1(n_860), .A2(n_581), .B(n_585), .C(n_573), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_835), .Y(n_1013) );
AOI221xp5_ASAP7_75t_L g1014 ( .A1(n_838), .A2(n_602), .B1(n_591), .B2(n_585), .C(n_581), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_841), .A2(n_585), .B1(n_602), .B2(n_581), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_842), .B(n_16), .Y(n_1016) );
AOI21xp5_ASAP7_75t_L g1017 ( .A1(n_810), .A2(n_599), .B(n_593), .Y(n_1017) );
A2O1A1Ixp33_ASAP7_75t_L g1018 ( .A1(n_807), .A2(n_599), .B(n_593), .C(n_24), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1019 ( .A(n_865), .B(n_22), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_844), .B(n_23), .Y(n_1020) );
AND2x4_ASAP7_75t_SL g1021 ( .A(n_846), .B(n_25), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_900), .A2(n_599), .B1(n_593), .B2(n_27), .Y(n_1022) );
AOI21xp5_ASAP7_75t_L g1023 ( .A1(n_870), .A2(n_599), .B(n_593), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_900), .A2(n_599), .B1(n_593), .B2(n_28), .Y(n_1024) );
INVx2_ASAP7_75t_L g1025 ( .A(n_913), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_901), .A2(n_599), .B1(n_593), .B2(n_29), .Y(n_1026) );
CKINVDCx10_ASAP7_75t_R g1027 ( .A(n_874), .Y(n_1027) );
AOI21xp5_ASAP7_75t_L g1028 ( .A1(n_883), .A2(n_827), .B(n_826), .Y(n_1028) );
OR2x2_ASAP7_75t_L g1029 ( .A(n_845), .B(n_26), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_816), .Y(n_1030) );
AOI221xp5_ASAP7_75t_L g1031 ( .A1(n_925), .A2(n_599), .B1(n_593), .B2(n_30), .C(n_31), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_901), .A2(n_599), .B1(n_593), .B2(n_30), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_847), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_899), .A2(n_599), .B1(n_593), .B2(n_35), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_837), .B(n_33), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_922), .B(n_34), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_913), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_918), .Y(n_1038) );
OAI22xp33_ASAP7_75t_L g1039 ( .A1(n_836), .A2(n_37), .B1(n_35), .B2(n_36), .Y(n_1039) );
AOI21xp5_ASAP7_75t_L g1040 ( .A1(n_883), .A2(n_151), .B(n_149), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_917), .A2(n_40), .B1(n_36), .B2(n_39), .Y(n_1041) );
INVx1_ASAP7_75t_SL g1042 ( .A(n_866), .Y(n_1042) );
BUFx3_ASAP7_75t_L g1043 ( .A(n_882), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_929), .A2(n_49), .B1(n_47), .B2(n_48), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_918), .Y(n_1045) );
AOI22xp33_ASAP7_75t_SL g1046 ( .A1(n_927), .A2(n_52), .B1(n_49), .B2(n_50), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1047 ( .A1(n_920), .A2(n_54), .B1(n_50), .B2(n_53), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_928), .Y(n_1048) );
AOI221xp5_ASAP7_75t_L g1049 ( .A1(n_853), .A2(n_55), .B1(n_57), .B2(n_59), .C(n_60), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_858), .B(n_55), .Y(n_1050) );
OAI22xp33_ASAP7_75t_L g1051 ( .A1(n_933), .A2(n_927), .B1(n_813), .B2(n_885), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_989), .B(n_858), .Y(n_1052) );
OAI22xp5_ASAP7_75t_SL g1053 ( .A1(n_963), .A2(n_927), .B1(n_904), .B2(n_894), .Y(n_1053) );
INVx1_ASAP7_75t_SL g1054 ( .A(n_1027), .Y(n_1054) );
OAI21xp5_ASAP7_75t_SL g1055 ( .A1(n_932), .A2(n_919), .B(n_908), .Y(n_1055) );
AOI33xp33_ASAP7_75t_L g1056 ( .A1(n_1036), .A2(n_804), .A3(n_814), .B1(n_60), .B2(n_61), .B3(n_62), .Y(n_1056) );
AO21x2_ASAP7_75t_L g1057 ( .A1(n_942), .A2(n_895), .B(n_827), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_941), .A2(n_808), .B1(n_885), .B2(n_813), .Y(n_1058) );
OAI221xp5_ASAP7_75t_SL g1059 ( .A1(n_1041), .A2(n_804), .B1(n_814), .B2(n_808), .C(n_931), .Y(n_1059) );
OR2x6_ASAP7_75t_L g1060 ( .A(n_946), .B(n_894), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_936), .Y(n_1061) );
CKINVDCx5p33_ASAP7_75t_R g1062 ( .A(n_960), .Y(n_1062) );
INVx2_ASAP7_75t_L g1063 ( .A(n_948), .Y(n_1063) );
OAI21xp5_ASAP7_75t_L g1064 ( .A1(n_1008), .A2(n_914), .B(n_931), .Y(n_1064) );
HB1xp67_ASAP7_75t_L g1065 ( .A(n_992), .Y(n_1065) );
INVx3_ASAP7_75t_L g1066 ( .A(n_997), .Y(n_1066) );
AO21x2_ASAP7_75t_L g1067 ( .A1(n_935), .A2(n_833), .B(n_826), .Y(n_1067) );
AOI22xp33_ASAP7_75t_SL g1068 ( .A1(n_1001), .A2(n_915), .B1(n_916), .B2(n_882), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_937), .A2(n_928), .B1(n_916), .B2(n_915), .Y(n_1069) );
NAND4xp25_ASAP7_75t_L g1070 ( .A(n_1019), .B(n_906), .C(n_910), .D(n_61), .Y(n_1070) );
BUFx2_ASAP7_75t_L g1071 ( .A(n_946), .Y(n_1071) );
AOI221xp5_ASAP7_75t_L g1072 ( .A1(n_985), .A2(n_910), .B1(n_906), .B2(n_833), .C(n_857), .Y(n_1072) );
NOR4xp25_ASAP7_75t_L g1073 ( .A(n_1039), .B(n_63), .C(n_57), .D(n_59), .Y(n_1073) );
AOI21x1_ASAP7_75t_L g1074 ( .A1(n_983), .A2(n_859), .B(n_857), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1030), .Y(n_1075) );
INVx2_ASAP7_75t_L g1076 ( .A(n_957), .Y(n_1076) );
AO21x2_ASAP7_75t_L g1077 ( .A1(n_951), .A2(n_867), .B(n_862), .Y(n_1077) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1025), .Y(n_1078) );
INVx2_ASAP7_75t_L g1079 ( .A(n_1037), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_939), .Y(n_1080) );
BUFx6f_ASAP7_75t_L g1081 ( .A(n_969), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_933), .A2(n_819), .B1(n_873), .B2(n_809), .Y(n_1082) );
AOI22xp33_ASAP7_75t_SL g1083 ( .A1(n_972), .A2(n_819), .B1(n_873), .B2(n_809), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1084 ( .A(n_938), .B(n_973), .Y(n_1084) );
NAND4xp25_ASAP7_75t_L g1085 ( .A(n_1010), .B(n_66), .C(n_64), .D(n_65), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_980), .B(n_986), .Y(n_1086) );
INVx2_ASAP7_75t_L g1087 ( .A(n_1038), .Y(n_1087) );
AOI22xp5_ASAP7_75t_L g1088 ( .A1(n_953), .A2(n_926), .B1(n_880), .B2(n_872), .Y(n_1088) );
INVx1_ASAP7_75t_SL g1089 ( .A(n_1042), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_945), .B(n_64), .Y(n_1090) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_955), .B(n_880), .Y(n_1091) );
AOI221xp5_ASAP7_75t_L g1092 ( .A1(n_978), .A2(n_873), .B1(n_819), .B2(n_68), .C(n_69), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_1000), .A2(n_68), .B1(n_65), .B2(n_67), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_998), .Y(n_1094) );
OAI222xp33_ASAP7_75t_L g1095 ( .A1(n_1039), .A2(n_67), .B1(n_70), .B2(n_71), .C1(n_73), .C2(n_74), .Y(n_1095) );
OAI21x1_ASAP7_75t_L g1096 ( .A1(n_964), .A2(n_155), .B(n_153), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1035), .B(n_71), .Y(n_1097) );
AO21x2_ASAP7_75t_L g1098 ( .A1(n_1005), .A2(n_75), .B(n_76), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1013), .Y(n_1099) );
INVx1_ASAP7_75t_SL g1100 ( .A(n_949), .Y(n_1100) );
AND2x4_ASAP7_75t_L g1101 ( .A(n_955), .B(n_157), .Y(n_1101) );
AND2x4_ASAP7_75t_L g1102 ( .A(n_955), .B(n_158), .Y(n_1102) );
OAI21xp5_ASAP7_75t_L g1103 ( .A1(n_1004), .A2(n_75), .B(n_76), .Y(n_1103) );
OAI221xp5_ASAP7_75t_L g1104 ( .A1(n_947), .A2(n_77), .B1(n_78), .B2(n_79), .C(n_80), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g1105 ( .A1(n_1006), .A2(n_78), .B1(n_79), .B2(n_80), .C(n_82), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_967), .B(n_83), .Y(n_1106) );
AO21x2_ASAP7_75t_L g1107 ( .A1(n_1005), .A2(n_83), .B(n_84), .Y(n_1107) );
OAI211xp5_ASAP7_75t_L g1108 ( .A1(n_1049), .A2(n_85), .B(n_86), .C(n_87), .Y(n_1108) );
INVx2_ASAP7_75t_SL g1109 ( .A(n_946), .Y(n_1109) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1045), .Y(n_1110) );
INVx2_ASAP7_75t_L g1111 ( .A(n_1048), .Y(n_1111) );
AOI221xp5_ASAP7_75t_L g1112 ( .A1(n_1006), .A2(n_85), .B1(n_86), .B2(n_87), .C(n_89), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_992), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1021), .B(n_90), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_994), .B(n_91), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1029), .Y(n_1116) );
OAI221xp5_ASAP7_75t_L g1117 ( .A1(n_1020), .A2(n_92), .B1(n_95), .B2(n_96), .C(n_97), .Y(n_1117) );
AOI33xp33_ASAP7_75t_L g1118 ( .A1(n_1044), .A2(n_97), .A3(n_98), .B1(n_99), .B2(n_100), .B3(n_101), .Y(n_1118) );
OAI321xp33_ASAP7_75t_L g1119 ( .A1(n_1044), .A2(n_103), .A3(n_104), .B1(n_105), .B2(n_106), .C(n_108), .Y(n_1119) );
OAI33xp33_ASAP7_75t_L g1120 ( .A1(n_1047), .A2(n_103), .A3(n_105), .B1(n_106), .B2(n_108), .B3(n_109), .Y(n_1120) );
OAI21xp5_ASAP7_75t_L g1121 ( .A1(n_956), .A2(n_110), .B(n_111), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1016), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1050), .Y(n_1123) );
NOR2xp33_ASAP7_75t_L g1124 ( .A(n_1033), .B(n_112), .Y(n_1124) );
OAI211xp5_ASAP7_75t_L g1125 ( .A1(n_991), .A2(n_112), .B(n_113), .C(n_114), .Y(n_1125) );
OA21x2_ASAP7_75t_L g1126 ( .A1(n_1023), .A2(n_165), .B(n_159), .Y(n_1126) );
OA21x2_ASAP7_75t_L g1127 ( .A1(n_1017), .A2(n_167), .B(n_166), .Y(n_1127) );
OA21x2_ASAP7_75t_L g1128 ( .A1(n_1028), .A2(n_169), .B(n_168), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_970), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_943), .B(n_113), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_971), .B(n_115), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_952), .B(n_115), .Y(n_1132) );
NAND3xp33_ASAP7_75t_L g1133 ( .A(n_1046), .B(n_968), .C(n_979), .Y(n_1133) );
AOI33xp33_ASAP7_75t_L g1134 ( .A1(n_993), .A2(n_116), .A3(n_117), .B1(n_118), .B2(n_119), .B3(n_120), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_981), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1043), .B(n_116), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_987), .Y(n_1137) );
OR2x2_ASAP7_75t_L g1138 ( .A(n_993), .B(n_117), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_995), .B(n_118), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_954), .B(n_120), .Y(n_1140) );
AOI22xp33_ASAP7_75t_SL g1141 ( .A1(n_965), .A2(n_121), .B1(n_122), .B2(n_123), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_990), .Y(n_1142) );
AOI22xp5_ASAP7_75t_L g1143 ( .A1(n_956), .A2(n_124), .B1(n_125), .B2(n_126), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_950), .B(n_127), .Y(n_1144) );
INVx2_ASAP7_75t_SL g1145 ( .A(n_969), .Y(n_1145) );
AOI222xp33_ASAP7_75t_L g1146 ( .A1(n_1031), .A2(n_127), .B1(n_128), .B2(n_129), .C1(n_130), .C2(n_132), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_962), .B(n_128), .Y(n_1147) );
OAI221xp5_ASAP7_75t_L g1148 ( .A1(n_940), .A2(n_133), .B1(n_135), .B2(n_137), .C(n_138), .Y(n_1148) );
OAI321xp33_ASAP7_75t_L g1149 ( .A1(n_1034), .A2(n_138), .A3(n_139), .B1(n_140), .B2(n_141), .C(n_142), .Y(n_1149) );
AOI21x1_ASAP7_75t_L g1150 ( .A1(n_961), .A2(n_146), .B(n_340), .Y(n_1150) );
OAI21xp5_ASAP7_75t_SL g1151 ( .A1(n_958), .A2(n_175), .B(n_177), .Y(n_1151) );
BUFx2_ASAP7_75t_L g1152 ( .A(n_944), .Y(n_1152) );
OR2x2_ASAP7_75t_L g1153 ( .A(n_1022), .B(n_1024), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_1024), .A2(n_178), .B1(n_180), .B2(n_182), .Y(n_1154) );
INVx2_ASAP7_75t_L g1155 ( .A(n_1063), .Y(n_1155) );
OAI221xp5_ASAP7_75t_L g1156 ( .A1(n_1070), .A2(n_1034), .B1(n_1032), .B2(n_1026), .C(n_966), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1061), .Y(n_1157) );
AO31x2_ASAP7_75t_L g1158 ( .A1(n_1082), .A2(n_1018), .A3(n_976), .B(n_1040), .Y(n_1158) );
OAI33xp33_ASAP7_75t_L g1159 ( .A1(n_1116), .A2(n_934), .A3(n_944), .B1(n_975), .B2(n_999), .B3(n_959), .Y(n_1159) );
AOI33xp33_ASAP7_75t_L g1160 ( .A1(n_1080), .A2(n_1032), .A3(n_1026), .B1(n_988), .B2(n_1007), .B3(n_1002), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1075), .Y(n_1161) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1063), .Y(n_1162) );
OAI21xp5_ASAP7_75t_L g1163 ( .A1(n_1085), .A2(n_1009), .B(n_1002), .Y(n_1163) );
INVx3_ASAP7_75t_L g1164 ( .A(n_1081), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1086), .B(n_974), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1079), .B(n_969), .Y(n_1166) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1076), .Y(n_1167) );
INVx3_ASAP7_75t_L g1168 ( .A(n_1081), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1094), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1099), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_1058), .A2(n_977), .B1(n_984), .B2(n_1007), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1087), .B(n_1110), .Y(n_1172) );
INVxp67_ASAP7_75t_SL g1173 ( .A(n_1065), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_1153), .A2(n_1011), .B1(n_996), .B2(n_1003), .Y(n_1174) );
INVx2_ASAP7_75t_SL g1175 ( .A(n_1060), .Y(n_1175) );
AOI221xp5_ASAP7_75t_L g1176 ( .A1(n_1073), .A2(n_982), .B1(n_1012), .B2(n_1015), .C(n_1014), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1084), .B(n_1015), .Y(n_1177) );
AOI21x1_ASAP7_75t_L g1178 ( .A1(n_1074), .A2(n_185), .B(n_186), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1110), .B(n_189), .Y(n_1179) );
HB1xp67_ASAP7_75t_L g1180 ( .A(n_1111), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1113), .Y(n_1181) );
INVxp67_ASAP7_75t_L g1182 ( .A(n_1100), .Y(n_1182) );
NOR2xp67_ASAP7_75t_L g1183 ( .A(n_1151), .B(n_195), .Y(n_1183) );
AND2x4_ASAP7_75t_L g1184 ( .A(n_1129), .B(n_196), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1135), .B(n_197), .Y(n_1185) );
OAI31xp33_ASAP7_75t_SL g1186 ( .A1(n_1068), .A2(n_198), .A3(n_202), .B(n_203), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1076), .Y(n_1187) );
HB1xp67_ASAP7_75t_L g1188 ( .A(n_1078), .Y(n_1188) );
OR2x2_ASAP7_75t_L g1189 ( .A(n_1123), .B(n_1089), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1056), .B(n_338), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1078), .Y(n_1191) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1081), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1058), .B(n_212), .Y(n_1193) );
OAI31xp33_ASAP7_75t_L g1194 ( .A1(n_1095), .A2(n_213), .A3(n_214), .B(n_215), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1152), .B(n_218), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1056), .B(n_222), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1134), .Y(n_1197) );
NAND2x1p5_ASAP7_75t_L g1198 ( .A(n_1101), .B(n_227), .Y(n_1198) );
AOI22xp5_ASAP7_75t_L g1199 ( .A1(n_1124), .A2(n_230), .B1(n_231), .B2(n_235), .Y(n_1199) );
NAND3xp33_ASAP7_75t_SL g1200 ( .A(n_1054), .B(n_239), .C(n_241), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1106), .B(n_244), .Y(n_1201) );
NAND3xp33_ASAP7_75t_L g1202 ( .A(n_1118), .B(n_246), .C(n_247), .Y(n_1202) );
HB1xp67_ASAP7_75t_L g1203 ( .A(n_1052), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1090), .B(n_249), .Y(n_1204) );
NAND3xp33_ASAP7_75t_L g1205 ( .A(n_1118), .B(n_251), .C(n_252), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1134), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_1144), .A2(n_253), .B1(n_254), .B2(n_255), .Y(n_1207) );
OAI31xp33_ASAP7_75t_L g1208 ( .A1(n_1108), .A2(n_258), .A3(n_260), .B(n_262), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_1120), .A2(n_265), .B1(n_270), .B2(n_271), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1130), .Y(n_1210) );
NAND3xp33_ASAP7_75t_L g1211 ( .A(n_1093), .B(n_278), .C(n_281), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1136), .Y(n_1212) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1081), .Y(n_1213) );
AND2x4_ASAP7_75t_L g1214 ( .A(n_1109), .B(n_283), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1122), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1131), .Y(n_1216) );
AND2x4_ASAP7_75t_L g1217 ( .A(n_1109), .B(n_284), .Y(n_1217) );
AOI33xp33_ASAP7_75t_L g1218 ( .A1(n_1132), .A2(n_285), .A3(n_287), .B1(n_289), .B2(n_290), .B3(n_291), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1071), .Y(n_1219) );
AND2x4_ASAP7_75t_L g1220 ( .A(n_1145), .B(n_292), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1057), .B(n_294), .Y(n_1221) );
BUFx2_ASAP7_75t_L g1222 ( .A(n_1060), .Y(n_1222) );
AOI211xp5_ASAP7_75t_L g1223 ( .A1(n_1104), .A2(n_295), .B(n_296), .C(n_297), .Y(n_1223) );
NAND3xp33_ASAP7_75t_L g1224 ( .A(n_1093), .B(n_302), .C(n_304), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1077), .B(n_305), .Y(n_1225) );
NOR2xp33_ASAP7_75t_L g1226 ( .A(n_1124), .B(n_307), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1147), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1098), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1115), .B(n_308), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1098), .Y(n_1230) );
INVx5_ASAP7_75t_L g1231 ( .A(n_1101), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1097), .B(n_309), .Y(n_1232) );
OAI221xp5_ASAP7_75t_SL g1233 ( .A1(n_1117), .A2(n_310), .B1(n_312), .B2(n_313), .C(n_314), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1107), .Y(n_1234) );
AOI21xp5_ASAP7_75t_L g1235 ( .A1(n_1051), .A2(n_315), .B(n_316), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1107), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_1120), .A2(n_317), .B1(n_318), .B2(n_320), .Y(n_1237) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1067), .Y(n_1238) );
CKINVDCx16_ASAP7_75t_R g1239 ( .A(n_1203), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_1197), .A2(n_1092), .B1(n_1141), .B2(n_1112), .Y(n_1240) );
NOR3xp33_ASAP7_75t_L g1241 ( .A(n_1200), .B(n_1119), .C(n_1149), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1157), .Y(n_1242) );
AND2x4_ASAP7_75t_L g1243 ( .A(n_1231), .B(n_1067), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1215), .B(n_1068), .Y(n_1244) );
NAND3xp33_ASAP7_75t_L g1245 ( .A(n_1186), .B(n_1105), .C(n_1146), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1161), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1169), .Y(n_1247) );
OAI31xp33_ASAP7_75t_L g1248 ( .A1(n_1226), .A2(n_1114), .A3(n_1125), .B(n_1148), .Y(n_1248) );
HB1xp67_ASAP7_75t_L g1249 ( .A(n_1180), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1181), .B(n_1064), .Y(n_1250) );
OR2x6_ASAP7_75t_L g1251 ( .A(n_1198), .B(n_1101), .Y(n_1251) );
INVx2_ASAP7_75t_L g1252 ( .A(n_1155), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1170), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1173), .B(n_1069), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1172), .B(n_1069), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1227), .B(n_1139), .Y(n_1256) );
AND2x4_ASAP7_75t_L g1257 ( .A(n_1231), .B(n_1102), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1216), .B(n_1172), .Y(n_1258) );
AND2x2_ASAP7_75t_SL g1259 ( .A(n_1214), .B(n_1102), .Y(n_1259) );
NOR2xp33_ASAP7_75t_L g1260 ( .A(n_1210), .B(n_1059), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1188), .B(n_1088), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1189), .Y(n_1262) );
OAI221xp5_ASAP7_75t_SL g1263 ( .A1(n_1206), .A2(n_1055), .B1(n_1143), .B2(n_1140), .C(n_1138), .Y(n_1263) );
AND2x4_ASAP7_75t_L g1264 ( .A(n_1231), .B(n_1102), .Y(n_1264) );
INVx2_ASAP7_75t_L g1265 ( .A(n_1155), .Y(n_1265) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1162), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1187), .Y(n_1267) );
OAI221xp5_ASAP7_75t_L g1268 ( .A1(n_1182), .A2(n_1121), .B1(n_1053), .B2(n_1103), .C(n_1133), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1191), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1212), .B(n_1072), .Y(n_1270) );
INVx2_ASAP7_75t_SL g1271 ( .A(n_1231), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1219), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1162), .Y(n_1273) );
INVx2_ASAP7_75t_L g1274 ( .A(n_1167), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1166), .B(n_1083), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_1156), .A2(n_1142), .B1(n_1137), .B2(n_1154), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1228), .B(n_1066), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1230), .B(n_1083), .Y(n_1278) );
AOI33xp33_ASAP7_75t_L g1279 ( .A1(n_1209), .A2(n_1091), .A3(n_1062), .B1(n_1150), .B2(n_1126), .B3(n_326), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1165), .B(n_1091), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1234), .B(n_1091), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1177), .B(n_1126), .Y(n_1282) );
AND2x4_ASAP7_75t_L g1283 ( .A(n_1175), .B(n_1096), .Y(n_1283) );
HB1xp67_ASAP7_75t_L g1284 ( .A(n_1222), .Y(n_1284) );
OR2x6_ASAP7_75t_L g1285 ( .A(n_1198), .B(n_1096), .Y(n_1285) );
INVx2_ASAP7_75t_L g1286 ( .A(n_1238), .Y(n_1286) );
INVx2_ASAP7_75t_SL g1287 ( .A(n_1164), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1179), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1236), .B(n_1128), .Y(n_1289) );
AND4x1_ASAP7_75t_L g1290 ( .A(n_1218), .B(n_321), .C(n_322), .D(n_323), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1204), .B(n_1127), .Y(n_1291) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1238), .Y(n_1292) );
BUFx2_ASAP7_75t_L g1293 ( .A(n_1214), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1195), .Y(n_1294) );
AND2x4_ASAP7_75t_L g1295 ( .A(n_1192), .B(n_1213), .Y(n_1295) );
INVxp33_ASAP7_75t_L g1296 ( .A(n_1195), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1221), .B(n_1127), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1217), .Y(n_1298) );
AO211x2_ASAP7_75t_L g1299 ( .A1(n_1245), .A2(n_1205), .B(n_1202), .C(n_1163), .Y(n_1299) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_1239), .B(n_1192), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1249), .B(n_1213), .Y(n_1301) );
BUFx2_ASAP7_75t_L g1302 ( .A(n_1251), .Y(n_1302) );
NOR2xp33_ASAP7_75t_L g1303 ( .A(n_1260), .B(n_1159), .Y(n_1303) );
OAI22xp5_ASAP7_75t_L g1304 ( .A1(n_1259), .A2(n_1217), .B1(n_1183), .B2(n_1209), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1242), .Y(n_1305) );
OAI21xp33_ASAP7_75t_L g1306 ( .A1(n_1260), .A2(n_1218), .B(n_1237), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1246), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1247), .Y(n_1308) );
INVxp67_ASAP7_75t_L g1309 ( .A(n_1278), .Y(n_1309) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1262), .B(n_1164), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1253), .Y(n_1311) );
OAI332xp33_ASAP7_75t_L g1312 ( .A1(n_1268), .A2(n_1190), .A3(n_1196), .B1(n_1229), .B2(n_1171), .B3(n_1160), .C1(n_1194), .C2(n_1223), .Y(n_1312) );
INVx1_ASAP7_75t_SL g1313 ( .A(n_1258), .Y(n_1313) );
OAI221xp5_ASAP7_75t_L g1314 ( .A1(n_1248), .A2(n_1233), .B1(n_1207), .B2(n_1208), .C(n_1237), .Y(n_1314) );
OR2x2_ASAP7_75t_L g1315 ( .A(n_1280), .B(n_1168), .Y(n_1315) );
AND2x4_ASAP7_75t_L g1316 ( .A(n_1281), .B(n_1217), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1284), .B(n_1225), .Y(n_1317) );
AOI221x1_ASAP7_75t_L g1318 ( .A1(n_1241), .A2(n_1235), .B1(n_1184), .B2(n_1211), .C(n_1224), .Y(n_1318) );
OR2x2_ASAP7_75t_L g1319 ( .A(n_1272), .B(n_1168), .Y(n_1319) );
INVx3_ASAP7_75t_L g1320 ( .A(n_1251), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1255), .B(n_1275), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1267), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1250), .B(n_1225), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1269), .B(n_1158), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1255), .B(n_1201), .Y(n_1325) );
AND2x4_ASAP7_75t_L g1326 ( .A(n_1281), .B(n_1220), .Y(n_1326) );
NOR2xp33_ASAP7_75t_L g1327 ( .A(n_1244), .B(n_1232), .Y(n_1327) );
AND2x4_ASAP7_75t_L g1328 ( .A(n_1251), .B(n_1220), .Y(n_1328) );
A2O1A1Ixp33_ASAP7_75t_L g1329 ( .A1(n_1296), .A2(n_1193), .B(n_1160), .C(n_1199), .Y(n_1329) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1254), .B(n_1184), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1275), .B(n_1184), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1261), .B(n_1185), .Y(n_1332) );
AND2x2_ASAP7_75t_SL g1333 ( .A(n_1293), .B(n_1220), .Y(n_1333) );
BUFx2_ASAP7_75t_L g1334 ( .A(n_1251), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1309), .B(n_1278), .Y(n_1335) );
NOR2xp33_ASAP7_75t_L g1336 ( .A(n_1303), .B(n_1263), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1309), .B(n_1273), .Y(n_1337) );
OR2x2_ASAP7_75t_L g1338 ( .A(n_1313), .B(n_1277), .Y(n_1338) );
OAI221xp5_ASAP7_75t_L g1339 ( .A1(n_1303), .A2(n_1276), .B1(n_1270), .B2(n_1240), .C(n_1256), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1321), .B(n_1294), .Y(n_1340) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1305), .Y(n_1341) );
INVxp67_ASAP7_75t_L g1342 ( .A(n_1300), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1324), .B(n_1282), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1307), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1324), .B(n_1266), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1308), .Y(n_1346) );
AND2x2_ASAP7_75t_SL g1347 ( .A(n_1333), .B(n_1257), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1311), .Y(n_1348) );
INVxp67_ASAP7_75t_SL g1349 ( .A(n_1301), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1322), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1310), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1319), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1315), .Y(n_1353) );
AOI22xp5_ASAP7_75t_L g1354 ( .A1(n_1306), .A2(n_1264), .B1(n_1298), .B2(n_1297), .Y(n_1354) );
AND2x4_ASAP7_75t_L g1355 ( .A(n_1302), .B(n_1243), .Y(n_1355) );
XOR2x2_ASAP7_75t_L g1356 ( .A(n_1333), .B(n_1290), .Y(n_1356) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1334), .Y(n_1357) );
NAND4xp25_ASAP7_75t_L g1358 ( .A(n_1318), .B(n_1329), .C(n_1314), .D(n_1327), .Y(n_1358) );
A2O1A1Ixp33_ASAP7_75t_L g1359 ( .A1(n_1328), .A2(n_1264), .B(n_1279), .C(n_1271), .Y(n_1359) );
INVxp67_ASAP7_75t_L g1360 ( .A(n_1317), .Y(n_1360) );
AND2x4_ASAP7_75t_L g1361 ( .A(n_1320), .B(n_1243), .Y(n_1361) );
NOR2xp33_ASAP7_75t_L g1362 ( .A(n_1312), .B(n_1287), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1325), .B(n_1288), .Y(n_1363) );
AOI211xp5_ASAP7_75t_SL g1364 ( .A1(n_1304), .A2(n_1291), .B(n_1243), .C(n_1283), .Y(n_1364) );
INVxp67_ASAP7_75t_L g1365 ( .A(n_1330), .Y(n_1365) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_1299), .A2(n_1283), .B1(n_1285), .B2(n_1176), .Y(n_1366) );
INVx2_ASAP7_75t_L g1367 ( .A(n_1326), .Y(n_1367) );
OAI22xp5_ASAP7_75t_L g1368 ( .A1(n_1316), .A2(n_1265), .B1(n_1252), .B2(n_1274), .Y(n_1368) );
OAI211xp5_ASAP7_75t_L g1369 ( .A1(n_1323), .A2(n_1174), .B(n_1289), .C(n_1292), .Y(n_1369) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_1358), .A2(n_1336), .B1(n_1362), .B2(n_1366), .Y(n_1370) );
OAI31xp33_ASAP7_75t_L g1371 ( .A1(n_1364), .A2(n_1359), .A3(n_1369), .B(n_1339), .Y(n_1371) );
OAI21xp33_ASAP7_75t_L g1372 ( .A1(n_1335), .A2(n_1354), .B(n_1357), .Y(n_1372) );
INVx1_ASAP7_75t_SL g1373 ( .A(n_1338), .Y(n_1373) );
XNOR2xp5_ASAP7_75t_L g1374 ( .A(n_1356), .B(n_1347), .Y(n_1374) );
OAI21xp5_ASAP7_75t_L g1375 ( .A1(n_1349), .A2(n_1360), .B(n_1368), .Y(n_1375) );
NAND2xp5_ASAP7_75t_SL g1376 ( .A(n_1355), .B(n_1361), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1352), .B(n_1343), .Y(n_1377) );
NOR2xp67_ASAP7_75t_L g1378 ( .A(n_1374), .B(n_1342), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1377), .Y(n_1379) );
AO22x2_ASAP7_75t_L g1380 ( .A1(n_1373), .A2(n_1341), .B1(n_1350), .B2(n_1344), .Y(n_1380) );
AOI221xp5_ASAP7_75t_L g1381 ( .A1(n_1370), .A2(n_1348), .B1(n_1346), .B2(n_1365), .C(n_1353), .Y(n_1381) );
NAND4xp75_ASAP7_75t_L g1382 ( .A(n_1371), .B(n_1331), .C(n_1337), .D(n_1332), .Y(n_1382) );
NAND4xp25_ASAP7_75t_L g1383 ( .A(n_1378), .B(n_1375), .C(n_1372), .D(n_1376), .Y(n_1383) );
OR3x1_ASAP7_75t_L g1384 ( .A(n_1379), .B(n_1351), .C(n_1367), .Y(n_1384) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1380), .Y(n_1385) );
NOR3xp33_ASAP7_75t_L g1386 ( .A(n_1382), .B(n_1178), .C(n_1345), .Y(n_1386) );
AND3x1_ASAP7_75t_L g1387 ( .A(n_1381), .B(n_1340), .C(n_1363), .Y(n_1387) );
AND3x4_ASAP7_75t_L g1388 ( .A(n_1386), .B(n_1316), .C(n_1326), .Y(n_1388) );
INVx4_ASAP7_75t_L g1389 ( .A(n_1385), .Y(n_1389) );
NOR3xp33_ASAP7_75t_L g1390 ( .A(n_1389), .B(n_1383), .C(n_1387), .Y(n_1390) );
NAND2x1p5_ASAP7_75t_SL g1391 ( .A(n_1388), .B(n_1384), .Y(n_1391) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_1390), .A2(n_1295), .B1(n_1286), .B2(n_1265), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g1393 ( .A1(n_1392), .A2(n_1390), .B1(n_1391), .B2(n_1295), .Y(n_1393) );
HB1xp67_ASAP7_75t_L g1394 ( .A(n_1393), .Y(n_1394) );
AOI221xp5_ASAP7_75t_L g1395 ( .A1(n_1394), .A2(n_1158), .B1(n_328), .B2(n_330), .C(n_332), .Y(n_1395) );
endmodule