module real_jpeg_23862_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_286;
wire n_176;
wire n_288;
wire n_292;
wire n_166;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_197;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_184;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_258;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_0),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_0),
.A2(n_46),
.B1(n_69),
.B2(n_70),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_46),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_2),
.A2(n_62),
.B1(n_78),
.B2(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_2),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_2),
.A2(n_69),
.B1(n_70),
.B2(n_117),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_117),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_117),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_5),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_5),
.B(n_79),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_5),
.B(n_31),
.C(n_50),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_160),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_5),
.B(n_123),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_5),
.A2(n_95),
.B1(n_96),
.B2(n_232),
.Y(n_235)
);

INVx8_ASAP7_75t_SL g68 ( 
.A(n_6),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_55),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_7),
.A2(n_55),
.B1(n_69),
.B2(n_70),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_8),
.A2(n_32),
.B1(n_61),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_8),
.A2(n_32),
.B1(n_69),
.B2(n_70),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_8),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_9),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_9),
.A2(n_60),
.B1(n_69),
.B2(n_70),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_60),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_60),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_10),
.A2(n_35),
.B1(n_69),
.B2(n_70),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_10),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_10),
.A2(n_35),
.B1(n_78),
.B2(n_138),
.Y(n_137)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_11),
.B(n_69),
.C(n_72),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_13),
.A2(n_61),
.B1(n_63),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_13),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_13),
.A2(n_69),
.B1(n_70),
.B2(n_163),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_163),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_163),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_15),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_147),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_145),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_118),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_19),
.B(n_118),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_92),
.C(n_103),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_20),
.A2(n_21),
.B1(n_92),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_56),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_22),
.B(n_80),
.C(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_23),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_25),
.A2(n_95),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_27),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_29),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_29),
.A2(n_95),
.B(n_108),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_37),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_31),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_30),
.B(n_237),
.Y(n_236)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_33),
.A2(n_177),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_34),
.B(n_37),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_36),
.A2(n_107),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_36),
.A2(n_192),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_37),
.Y(n_233)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_38),
.Y(n_192)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_42),
.A2(n_52),
.B(n_110),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_44),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_44),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_43),
.A2(n_84),
.B(n_247),
.C(n_249),
.Y(n_246)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_44),
.B(n_207),
.Y(n_206)
);

NOR3xp33_ASAP7_75t_L g249 ( 
.A(n_44),
.B(n_69),
.C(n_83),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_47),
.B(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_47),
.A2(n_100),
.B(n_127),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_47),
.A2(n_53),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_47),
.A2(n_53),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_48),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_48),
.A2(n_52),
.B1(n_211),
.B2(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_48),
.A2(n_126),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_52),
.B(n_160),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_53),
.B(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_54),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_80),
.B1(n_81),
.B2(n_91),
.Y(n_56)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_64),
.B(n_75),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_59),
.A2(n_65),
.B1(n_79),
.B2(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_67),
.B1(n_72),
.B2(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_64),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_64),
.A2(n_66),
.B1(n_162),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_65),
.A2(n_79),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_73),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_67),
.A2(n_70),
.B(n_159),
.C(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_70),
.B1(n_83),
.B2(n_84),
.Y(n_88)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

HAxp5_ASAP7_75t_SL g248 ( 
.A(n_70),
.B(n_160),
.CON(n_248),
.SN(n_248)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_76),
.Y(n_135)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

HAxp5_ASAP7_75t_SL g159 ( 
.A(n_78),
.B(n_160),
.CON(n_159),
.SN(n_159)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_79),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B(n_86),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_82),
.A2(n_171),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_85),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_87),
.A2(n_123),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_87),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_87),
.A2(n_123),
.B1(n_197),
.B2(n_248),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_92),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_102),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_94),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_97),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_106),
.B(n_108),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_95),
.A2(n_225),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_103),
.B(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_112),
.C(n_115),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_104),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_109),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_112),
.B(n_115),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_113),
.B(n_123),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_116),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_118)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_129),
.B1(n_140),
.B2(n_141),
.Y(n_119)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_125),
.B(n_128),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_139),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_289),
.B(n_294),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_199),
.B(n_280),
.C(n_288),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_184),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_150),
.B(n_184),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_164),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_152),
.B(n_153),
.C(n_164),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.C(n_158),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_160),
.B(n_238),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_173),
.B2(n_183),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_167),
.B(n_169),
.C(n_183),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B(n_172),
.Y(n_169)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_181),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_175),
.B1(n_181),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_181),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_189),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_185),
.B(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_187),
.B(n_189),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_190),
.Y(n_265)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_195),
.B(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_279),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_274),
.B(n_278),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_259),
.B(n_273),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_242),
.B(n_258),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_221),
.B(n_241),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_212),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_208),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_213),
.B(n_216),
.C(n_219),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_214),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_220),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_228),
.B(n_240),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_227),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_234),
.B(n_239),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_231),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_257),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_257),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_253),
.C(n_254),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_250),
.B2(n_251),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_251),
.Y(n_268)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_256),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_261),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_269),
.C(n_271),
.Y(n_277)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_277),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.C(n_287),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);


endmodule