module fake_jpeg_27583_n_101 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_21),
.Y(n_28)
);

INVx5_ASAP7_75t_SL g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_29),
.B(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_6),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_5),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_18),
.B1(n_14),
.B2(n_16),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_38),
.B(n_42),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_20),
.B1(n_16),
.B2(n_23),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_20),
.B1(n_18),
.B2(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_24),
.A2(n_19),
.B1(n_13),
.B2(n_12),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_35),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_53),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_12),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_19),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_37),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_66),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_39),
.B1(n_42),
.B2(n_37),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_55),
.B1(n_39),
.B2(n_28),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_59),
.B1(n_61),
.B2(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_65),
.B(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

A2O1A1O1Ixp25_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_31),
.B(n_40),
.C(n_8),
.D(n_7),
.Y(n_81)
);

NOR2xp67_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_77),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_9),
.C(n_1),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_75),
.C(n_78),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_88),
.Y(n_92)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_89),
.A2(n_90),
.B1(n_81),
.B2(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_82),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_94),
.B(n_88),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_89),
.B(n_83),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_84),
.B1(n_74),
.B2(n_2),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_96),
.A2(n_0),
.B1(n_1),
.B2(n_92),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_0),
.B1(n_1),
.B2(n_97),
.C(n_99),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_0),
.Y(n_101)
);


endmodule