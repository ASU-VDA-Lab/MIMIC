module real_jpeg_5358_n_10 (n_8, n_0, n_73, n_2, n_76, n_9, n_79, n_78, n_75, n_6, n_7, n_3, n_77, n_5, n_4, n_81, n_1, n_74, n_80, n_10);

input n_8;
input n_0;
input n_73;
input n_2;
input n_76;
input n_9;
input n_79;
input n_78;
input n_75;
input n_6;
input n_7;
input n_3;
input n_77;
input n_5;
input n_4;
input n_81;
input n_1;
input n_74;
input n_80;

output n_10;

wire n_54;
wire n_37;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_67;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_57;
wire n_43;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_16;

INVx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_0),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_2),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_2),
.B(n_27),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_3),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_4),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_4),
.B(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_7),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_7),
.B(n_54),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_9),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_9),
.B(n_67),
.Y(n_69)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_22),
.B1(n_70),
.B2(n_71),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_21),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_17),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_17),
.B(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

OAI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_66),
.B(n_69),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_61),
.B(n_65),
.Y(n_23)
);

AO221x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.C(n_60),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AO21x1_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_42),
.B(n_57),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_41),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_53),
.B(n_56),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B(n_52),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_64),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_73),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_74),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_75),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_76),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_77),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_78),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_79),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_80),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_81),
.Y(n_68)
);


endmodule