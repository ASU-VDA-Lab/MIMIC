module fake_aes_272_n_868 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_115, n_97, n_80, n_107, n_60, n_114, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_113, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_868);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_113;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_868;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_638;
wire n_540;
wire n_563;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_822;
wire n_823;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g116 ( .A(n_36), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_15), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_89), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_41), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_51), .Y(n_120) );
BUFx2_ASAP7_75t_SL g121 ( .A(n_56), .Y(n_121) );
BUFx2_ASAP7_75t_L g122 ( .A(n_114), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_100), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_43), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_28), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_37), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_72), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_44), .Y(n_128) );
CKINVDCx16_ASAP7_75t_R g129 ( .A(n_53), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_30), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_42), .Y(n_131) );
OR2x2_ASAP7_75t_L g132 ( .A(n_107), .B(n_80), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_59), .Y(n_133) );
CKINVDCx14_ASAP7_75t_R g134 ( .A(n_98), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_115), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_12), .Y(n_136) );
INVxp67_ASAP7_75t_SL g137 ( .A(n_75), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_39), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_23), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_34), .B(n_111), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_82), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_60), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_105), .Y(n_143) );
INVx1_ASAP7_75t_SL g144 ( .A(n_109), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_76), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_65), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_102), .Y(n_147) );
INVxp33_ASAP7_75t_SL g148 ( .A(n_92), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_47), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_45), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_29), .Y(n_151) );
OR2x2_ASAP7_75t_L g152 ( .A(n_48), .B(n_70), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_85), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_61), .Y(n_154) );
INVx4_ASAP7_75t_R g155 ( .A(n_3), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_6), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_38), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_2), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_11), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_6), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_99), .Y(n_161) );
INVxp67_ASAP7_75t_SL g162 ( .A(n_1), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_83), .Y(n_163) );
CKINVDCx16_ASAP7_75t_R g164 ( .A(n_62), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_71), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_58), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_78), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_9), .Y(n_168) );
INVxp33_ASAP7_75t_L g169 ( .A(n_77), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_87), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_64), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_9), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_125), .Y(n_173) );
CKINVDCx8_ASAP7_75t_R g174 ( .A(n_129), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_122), .B(n_0), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_122), .B(n_0), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_125), .B(n_1), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_119), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_169), .B(n_2), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_128), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_127), .B(n_3), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_164), .B(n_4), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_146), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_128), .Y(n_184) );
INVx6_ASAP7_75t_L g185 ( .A(n_119), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_134), .B(n_4), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g187 ( .A(n_154), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_131), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_131), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_119), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_136), .B(n_5), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_119), .Y(n_192) );
AND2x6_ASAP7_75t_L g193 ( .A(n_170), .B(n_52), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_118), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_119), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_156), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_170), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_161), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_171), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_161), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_130), .B(n_7), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_118), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_177), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_175), .B(n_160), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_202), .B(n_124), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_198), .Y(n_206) );
BUFx10_ASAP7_75t_L g207 ( .A(n_194), .Y(n_207) );
NAND2xp33_ASAP7_75t_L g208 ( .A(n_193), .B(n_124), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_174), .A2(n_172), .B1(n_136), .B2(n_168), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_186), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_177), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_202), .B(n_148), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_177), .Y(n_213) );
BUFx10_ASAP7_75t_L g214 ( .A(n_193), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_183), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_177), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_177), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_174), .B(n_116), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_179), .B(n_133), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_191), .A2(n_168), .B1(n_172), .B2(n_117), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_187), .Y(n_221) );
BUFx2_ASAP7_75t_L g222 ( .A(n_186), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_180), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_193), .Y(n_224) );
INVx4_ASAP7_75t_L g225 ( .A(n_193), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_175), .A2(n_159), .B1(n_151), .B2(n_139), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_180), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_184), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_184), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_188), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_198), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_175), .B(n_160), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_193), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_179), .B(n_133), .Y(n_234) );
NOR2xp33_ASAP7_75t_SL g235 ( .A(n_174), .B(n_142), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_188), .B(n_120), .Y(n_236) );
NAND2xp33_ASAP7_75t_L g237 ( .A(n_193), .B(n_142), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_189), .Y(n_238) );
BUFx6f_ASAP7_75t_SL g239 ( .A(n_193), .Y(n_239) );
BUFx8_ASAP7_75t_SL g240 ( .A(n_182), .Y(n_240) );
INVx1_ASAP7_75t_SL g241 ( .A(n_182), .Y(n_241) );
BUFx10_ASAP7_75t_L g242 ( .A(n_193), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_189), .Y(n_243) );
BUFx2_ASAP7_75t_L g244 ( .A(n_186), .Y(n_244) );
INVx4_ASAP7_75t_L g245 ( .A(n_193), .Y(n_245) );
INVx4_ASAP7_75t_L g246 ( .A(n_198), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_198), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_197), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_215), .Y(n_249) );
NAND3xp33_ASAP7_75t_L g250 ( .A(n_208), .B(n_182), .C(n_179), .Y(n_250) );
AND2x4_ASAP7_75t_SL g251 ( .A(n_207), .B(n_158), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_219), .B(n_176), .Y(n_252) );
AND2x6_ASAP7_75t_L g253 ( .A(n_233), .B(n_191), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_203), .Y(n_254) );
OAI21xp33_ASAP7_75t_L g255 ( .A1(n_234), .A2(n_176), .B(n_191), .Y(n_255) );
NOR2xp33_ASAP7_75t_R g256 ( .A(n_221), .B(n_187), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_204), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_233), .Y(n_258) );
INVx5_ASAP7_75t_L g259 ( .A(n_246), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_204), .B(n_181), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_224), .B(n_197), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_203), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_223), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_211), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_224), .B(n_199), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_209), .A2(n_241), .B1(n_222), .B2(n_244), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_204), .B(n_199), .Y(n_267) );
NOR2xp33_ASAP7_75t_R g268 ( .A(n_235), .B(n_143), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_224), .B(n_132), .Y(n_269) );
NAND2x1p5_ASAP7_75t_L g270 ( .A(n_222), .B(n_132), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_204), .B(n_181), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_245), .B(n_152), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_232), .B(n_201), .Y(n_273) );
INVx4_ASAP7_75t_L g274 ( .A(n_225), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_210), .A2(n_201), .B1(n_173), .B2(n_162), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_232), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_223), .Y(n_277) );
NOR2x1_ASAP7_75t_L g278 ( .A(n_205), .B(n_152), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_210), .B(n_143), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_244), .B(n_211), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_213), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_227), .B(n_145), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_213), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_216), .B(n_173), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_240), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_227), .B(n_145), .Y(n_286) );
AND3x2_ASAP7_75t_SL g287 ( .A(n_207), .B(n_196), .C(n_155), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_216), .Y(n_288) );
NOR2xp33_ASAP7_75t_R g289 ( .A(n_207), .B(n_237), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_268), .B(n_245), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_260), .B(n_212), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_263), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_259), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_252), .B(n_207), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_260), .A2(n_217), .B1(n_220), .B2(n_226), .Y(n_295) );
NAND2x1p5_ASAP7_75t_L g296 ( .A(n_274), .B(n_225), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_259), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_260), .B(n_228), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_270), .B(n_217), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_251), .Y(n_300) );
AO32x2_ASAP7_75t_L g301 ( .A1(n_257), .A2(n_225), .A3(n_245), .B1(n_246), .B2(n_121), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_253), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_259), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_259), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_259), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_274), .Y(n_306) );
AND2x2_ASAP7_75t_SL g307 ( .A(n_251), .B(n_225), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_253), .Y(n_308) );
NOR2x1_ASAP7_75t_L g309 ( .A(n_250), .B(n_248), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_249), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_268), .B(n_214), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_274), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_271), .B(n_248), .Y(n_313) );
INVx4_ASAP7_75t_L g314 ( .A(n_253), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_280), .B(n_228), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_270), .B(n_196), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_266), .A2(n_230), .B1(n_243), .B2(n_229), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_263), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_253), .Y(n_319) );
OAI21xp33_ASAP7_75t_SL g320 ( .A1(n_254), .A2(n_230), .B(n_229), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_276), .A2(n_243), .B(n_238), .C(n_236), .Y(n_321) );
INVx4_ASAP7_75t_L g322 ( .A(n_253), .Y(n_322) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_255), .A2(n_238), .B(n_218), .C(n_171), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_279), .Y(n_324) );
A2O1A1Ixp33_ASAP7_75t_SL g325 ( .A1(n_294), .A2(n_275), .B(n_273), .C(n_277), .Y(n_325) );
OA21x2_ASAP7_75t_L g326 ( .A1(n_323), .A2(n_147), .B(n_153), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_321), .A2(n_278), .B(n_269), .Y(n_327) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_317), .A2(n_269), .B(n_272), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_320), .A2(n_318), .B(n_313), .C(n_277), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_318), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_299), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_295), .B(n_298), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_305), .Y(n_333) );
AO31x2_ASAP7_75t_L g334 ( .A1(n_292), .A2(n_283), .A3(n_288), .B(n_262), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_292), .Y(n_335) );
OAI21xp5_ASAP7_75t_L g336 ( .A1(n_309), .A2(n_264), .B(n_281), .Y(n_336) );
AO31x2_ASAP7_75t_L g337 ( .A1(n_315), .A2(n_178), .A3(n_200), .B(n_192), .Y(n_337) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_291), .A2(n_267), .B(n_272), .C(n_280), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_299), .B(n_280), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_309), .A2(n_135), .B(n_149), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_299), .B(n_284), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_299), .B(n_284), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_314), .Y(n_343) );
OAI21x1_ASAP7_75t_L g344 ( .A1(n_290), .A2(n_135), .B(n_149), .Y(n_344) );
AO21x2_ASAP7_75t_L g345 ( .A1(n_311), .A2(n_138), .B(n_123), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_305), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_297), .A2(n_130), .B(n_126), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_297), .A2(n_157), .B(n_141), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_305), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_306), .Y(n_350) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_324), .A2(n_192), .B(n_178), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_314), .Y(n_352) );
OR2x6_ASAP7_75t_L g353 ( .A(n_339), .B(n_314), .Y(n_353) );
INVx6_ASAP7_75t_L g354 ( .A(n_341), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_341), .B(n_316), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_332), .A2(n_316), .B1(n_307), .B2(n_284), .Y(n_356) );
OA21x2_ASAP7_75t_L g357 ( .A1(n_340), .A2(n_200), .B(n_178), .Y(n_357) );
OA21x2_ASAP7_75t_L g358 ( .A1(n_340), .A2(n_192), .B(n_200), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_339), .B(n_307), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_340), .A2(n_296), .B(n_297), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_332), .A2(n_256), .B1(n_285), .B2(n_300), .C(n_310), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_342), .A2(n_307), .B1(n_322), .B2(n_302), .Y(n_362) );
BUFx4f_ASAP7_75t_L g363 ( .A(n_343), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_329), .A2(n_261), .B(n_265), .Y(n_364) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_331), .A2(n_287), .B(n_173), .C(n_144), .Y(n_365) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_331), .A2(n_256), .B(n_300), .C(n_287), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_325), .A2(n_310), .B1(n_286), .B2(n_282), .C(n_302), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_342), .A2(n_322), .B1(n_319), .B2(n_308), .Y(n_368) );
A2O1A1Ixp33_ASAP7_75t_L g369 ( .A1(n_338), .A2(n_319), .B(n_308), .C(n_303), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g370 ( .A1(n_338), .A2(n_303), .B(n_304), .C(n_293), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_344), .A2(n_296), .B(n_312), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_341), .B(n_293), .Y(n_372) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_325), .A2(n_322), .B1(n_173), .B2(n_304), .C(n_306), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_330), .B(n_150), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_330), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_335), .B(n_306), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_334), .B(n_312), .Y(n_378) );
OA21x2_ASAP7_75t_L g379 ( .A1(n_344), .A2(n_137), .B(n_265), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g380 ( .A1(n_343), .A2(n_289), .B1(n_121), .B2(n_312), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_329), .A2(n_296), .B1(n_150), .B2(n_165), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_349), .B(n_165), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_328), .A2(n_289), .B1(n_161), .B2(n_163), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_337), .Y(n_384) );
OAI21x1_ASAP7_75t_L g385 ( .A1(n_344), .A2(n_261), .B(n_301), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_343), .A2(n_166), .B1(n_167), .B2(n_239), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_336), .A2(n_167), .B1(n_166), .B2(n_247), .C(n_231), .Y(n_387) );
INVx5_ASAP7_75t_SL g388 ( .A(n_346), .Y(n_388) );
CKINVDCx11_ASAP7_75t_R g389 ( .A(n_349), .Y(n_389) );
AOI22xp33_ASAP7_75t_SL g390 ( .A1(n_363), .A2(n_328), .B1(n_333), .B2(n_348), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_375), .B(n_334), .Y(n_391) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_363), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_376), .B(n_334), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_378), .B(n_334), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_375), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_384), .B(n_334), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_363), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_357), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_377), .Y(n_399) );
OA21x2_ASAP7_75t_L g400 ( .A1(n_370), .A2(n_347), .B(n_336), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_355), .B(n_334), .Y(n_401) );
NOR4xp25_ASAP7_75t_SL g402 ( .A(n_365), .B(n_326), .C(n_347), .D(n_348), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_388), .B(n_334), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_353), .B(n_346), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_382), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_370), .B(n_334), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_360), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_356), .A2(n_328), .B1(n_327), .B2(n_346), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_371), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_388), .B(n_346), .Y(n_411) );
NOR2x1_ASAP7_75t_SL g412 ( .A(n_353), .B(n_350), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_356), .A2(n_328), .B1(n_327), .B2(n_333), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_388), .B(n_328), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_371), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_385), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_357), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_353), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_353), .B(n_333), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_359), .B(n_327), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_385), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_372), .B(n_326), .Y(n_422) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_369), .A2(n_347), .B(n_348), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_374), .Y(n_424) );
BUFx3_ASAP7_75t_L g425 ( .A(n_389), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_354), .B(n_326), .Y(n_426) );
AO31x2_ASAP7_75t_L g427 ( .A1(n_381), .A2(n_350), .A3(n_326), .B(n_140), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_354), .B(n_326), .Y(n_428) );
INVxp67_ASAP7_75t_R g429 ( .A(n_389), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_357), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_358), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_354), .B(n_326), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_369), .B(n_350), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_358), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_368), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_383), .B(n_333), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_358), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_379), .Y(n_438) );
INVxp67_ASAP7_75t_L g439 ( .A(n_361), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_367), .A2(n_333), .B1(n_345), .B2(n_350), .Y(n_440) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_383), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_366), .B(n_351), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_379), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_379), .Y(n_444) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_364), .A2(n_345), .B(n_301), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_362), .B(n_351), .Y(n_446) );
AO21x2_ASAP7_75t_L g447 ( .A1(n_373), .A2(n_345), .B(n_301), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_387), .B(n_351), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_380), .Y(n_449) );
NAND2x1_ASAP7_75t_L g450 ( .A(n_386), .B(n_352), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_375), .B(n_352), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_375), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_363), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_378), .B(n_351), .Y(n_454) );
NOR2x1_ASAP7_75t_L g455 ( .A(n_425), .B(n_453), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_391), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_450), .A2(n_351), .B(n_345), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_391), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_394), .B(n_337), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_394), .B(n_337), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_398), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_395), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_452), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_398), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_399), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_399), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_396), .B(n_337), .Y(n_467) );
OAI31xp33_ASAP7_75t_L g468 ( .A1(n_439), .A2(n_352), .A3(n_10), .B(n_11), .Y(n_468) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_443), .A2(n_345), .B(n_301), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_396), .B(n_337), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_425), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_398), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_403), .B(n_337), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_393), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_393), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_424), .B(n_337), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g477 ( .A(n_405), .B(n_161), .C(n_163), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_407), .Y(n_478) );
OAI21x1_ASAP7_75t_L g479 ( .A1(n_444), .A2(n_352), .B(n_351), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_401), .B(n_337), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_417), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_417), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_403), .B(n_352), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_453), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_411), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_404), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_411), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_425), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_414), .B(n_161), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_431), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_401), .B(n_163), .Y(n_491) );
AO31x2_ASAP7_75t_L g492 ( .A1(n_406), .A2(n_301), .A3(n_190), .B(n_195), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_454), .B(n_163), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_431), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_454), .B(n_163), .Y(n_495) );
OAI21xp5_ASAP7_75t_SL g496 ( .A1(n_397), .A2(n_8), .B(n_10), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_417), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_437), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_449), .A2(n_239), .B1(n_185), .B2(n_214), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_422), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_414), .B(n_12), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_430), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_426), .B(n_13), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_426), .B(n_13), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_420), .B(n_14), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_428), .B(n_14), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_422), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_392), .B(n_15), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_420), .B(n_16), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_428), .B(n_16), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_432), .B(n_17), .Y(n_511) );
AND2x2_ASAP7_75t_SL g512 ( .A(n_436), .B(n_17), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_432), .B(n_18), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_409), .B(n_18), .Y(n_514) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_449), .A2(n_190), .B1(n_195), .B2(n_206), .C(n_231), .Y(n_515) );
NAND2xp33_ASAP7_75t_SL g516 ( .A(n_418), .B(n_239), .Y(n_516) );
INVx4_ASAP7_75t_L g517 ( .A(n_419), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_451), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_441), .B(n_19), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_443), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_406), .A2(n_190), .B1(n_195), .B2(n_206), .C(n_247), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_451), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_430), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_430), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_451), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_412), .Y(n_526) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_443), .A2(n_190), .B(n_195), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_413), .B(n_19), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_451), .Y(n_529) );
INVx4_ASAP7_75t_L g530 ( .A(n_419), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_404), .B(n_20), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_434), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_404), .B(n_20), .Y(n_533) );
OAI31xp33_ASAP7_75t_L g534 ( .A1(n_442), .A2(n_21), .A3(n_22), .B(n_23), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_434), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_407), .B(n_21), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_418), .B(n_22), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_444), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_444), .Y(n_539) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_434), .A2(n_190), .B(n_195), .Y(n_540) );
OAI31xp33_ASAP7_75t_L g541 ( .A1(n_442), .A2(n_24), .A3(n_25), .B(n_26), .Y(n_541) );
NAND2x1p5_ASAP7_75t_L g542 ( .A(n_418), .B(n_258), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_404), .B(n_24), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_444), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_438), .A2(n_190), .B1(n_195), .B2(n_246), .C(n_28), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_408), .B(n_25), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_416), .Y(n_547) );
INVxp67_ASAP7_75t_SL g548 ( .A(n_412), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_418), .B(n_26), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_408), .B(n_445), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g551 ( .A1(n_438), .A2(n_195), .B1(n_190), .B2(n_246), .C(n_27), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_445), .B(n_27), .Y(n_552) );
AOI33xp33_ASAP7_75t_L g553 ( .A1(n_390), .A2(n_29), .A3(n_185), .B1(n_32), .B2(n_33), .B3(n_35), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_419), .Y(n_554) );
INVx4_ASAP7_75t_L g555 ( .A(n_419), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_416), .Y(n_556) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_440), .A2(n_185), .B1(n_258), .B2(n_46), .C(n_49), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_410), .Y(n_558) );
NAND4xp25_ASAP7_75t_L g559 ( .A(n_446), .B(n_185), .C(n_40), .D(n_50), .Y(n_559) );
NOR3xp33_ASAP7_75t_L g560 ( .A(n_450), .B(n_185), .C(n_54), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_503), .B(n_429), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_458), .B(n_415), .Y(n_562) );
BUFx3_ASAP7_75t_L g563 ( .A(n_484), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_462), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_463), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_461), .Y(n_566) );
BUFx2_ASAP7_75t_L g567 ( .A(n_455), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_552), .B(n_402), .C(n_415), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_465), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_466), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_471), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_461), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_456), .B(n_445), .Y(n_573) );
INVx6_ASAP7_75t_L g574 ( .A(n_517), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_536), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_536), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_503), .B(n_429), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_504), .B(n_436), .Y(n_578) );
BUFx3_ASAP7_75t_L g579 ( .A(n_493), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_456), .B(n_445), .Y(n_580) );
NAND2x1_ASAP7_75t_L g581 ( .A(n_517), .B(n_436), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_490), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_488), .Y(n_583) );
NAND2xp33_ASAP7_75t_SL g584 ( .A(n_517), .B(n_446), .Y(n_584) );
OR2x6_ASAP7_75t_L g585 ( .A(n_526), .B(n_436), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_504), .B(n_435), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_490), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_496), .B(n_435), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_506), .B(n_410), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_464), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_506), .B(n_423), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_510), .B(n_423), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_494), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_494), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_474), .B(n_427), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_510), .B(n_423), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_464), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_498), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_512), .B(n_433), .Y(n_599) );
INVxp67_ASAP7_75t_SL g600 ( .A(n_472), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_511), .B(n_423), .Y(n_601) );
AOI321xp33_ASAP7_75t_L g602 ( .A1(n_528), .A2(n_448), .A3(n_421), .B1(n_433), .B2(n_402), .C(n_427), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_511), .B(n_400), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_513), .B(n_400), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_498), .Y(n_605) );
NOR2xp67_ASAP7_75t_L g606 ( .A(n_559), .B(n_421), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_458), .B(n_427), .Y(n_607) );
NOR2xp33_ASAP7_75t_R g608 ( .A(n_516), .B(n_448), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_478), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_478), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_480), .B(n_427), .Y(n_611) );
INVxp33_ASAP7_75t_L g612 ( .A(n_491), .Y(n_612) );
CKINVDCx16_ASAP7_75t_R g613 ( .A(n_513), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_480), .B(n_427), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_501), .B(n_400), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_501), .B(n_400), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_472), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_519), .B(n_447), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_475), .B(n_427), .Y(n_619) );
NAND4xp25_ASAP7_75t_L g620 ( .A(n_534), .B(n_447), .C(n_55), .D(n_57), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_500), .B(n_507), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_546), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_459), .B(n_447), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_459), .B(n_447), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_546), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_475), .B(n_31), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_460), .B(n_63), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_485), .B(n_66), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_530), .B(n_67), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_512), .A2(n_242), .B1(n_214), .B2(n_73), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_460), .B(n_68), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_476), .B(n_69), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_531), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_491), .B(n_74), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_487), .Y(n_635) );
AND2x4_ASAP7_75t_L g636 ( .A(n_530), .B(n_79), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_531), .B(n_81), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_558), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_481), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_533), .B(n_84), .Y(n_640) );
AOI211xp5_ASAP7_75t_L g641 ( .A1(n_552), .A2(n_86), .B(n_88), .C(n_90), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_493), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_533), .B(n_91), .Y(n_643) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_481), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_482), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_543), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_530), .B(n_93), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_467), .B(n_94), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_486), .B(n_95), .Y(n_649) );
AND2x4_ASAP7_75t_SL g650 ( .A(n_555), .B(n_96), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_543), .Y(n_651) );
NAND3xp33_ASAP7_75t_SL g652 ( .A(n_553), .B(n_97), .C(n_101), .Y(n_652) );
AOI321xp33_ASAP7_75t_L g653 ( .A1(n_528), .A2(n_103), .A3(n_104), .B1(n_106), .B2(n_108), .C(n_110), .Y(n_653) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_495), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_505), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_537), .A2(n_214), .B1(n_242), .B2(n_112), .Y(n_656) );
NAND2xp33_ASAP7_75t_R g657 ( .A(n_495), .B(n_113), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_508), .B(n_242), .Y(n_658) );
NOR2xp33_ASAP7_75t_SL g659 ( .A(n_548), .B(n_242), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_489), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_489), .B(n_470), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_489), .B(n_470), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_505), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_468), .A2(n_541), .B1(n_514), .B2(n_473), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_482), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_509), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_467), .B(n_509), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_473), .B(n_554), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_556), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_473), .B(n_555), .Y(n_670) );
INVxp67_ASAP7_75t_SL g671 ( .A(n_497), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_556), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_520), .Y(n_673) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_497), .Y(n_674) );
NOR3xp33_ASAP7_75t_SL g675 ( .A(n_549), .B(n_477), .C(n_557), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_520), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_555), .B(n_483), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_667), .B(n_486), .Y(n_678) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_588), .B(n_514), .C(n_550), .D(n_551), .Y(n_679) );
OAI21xp33_ASAP7_75t_L g680 ( .A1(n_618), .A2(n_550), .B(n_539), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_564), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_661), .B(n_486), .Y(n_682) );
INVxp67_ASAP7_75t_L g683 ( .A(n_638), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_565), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_635), .B(n_524), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g686 ( .A(n_618), .B(n_545), .C(n_544), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_665), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_613), .B(n_524), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_571), .Y(n_689) );
AND3x1_ASAP7_75t_L g690 ( .A(n_561), .B(n_560), .C(n_457), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_569), .Y(n_691) );
NOR2x1_ASAP7_75t_L g692 ( .A(n_567), .B(n_540), .Y(n_692) );
INVx1_ASAP7_75t_SL g693 ( .A(n_583), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_588), .B(n_522), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_662), .B(n_483), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g696 ( .A1(n_620), .A2(n_525), .B(n_518), .C(n_529), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_585), .B(n_544), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_668), .B(n_483), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_655), .B(n_547), .Y(n_699) );
AOI222xp33_ASAP7_75t_L g700 ( .A1(n_599), .A2(n_539), .B1(n_538), .B2(n_521), .C1(n_515), .C2(n_547), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_670), .B(n_523), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_663), .B(n_538), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_621), .B(n_523), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_666), .B(n_502), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_570), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_665), .Y(n_706) );
OAI31xp33_ASAP7_75t_L g707 ( .A1(n_584), .A2(n_516), .A3(n_542), .B(n_502), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_582), .Y(n_708) );
BUFx2_ASAP7_75t_SL g709 ( .A(n_577), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_642), .B(n_654), .Y(n_710) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_674), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_587), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_593), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_578), .B(n_535), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_594), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_575), .B(n_535), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_677), .B(n_532), .Y(n_717) );
INVxp67_ASAP7_75t_L g718 ( .A(n_638), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_674), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_576), .B(n_532), .Y(n_720) );
INVx1_ASAP7_75t_SL g721 ( .A(n_574), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_603), .B(n_492), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_598), .Y(n_723) );
NOR2xp33_ASAP7_75t_SL g724 ( .A(n_650), .B(n_542), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_622), .B(n_469), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_625), .B(n_469), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_585), .B(n_492), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_586), .B(n_492), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_563), .B(n_492), .Y(n_729) );
INVxp67_ASAP7_75t_L g730 ( .A(n_609), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_563), .B(n_492), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_589), .B(n_469), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_605), .Y(n_733) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_609), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_633), .B(n_479), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_646), .B(n_542), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_651), .B(n_479), .Y(n_737) );
INVxp67_ASAP7_75t_L g738 ( .A(n_610), .Y(n_738) );
NAND2x1_ASAP7_75t_L g739 ( .A(n_574), .B(n_540), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_660), .B(n_527), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_642), .B(n_527), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_579), .B(n_499), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_669), .Y(n_743) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_600), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_672), .B(n_623), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_624), .B(n_573), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_566), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_599), .B(n_612), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_585), .B(n_581), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_579), .B(n_612), .Y(n_750) );
INVx2_ASAP7_75t_SL g751 ( .A(n_574), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_608), .B(n_606), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_673), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_654), .B(n_592), .Y(n_754) );
INVx1_ASAP7_75t_SL g755 ( .A(n_650), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_676), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_562), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_580), .B(n_596), .Y(n_758) );
OR2x2_ASAP7_75t_L g759 ( .A(n_611), .B(n_614), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_600), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g761 ( .A1(n_680), .A2(n_679), .B1(n_694), .B2(n_748), .C(n_746), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_711), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_754), .B(n_601), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_739), .A2(n_584), .B(n_652), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_694), .A2(n_657), .B1(n_664), .B2(n_591), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_748), .A2(n_664), .B1(n_616), .B2(n_615), .C(n_652), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_728), .A2(n_608), .B1(n_568), .B2(n_604), .Y(n_767) );
OAI211xp5_ASAP7_75t_L g768 ( .A1(n_696), .A2(n_653), .B(n_641), .C(n_630), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_755), .A2(n_752), .B1(n_688), .B2(n_709), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g770 ( .A1(n_690), .A2(n_602), .B1(n_657), .B2(n_675), .C(n_630), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_711), .Y(n_771) );
A2O1A1Ixp33_ASAP7_75t_L g772 ( .A1(n_707), .A2(n_675), .B(n_636), .C(n_629), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_682), .B(n_610), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_752), .A2(n_640), .B1(n_637), .B2(n_643), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_691), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_736), .A2(n_628), .B1(n_595), .B2(n_648), .Y(n_776) );
NAND3xp33_ASAP7_75t_L g777 ( .A(n_683), .B(n_619), .C(n_632), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_732), .B(n_607), .Y(n_778) );
AOI32xp33_ASAP7_75t_L g779 ( .A1(n_724), .A2(n_636), .A3(n_647), .B1(n_629), .B2(n_649), .Y(n_779) );
AOI22xp33_ASAP7_75t_SL g780 ( .A1(n_749), .A2(n_631), .B1(n_627), .B2(n_647), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_705), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_681), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g783 ( .A1(n_683), .A2(n_649), .B(n_626), .Y(n_783) );
O2A1O1Ixp33_ASAP7_75t_L g784 ( .A1(n_718), .A2(n_634), .B(n_649), .C(n_659), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_736), .A2(n_658), .B1(n_671), .B2(n_644), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_684), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_689), .B(n_658), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g788 ( .A(n_749), .B(n_566), .Y(n_788) );
OR2x2_ASAP7_75t_L g789 ( .A(n_759), .B(n_671), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_749), .A2(n_644), .B1(n_590), .B2(n_597), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_695), .B(n_572), .Y(n_791) );
INVxp67_ASAP7_75t_L g792 ( .A(n_710), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_687), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_718), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_742), .A2(n_572), .B1(n_590), .B2(n_597), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_745), .B(n_617), .Y(n_796) );
OAI21xp33_ASAP7_75t_SL g797 ( .A1(n_751), .A2(n_617), .B(n_639), .Y(n_797) );
NOR2x1_ASAP7_75t_L g798 ( .A(n_693), .B(n_639), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_751), .A2(n_645), .B1(n_656), .B2(n_721), .Y(n_799) );
OAI21xp5_ASAP7_75t_SL g800 ( .A1(n_727), .A2(n_645), .B(n_700), .Y(n_800) );
OR2x2_ASAP7_75t_L g801 ( .A(n_758), .B(n_703), .Y(n_801) );
OAI211xp5_ASAP7_75t_SL g802 ( .A1(n_730), .A2(n_738), .B(n_692), .C(n_686), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_701), .B(n_717), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_708), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_712), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_750), .B(n_698), .Y(n_806) );
OAI322xp33_ASAP7_75t_L g807 ( .A1(n_730), .A2(n_738), .A3(n_678), .B1(n_757), .B2(n_702), .C1(n_726), .C2(n_725), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_801), .B(n_685), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_761), .B(n_734), .Y(n_809) );
OAI311xp33_ASAP7_75t_L g810 ( .A1(n_766), .A2(n_741), .A3(n_735), .B1(n_737), .C1(n_729), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_763), .B(n_722), .Y(n_811) );
OAI22xp5_ASAP7_75t_SL g812 ( .A1(n_780), .A2(n_744), .B1(n_727), .B2(n_734), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_770), .A2(n_727), .B1(n_722), .B2(n_697), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_762), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_803), .B(n_714), .Y(n_815) );
INVxp67_ASAP7_75t_L g816 ( .A(n_798), .Y(n_816) );
INVxp67_ASAP7_75t_L g817 ( .A(n_794), .Y(n_817) );
OAI211xp5_ASAP7_75t_L g818 ( .A1(n_800), .A2(n_744), .B(n_699), .C(n_704), .Y(n_818) );
INVxp67_ASAP7_75t_SL g819 ( .A(n_789), .Y(n_819) );
INVxp67_ASAP7_75t_SL g820 ( .A(n_771), .Y(n_820) );
NAND3xp33_ASAP7_75t_L g821 ( .A(n_761), .B(n_760), .C(n_720), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_792), .B(n_715), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_795), .B(n_733), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_780), .A2(n_697), .B1(n_731), .B2(n_756), .Y(n_824) );
INVxp67_ASAP7_75t_L g825 ( .A(n_769), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_793), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_775), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_781), .Y(n_828) );
HAxp5_ASAP7_75t_SL g829 ( .A(n_765), .B(n_723), .CON(n_829), .SN(n_829) );
OAI21xp5_ASAP7_75t_L g830 ( .A1(n_772), .A2(n_716), .B(n_697), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_782), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_778), .B(n_743), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_808), .Y(n_833) );
NOR2x1_ASAP7_75t_L g834 ( .A(n_818), .B(n_802), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_809), .B(n_766), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_828), .Y(n_836) );
AOI211xp5_ASAP7_75t_SL g837 ( .A1(n_812), .A2(n_768), .B(n_764), .C(n_802), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_828), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_825), .A2(n_768), .B1(n_767), .B2(n_797), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_808), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_821), .B(n_786), .Y(n_841) );
AO22x1_ASAP7_75t_L g842 ( .A1(n_824), .A2(n_783), .B1(n_779), .B2(n_787), .Y(n_842) );
OA22x2_ASAP7_75t_L g843 ( .A1(n_829), .A2(n_774), .B1(n_785), .B2(n_788), .Y(n_843) );
OAI21xp5_ASAP7_75t_SL g844 ( .A1(n_829), .A2(n_784), .B(n_764), .Y(n_844) );
A2O1A1Ixp33_ASAP7_75t_SL g845 ( .A1(n_813), .A2(n_830), .B(n_816), .C(n_817), .Y(n_845) );
AOI211xp5_ASAP7_75t_SL g846 ( .A1(n_844), .A2(n_810), .B(n_799), .C(n_807), .Y(n_846) );
NOR2x1_ASAP7_75t_L g847 ( .A(n_844), .B(n_784), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_843), .A2(n_822), .B1(n_819), .B2(n_823), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_835), .A2(n_777), .B1(n_832), .B2(n_776), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_839), .A2(n_831), .B1(n_827), .B2(n_790), .Y(n_850) );
A2O1A1Ixp33_ASAP7_75t_L g851 ( .A1(n_837), .A2(n_811), .B(n_815), .C(n_773), .Y(n_851) );
NOR3xp33_ASAP7_75t_L g852 ( .A(n_834), .B(n_820), .C(n_814), .Y(n_852) );
NAND3xp33_ASAP7_75t_SL g853 ( .A(n_848), .B(n_837), .C(n_845), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_849), .B(n_841), .Y(n_854) );
NOR2x1_ASAP7_75t_L g855 ( .A(n_847), .B(n_833), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_850), .Y(n_856) );
OR4x2_ASAP7_75t_L g857 ( .A(n_853), .B(n_851), .C(n_842), .D(n_846), .Y(n_857) );
OR4x2_ASAP7_75t_L g858 ( .A(n_855), .B(n_852), .C(n_840), .D(n_811), .Y(n_858) );
OR3x1_ASAP7_75t_L g859 ( .A(n_856), .B(n_838), .C(n_836), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_857), .Y(n_860) );
AOI21xp5_ASAP7_75t_L g861 ( .A1(n_857), .A2(n_854), .B(n_814), .Y(n_861) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_861), .Y(n_862) );
OAI22xp5_ASAP7_75t_SL g863 ( .A1(n_860), .A2(n_859), .B1(n_858), .B2(n_805), .Y(n_863) );
A2O1A1Ixp33_ASAP7_75t_L g864 ( .A1(n_862), .A2(n_804), .B(n_815), .C(n_826), .Y(n_864) );
OAI221xp5_ASAP7_75t_L g865 ( .A1(n_863), .A2(n_826), .B1(n_796), .B2(n_713), .C(n_753), .Y(n_865) );
AOI222xp33_ASAP7_75t_SL g866 ( .A1(n_865), .A2(n_687), .B1(n_706), .B2(n_719), .C1(n_747), .C2(n_806), .Y(n_866) );
AND2x2_ASAP7_75t_SL g867 ( .A(n_866), .B(n_864), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_867), .A2(n_791), .B1(n_740), .B2(n_719), .Y(n_868) );
endmodule