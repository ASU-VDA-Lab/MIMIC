module fake_ariane_88_n_862 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_862);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_862;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_779;
wire n_731;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_782;
wire n_650;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_767;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

BUFx10_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_100),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_49),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_44),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_27),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_2),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_69),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_25),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_97),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_6),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_102),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_140),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_21),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_47),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_9),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_167),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_5),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_61),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_48),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_20),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_152),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_147),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_118),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_95),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_111),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_67),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_116),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_60),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_117),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_127),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_87),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_18),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_72),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_16),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_115),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_38),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_84),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_82),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_81),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_68),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_121),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_L g226 ( 
.A(n_35),
.B(n_124),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_79),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_64),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_4),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_76),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_107),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_158),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_94),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_14),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_88),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_141),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_9),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_130),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_106),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_136),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_137),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_120),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_57),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_0),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_138),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_86),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_45),
.B(n_108),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_22),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_20),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

BUFx8_ASAP7_75t_SL g251 ( 
.A(n_244),
.Y(n_251)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_178),
.A2(n_0),
.B(n_1),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_249),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_189),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_191),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_1),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_213),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_205),
.Y(n_263)
);

CKINVDCx6p67_ASAP7_75t_R g264 ( 
.A(n_193),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_233),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_176),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_205),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_224),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_176),
.B(n_2),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_224),
.A2(n_78),
.B(n_173),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_211),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_183),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_184),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

OAI21x1_ASAP7_75t_L g279 ( 
.A1(n_248),
.A2(n_77),
.B(n_172),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_185),
.B(n_3),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_192),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_194),
.Y(n_282)
);

OAI22x1_ASAP7_75t_SL g283 ( 
.A1(n_200),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_188),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_239),
.B(n_23),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_195),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_204),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_177),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_206),
.Y(n_291)
);

CKINVDCx11_ASAP7_75t_R g292 ( 
.A(n_180),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_210),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_220),
.A2(n_240),
.B(n_222),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_241),
.B(n_6),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_243),
.A2(n_7),
.B(n_8),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_179),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_226),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_181),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_197),
.B(n_7),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_260),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

INVx11_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_285),
.A2(n_216),
.B1(n_229),
.B2(n_234),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_253),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_254),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_254),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_260),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_209),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_266),
.B(n_232),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g320 ( 
.A(n_256),
.B(n_258),
.C(n_290),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_270),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_278),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_257),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_182),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_267),
.B(n_186),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_267),
.B(n_187),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_267),
.B(n_190),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_267),
.B(n_196),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_257),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_257),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_257),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_274),
.B(n_198),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_274),
.B(n_199),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_288),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_257),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_257),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_288),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_259),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_266),
.B(n_201),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_290),
.A2(n_247),
.B1(n_245),
.B2(n_242),
.Y(n_346)
);

AO21x2_ASAP7_75t_L g347 ( 
.A1(n_295),
.A2(n_238),
.B(n_236),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_259),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_274),
.B(n_202),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_281),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_281),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_274),
.B(n_203),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_350),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_305),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_314),
.B(n_298),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_350),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_350),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_306),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_347),
.A2(n_296),
.B1(n_252),
.B2(n_297),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_298),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_315),
.B(n_264),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_303),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_312),
.A2(n_295),
.B(n_280),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_306),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_302),
.B(n_269),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_307),
.B(n_271),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_308),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_269),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_315),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_269),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_312),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_339),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_312),
.B(n_269),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_339),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_307),
.B(n_271),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_302),
.B(n_276),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_308),
.B(n_296),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_296),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_318),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_313),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_318),
.B(n_296),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_331),
.B(n_276),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_319),
.B(n_276),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_319),
.B(n_293),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_346),
.A2(n_301),
.B1(n_264),
.B2(n_283),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_320),
.A2(n_344),
.B1(n_337),
.B2(n_349),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_316),
.A2(n_283),
.B1(n_273),
.B2(n_293),
.Y(n_392)
);

NAND3xp33_ASAP7_75t_SL g393 ( 
.A(n_332),
.B(n_275),
.C(n_255),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_347),
.A2(n_252),
.B1(n_297),
.B2(n_294),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_304),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_319),
.B(n_263),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_333),
.A2(n_252),
.B1(n_297),
.B2(n_284),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_352),
.B(n_263),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_313),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_321),
.B(n_277),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_310),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_342),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_327),
.B(n_263),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_327),
.B(n_263),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_321),
.B(n_292),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_311),
.B(n_263),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_311),
.B(n_263),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_317),
.B(n_281),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_322),
.B(n_323),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_322),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_317),
.B(n_281),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

A2O1A1Ixp33_ASAP7_75t_L g415 ( 
.A1(n_342),
.A2(n_272),
.B(n_279),
.C(n_294),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_325),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_355),
.B(n_324),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_383),
.B(n_325),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_375),
.B(n_326),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_372),
.B(n_345),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_368),
.A2(n_347),
.B1(n_277),
.B2(n_282),
.Y(n_423)
);

A2O1A1Ixp33_ASAP7_75t_L g424 ( 
.A1(n_411),
.A2(n_272),
.B(n_279),
.C(n_326),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_378),
.B(n_304),
.Y(n_425)
);

O2A1O1Ixp33_ASAP7_75t_L g426 ( 
.A1(n_375),
.A2(n_284),
.B(n_286),
.C(n_287),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_374),
.A2(n_351),
.B(n_334),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_390),
.A2(n_282),
.B1(n_291),
.B2(n_212),
.Y(n_428)
);

OR2x6_ASAP7_75t_L g429 ( 
.A(n_363),
.B(n_291),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_386),
.B(n_299),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_354),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_397),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_386),
.B(n_299),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_371),
.A2(n_252),
.B1(n_297),
.B2(n_286),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_400),
.A2(n_376),
.B(n_373),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_381),
.A2(n_351),
.B(n_348),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_251),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_377),
.B(n_286),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_407),
.B(n_281),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_356),
.Y(n_440)
);

BUFx12f_ASAP7_75t_L g441 ( 
.A(n_358),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_360),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_366),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_404),
.Y(n_444)
);

NOR2x1_ASAP7_75t_L g445 ( 
.A(n_393),
.B(n_286),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_392),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_385),
.A2(n_348),
.B(n_343),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_416),
.A2(n_281),
.B1(n_287),
.B2(n_289),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_377),
.B(n_379),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_387),
.A2(n_343),
.B(n_341),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_353),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_367),
.A2(n_341),
.B(n_340),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_379),
.B(n_287),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_367),
.A2(n_340),
.B(n_335),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_362),
.B(n_411),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_380),
.A2(n_370),
.B1(n_384),
.B2(n_401),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_389),
.B(n_207),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_398),
.A2(n_335),
.B(n_334),
.Y(n_460)
);

NAND3xp33_ASAP7_75t_L g461 ( 
.A(n_362),
.B(n_230),
.C(n_214),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_380),
.A2(n_328),
.B(n_336),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_365),
.A2(n_388),
.B(n_382),
.Y(n_463)
);

OAI21x1_ASAP7_75t_L g464 ( 
.A1(n_399),
.A2(n_328),
.B(n_289),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_412),
.A2(n_336),
.B(n_228),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_414),
.A2(n_336),
.B(n_231),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_418),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_357),
.A2(n_359),
.B(n_405),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_417),
.B(n_287),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_406),
.A2(n_336),
.B(n_227),
.Y(n_470)
);

AOI21x1_ASAP7_75t_L g471 ( 
.A1(n_410),
.A2(n_336),
.B(n_259),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_358),
.Y(n_472)
);

A2O1A1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_361),
.A2(n_289),
.B(n_225),
.C(n_235),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_415),
.A2(n_289),
.B(n_223),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_361),
.A2(n_221),
.B(n_219),
.C(n_208),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_358),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_417),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_364),
.B(n_259),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_402),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_369),
.B(n_259),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_395),
.B(n_259),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_395),
.B(n_261),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_408),
.A2(n_261),
.B(n_85),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_391),
.B(n_261),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_409),
.A2(n_261),
.B(n_89),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_395),
.B(n_8),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_410),
.A2(n_261),
.B(n_90),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_395),
.B(n_261),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_403),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_457),
.B(n_403),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_429),
.B(n_403),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_450),
.A2(n_403),
.B(n_413),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_463),
.A2(n_394),
.B(n_413),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_430),
.B(n_394),
.Y(n_494)
);

AO31x2_ASAP7_75t_L g495 ( 
.A1(n_473),
.A2(n_10),
.A3(n_11),
.B(n_12),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_433),
.B(n_10),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_429),
.B(n_11),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_446),
.B(n_12),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_464),
.A2(n_92),
.B(n_171),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_435),
.A2(n_83),
.B(n_170),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_432),
.B(n_24),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_471),
.A2(n_93),
.B(n_169),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_429),
.Y(n_503)
);

AND3x4_ASAP7_75t_L g504 ( 
.A(n_445),
.B(n_13),
.C(n_14),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_467),
.B(n_13),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_474),
.A2(n_96),
.B(n_168),
.Y(n_506)
);

A2O1A1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_428),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_427),
.A2(n_80),
.B(n_166),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_431),
.B(n_15),
.Y(n_509)
);

AOI21x1_ASAP7_75t_SL g510 ( 
.A1(n_438),
.A2(n_17),
.B(n_18),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_451),
.A2(n_99),
.B(n_26),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_432),
.B(n_28),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_468),
.A2(n_101),
.B(n_29),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_447),
.A2(n_103),
.B(n_30),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_440),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_442),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_460),
.A2(n_104),
.B(n_31),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_454),
.A2(n_105),
.B(n_32),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_444),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_477),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_436),
.A2(n_455),
.B(n_453),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_458),
.A2(n_110),
.B(n_33),
.Y(n_522)
);

AO31x2_ASAP7_75t_L g523 ( 
.A1(n_424),
.A2(n_19),
.A3(n_34),
.B(n_36),
.Y(n_523)
);

INVx3_ASAP7_75t_SL g524 ( 
.A(n_459),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_443),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_479),
.A2(n_19),
.B1(n_37),
.B2(n_39),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_469),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_448),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_421),
.A2(n_43),
.B(n_46),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_439),
.Y(n_530)
);

INVx6_ASAP7_75t_L g531 ( 
.A(n_441),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_419),
.B(n_50),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_462),
.A2(n_51),
.B(n_52),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_434),
.A2(n_53),
.B(n_54),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_448),
.A2(n_55),
.B(n_56),
.Y(n_535)
);

NAND2x1p5_ASAP7_75t_L g536 ( 
.A(n_476),
.B(n_58),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_422),
.A2(n_59),
.B(n_62),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_475),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_488),
.A2(n_70),
.B(n_71),
.Y(n_539)
);

A2O1A1Ixp33_ASAP7_75t_L g540 ( 
.A1(n_426),
.A2(n_73),
.B(n_74),
.C(n_75),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_425),
.B(n_98),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_465),
.A2(n_112),
.B(n_113),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_452),
.Y(n_543)
);

OAI21x1_ASAP7_75t_L g544 ( 
.A1(n_466),
.A2(n_119),
.B(n_125),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_420),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_423),
.B(n_126),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_456),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_437),
.B(n_128),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_472),
.A2(n_129),
.B(n_131),
.Y(n_549)
);

BUFx2_ASAP7_75t_SL g550 ( 
.A(n_519),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_547),
.Y(n_551)
);

OA21x2_ASAP7_75t_L g552 ( 
.A1(n_506),
.A2(n_483),
.B(n_485),
.Y(n_552)
);

CKINVDCx11_ASAP7_75t_R g553 ( 
.A(n_548),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_491),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_499),
.A2(n_487),
.B(n_470),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_545),
.B(n_449),
.Y(n_556)
);

OA21x2_ASAP7_75t_L g557 ( 
.A1(n_534),
.A2(n_521),
.B(n_493),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_546),
.A2(n_484),
.B(n_478),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_515),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_524),
.B(n_461),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_527),
.B(n_489),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_515),
.A2(n_496),
.B1(n_516),
.B2(n_525),
.Y(n_562)
);

AOI21x1_ASAP7_75t_L g563 ( 
.A1(n_492),
.A2(n_480),
.B(n_482),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_547),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_490),
.A2(n_489),
.B(n_476),
.Y(n_565)
);

AO21x2_ASAP7_75t_L g566 ( 
.A1(n_494),
.A2(n_481),
.B(n_486),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_520),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_509),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_541),
.A2(n_489),
.B1(n_476),
.B2(n_134),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_527),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_531),
.Y(n_571)
);

OAI21x1_ASAP7_75t_SL g572 ( 
.A1(n_522),
.A2(n_132),
.B(n_133),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_543),
.B(n_135),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_511),
.A2(n_139),
.B(n_143),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_491),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_541),
.A2(n_144),
.B1(n_146),
.B2(n_148),
.Y(n_576)
);

OAI21x1_ASAP7_75t_L g577 ( 
.A1(n_513),
.A2(n_149),
.B(n_153),
.Y(n_577)
);

AO22x2_ASAP7_75t_L g578 ( 
.A1(n_504),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_578)
);

OAI22xp33_ASAP7_75t_L g579 ( 
.A1(n_548),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_498),
.B(n_174),
.Y(n_580)
);

AOI22x1_ASAP7_75t_L g581 ( 
.A1(n_500),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_581)
);

AO21x2_ASAP7_75t_L g582 ( 
.A1(n_532),
.A2(n_165),
.B(n_538),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_497),
.B(n_503),
.Y(n_583)
);

OA21x2_ASAP7_75t_L g584 ( 
.A1(n_514),
.A2(n_517),
.B(n_502),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_505),
.Y(n_585)
);

OA21x2_ASAP7_75t_L g586 ( 
.A1(n_542),
.A2(n_544),
.B(n_539),
.Y(n_586)
);

OAI22xp33_ASAP7_75t_L g587 ( 
.A1(n_497),
.A2(n_531),
.B1(n_530),
.B2(n_501),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_510),
.A2(n_533),
.B(n_508),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_518),
.A2(n_529),
.B(n_535),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_523),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_523),
.B(n_536),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_523),
.Y(n_592)
);

NAND2x1_ASAP7_75t_L g593 ( 
.A(n_512),
.B(n_537),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_540),
.A2(n_507),
.B(n_528),
.Y(n_594)
);

INVx3_ASAP7_75t_SL g595 ( 
.A(n_495),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_549),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_526),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_559),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_571),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_578),
.B(n_570),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_567),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_568),
.B(n_495),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_570),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_554),
.B(n_495),
.Y(n_604)
);

AO21x1_ASAP7_75t_SL g605 ( 
.A1(n_594),
.A2(n_569),
.B(n_585),
.Y(n_605)
);

NAND2x1p5_ASAP7_75t_L g606 ( 
.A(n_554),
.B(n_575),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_551),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_550),
.B(n_583),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_551),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_564),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_564),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_553),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_588),
.A2(n_589),
.B(n_555),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_560),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_562),
.A2(n_561),
.B(n_565),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_556),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_561),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_575),
.Y(n_618)
);

OR2x6_ASAP7_75t_L g619 ( 
.A(n_575),
.B(n_578),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_578),
.B(n_575),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_573),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_573),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_563),
.Y(n_623)
);

O2A1O1Ixp33_ASAP7_75t_SL g624 ( 
.A1(n_579),
.A2(n_593),
.B(n_576),
.C(n_587),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_587),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_590),
.Y(n_626)
);

BUFx2_ASAP7_75t_SL g627 ( 
.A(n_571),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_590),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_588),
.A2(n_589),
.B(n_555),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_580),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_592),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_560),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_592),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_579),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_591),
.Y(n_635)
);

NAND2x1p5_ASAP7_75t_L g636 ( 
.A(n_597),
.B(n_596),
.Y(n_636)
);

O2A1O1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_572),
.A2(n_582),
.B(n_557),
.C(n_595),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_595),
.B(n_581),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_566),
.B(n_557),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_557),
.B(n_558),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_577),
.B(n_553),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_635),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_635),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_604),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_600),
.B(n_591),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_603),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_600),
.B(n_591),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_619),
.B(n_577),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_616),
.B(n_591),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_619),
.B(n_558),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_618),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_601),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_SL g653 ( 
.A1(n_619),
.A2(n_591),
.B1(n_582),
.B2(n_574),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_602),
.B(n_574),
.Y(n_654)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_636),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_602),
.B(n_619),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_603),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_626),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_620),
.B(n_574),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_620),
.B(n_586),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_621),
.B(n_584),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_604),
.B(n_586),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_626),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_628),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_604),
.B(n_586),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_628),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_635),
.B(n_584),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_598),
.B(n_584),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_617),
.B(n_552),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_631),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_608),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_634),
.B(n_552),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_599),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_641),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_610),
.B(n_552),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_632),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_610),
.B(n_611),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_636),
.B(n_639),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_611),
.B(n_607),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_609),
.B(n_622),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_639),
.B(n_632),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_605),
.B(n_630),
.Y(n_682)
);

INVx5_ASAP7_75t_L g683 ( 
.A(n_641),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_631),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_625),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_614),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_633),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_599),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_640),
.B(n_633),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_615),
.B(n_641),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_612),
.B(n_627),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_623),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_662),
.B(n_640),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_662),
.B(n_641),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_671),
.B(n_606),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_665),
.B(n_623),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_652),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_642),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_665),
.B(n_613),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_644),
.B(n_613),
.Y(n_700)
);

NOR2xp67_ASAP7_75t_L g701 ( 
.A(n_676),
.B(n_638),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_680),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_667),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_644),
.B(n_629),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_680),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_686),
.B(n_606),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_688),
.B(n_685),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_660),
.B(n_629),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_679),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_682),
.B(n_624),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_683),
.B(n_638),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_679),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_681),
.B(n_624),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_658),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_658),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_668),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_666),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_666),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_677),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_677),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_683),
.B(n_637),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_682),
.B(n_681),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_660),
.B(n_678),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_668),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_669),
.B(n_690),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_678),
.B(n_672),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_670),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_669),
.B(n_651),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_683),
.B(n_674),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_646),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_646),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_657),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_663),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_693),
.B(n_690),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_707),
.B(n_651),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_693),
.B(n_659),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_697),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_725),
.B(n_659),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_723),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_702),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_705),
.Y(n_741)
);

AND2x4_ASAP7_75t_SL g742 ( 
.A(n_698),
.B(n_711),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_710),
.B(n_706),
.Y(n_743)
);

NAND2x1p5_ASAP7_75t_L g744 ( 
.A(n_701),
.B(n_683),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_733),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_733),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_709),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_712),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_725),
.B(n_654),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_703),
.B(n_683),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_719),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_728),
.B(n_654),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_720),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_724),
.B(n_656),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_703),
.B(n_674),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_723),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_699),
.B(n_656),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_726),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_694),
.B(n_674),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_714),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_713),
.B(n_698),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_699),
.B(n_672),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_726),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_722),
.B(n_661),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_698),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_694),
.B(n_667),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_716),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_757),
.B(n_716),
.Y(n_768)
);

OAI322xp33_ASAP7_75t_L g769 ( 
.A1(n_764),
.A2(n_743),
.A3(n_756),
.B1(n_737),
.B2(n_763),
.C1(n_758),
.C2(n_741),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_739),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_743),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_735),
.B(n_713),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_757),
.B(n_749),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_744),
.B(n_648),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_760),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_767),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_749),
.B(n_708),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_746),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_746),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_745),
.Y(n_780)
);

CKINVDCx16_ASAP7_75t_R g781 ( 
.A(n_754),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_752),
.B(n_708),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_736),
.B(n_696),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_751),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_736),
.B(n_696),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_755),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_738),
.B(n_762),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_753),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_762),
.B(n_700),
.Y(n_789)
);

NAND2x1_ASAP7_75t_L g790 ( 
.A(n_770),
.B(n_755),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_780),
.Y(n_791)
);

OAI322xp33_ASAP7_75t_L g792 ( 
.A1(n_771),
.A2(n_740),
.A3(n_748),
.B1(n_747),
.B2(n_761),
.C1(n_738),
.C2(n_754),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_781),
.B(n_691),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_778),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_779),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_776),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_784),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_773),
.B(n_766),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_774),
.A2(n_647),
.B1(n_645),
.B2(n_653),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_788),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_774),
.A2(n_734),
.B1(n_711),
.B2(n_750),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_769),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_793),
.B(n_769),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_802),
.A2(n_801),
.B1(n_648),
.B2(n_774),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_791),
.B(n_772),
.Y(n_805)
);

OAI322xp33_ASAP7_75t_L g806 ( 
.A1(n_797),
.A2(n_782),
.A3(n_787),
.B1(n_785),
.B2(n_789),
.C1(n_777),
.C2(n_783),
.Y(n_806)
);

OAI31xp33_ASAP7_75t_L g807 ( 
.A1(n_799),
.A2(n_734),
.A3(n_786),
.B(n_645),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_791),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_796),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_790),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_803),
.B(n_800),
.Y(n_811)
);

AOI222xp33_ASAP7_75t_L g812 ( 
.A1(n_804),
.A2(n_805),
.B1(n_809),
.B2(n_808),
.C1(n_794),
.C2(n_795),
.Y(n_812)
);

OAI21xp33_ASAP7_75t_SL g813 ( 
.A1(n_810),
.A2(n_798),
.B(n_768),
.Y(n_813)
);

AOI322xp5_ASAP7_75t_L g814 ( 
.A1(n_804),
.A2(n_792),
.A3(n_647),
.B1(n_761),
.B2(n_786),
.C1(n_766),
.C2(n_721),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_807),
.A2(n_721),
.B1(n_648),
.B2(n_649),
.Y(n_815)
);

OAI221xp5_ASAP7_75t_L g816 ( 
.A1(n_806),
.A2(n_648),
.B1(n_695),
.B2(n_775),
.C(n_744),
.Y(n_816)
);

XNOR2x1_ASAP7_75t_L g817 ( 
.A(n_804),
.B(n_711),
.Y(n_817)
);

OAI211xp5_ASAP7_75t_SL g818 ( 
.A1(n_811),
.A2(n_765),
.B(n_643),
.C(n_650),
.Y(n_818)
);

NAND4xp25_ASAP7_75t_L g819 ( 
.A(n_812),
.B(n_704),
.C(n_700),
.D(n_673),
.Y(n_819)
);

AOI211xp5_ASAP7_75t_SL g820 ( 
.A1(n_816),
.A2(n_704),
.B(n_755),
.C(n_667),
.Y(n_820)
);

NOR3xp33_ASAP7_75t_L g821 ( 
.A(n_813),
.B(n_673),
.C(n_765),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_814),
.B(n_673),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_822),
.Y(n_823)
);

AND4x1_ASAP7_75t_L g824 ( 
.A(n_820),
.B(n_815),
.C(n_817),
.D(n_742),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_818),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_823),
.B(n_821),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_825),
.B(n_819),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_825),
.Y(n_828)
);

NOR2x1_ASAP7_75t_L g829 ( 
.A(n_825),
.B(n_750),
.Y(n_829)
);

XNOR2x1_ASAP7_75t_L g830 ( 
.A(n_828),
.B(n_824),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_829),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_826),
.Y(n_832)
);

INVx3_ASAP7_75t_SL g833 ( 
.A(n_827),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_828),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_828),
.Y(n_835)
);

AO22x2_ASAP7_75t_L g836 ( 
.A1(n_832),
.A2(n_835),
.B1(n_834),
.B2(n_831),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_830),
.A2(n_655),
.B(n_742),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_832),
.B(n_833),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_831),
.Y(n_839)
);

AO22x2_ASAP7_75t_L g840 ( 
.A1(n_832),
.A2(n_759),
.B1(n_721),
.B2(n_750),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_830),
.A2(n_759),
.B1(n_642),
.B2(n_643),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_832),
.B(n_759),
.Y(n_842)
);

AO22x2_ASAP7_75t_L g843 ( 
.A1(n_832),
.A2(n_729),
.B1(n_643),
.B2(n_650),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_839),
.A2(n_698),
.B1(n_642),
.B2(n_675),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_838),
.A2(n_698),
.B(n_642),
.Y(n_845)
);

AOI32xp33_ASAP7_75t_L g846 ( 
.A1(n_836),
.A2(n_729),
.A3(n_675),
.B1(n_760),
.B2(n_730),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_841),
.A2(n_642),
.B1(n_729),
.B2(n_732),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_842),
.B(n_731),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_845),
.A2(n_837),
.B(n_840),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_846),
.A2(n_843),
.B(n_692),
.Y(n_850)
);

XNOR2x1_ASAP7_75t_SL g851 ( 
.A(n_844),
.B(n_687),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_847),
.A2(n_692),
.B(n_689),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_L g853 ( 
.A1(n_849),
.A2(n_848),
.B1(n_689),
.B2(n_657),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_852),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_850),
.A2(n_714),
.B1(n_727),
.B2(n_718),
.Y(n_855)
);

OAI21xp33_ASAP7_75t_L g856 ( 
.A1(n_851),
.A2(n_663),
.B(n_664),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_853),
.A2(n_664),
.B1(n_684),
.B2(n_687),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_854),
.Y(n_858)
);

OAI22x1_ASAP7_75t_L g859 ( 
.A1(n_855),
.A2(n_717),
.B1(n_727),
.B2(n_718),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_858),
.B(n_856),
.Y(n_860)
);

OR2x6_ASAP7_75t_L g861 ( 
.A(n_860),
.B(n_857),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_861),
.A2(n_859),
.B1(n_715),
.B2(n_717),
.Y(n_862)
);


endmodule