module fake_jpeg_28653_n_523 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_523);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_523;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_66),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_24),
.B(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_68),
.Y(n_158)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_79),
.Y(n_110)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_16),
.B(n_6),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_95),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_88),
.Y(n_154)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_101),
.Y(n_113)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_66),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_118),
.A2(n_37),
.B1(n_39),
.B2(n_49),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_79),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_124),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_25),
.B1(n_24),
.B2(n_49),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_122),
.A2(n_131),
.B(n_133),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_26),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_81),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_148),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_54),
.B(n_36),
.C(n_43),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_36),
.C(n_43),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_22),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_136),
.B(n_48),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_59),
.B(n_22),
.C(n_41),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_16),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_87),
.A2(n_51),
.B1(n_17),
.B2(n_27),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_142),
.A2(n_150),
.B1(n_50),
.B2(n_63),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_90),
.B(n_18),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_93),
.A2(n_17),
.B1(n_27),
.B2(n_50),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_96),
.B(n_41),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_18),
.Y(n_178)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_162),
.B(n_211),
.Y(n_250)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_122),
.Y(n_165)
);

BUFx4f_ASAP7_75t_SL g238 ( 
.A(n_165),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_107),
.A2(n_110),
.B1(n_102),
.B2(n_157),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_166),
.A2(n_196),
.B1(n_208),
.B2(n_158),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_105),
.A2(n_98),
.B1(n_86),
.B2(n_85),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_171),
.A2(n_209),
.B1(n_139),
.B2(n_108),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_172),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_173),
.B(n_210),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_107),
.B(n_110),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_176),
.Y(n_220)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_179),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_136),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_180),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_142),
.A2(n_84),
.B1(n_76),
.B2(n_75),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_184),
.B1(n_200),
.B2(n_108),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_28),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_185),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_150),
.A2(n_73),
.B1(n_68),
.B2(n_67),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_118),
.A2(n_37),
.B(n_50),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_165),
.B(n_189),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_118),
.B(n_35),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_191),
.Y(n_229)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_111),
.B(n_26),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_198),
.Y(n_235)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_140),
.B(n_28),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_197),
.Y(n_231)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_201),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_127),
.A2(n_62),
.B1(n_151),
.B2(n_153),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_109),
.B(n_114),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_203),
.Y(n_242)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_103),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_132),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_206),
.Y(n_239)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_144),
.B(n_48),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_105),
.A2(n_27),
.B1(n_31),
.B2(n_42),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_146),
.A2(n_27),
.B1(n_50),
.B2(n_46),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_152),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_165),
.A2(n_113),
.B1(n_132),
.B2(n_154),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_214),
.A2(n_208),
.B1(n_176),
.B2(n_166),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_215),
.A2(n_9),
.B(n_13),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_204),
.A2(n_138),
.B1(n_156),
.B2(n_145),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_232),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_139),
.C(n_158),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_169),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_162),
.B1(n_167),
.B2(n_200),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_194),
.A2(n_126),
.B1(n_123),
.B2(n_117),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_123),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_251),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_172),
.A2(n_126),
.B1(n_50),
.B2(n_48),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_245),
.A2(n_247),
.B1(n_177),
.B2(n_161),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_211),
.A2(n_48),
.B1(n_49),
.B2(n_38),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_48),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_184),
.B(n_182),
.C(n_162),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_252),
.A2(n_287),
.B(n_249),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_227),
.B(n_164),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_253),
.B(n_285),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_254),
.A2(n_273),
.B1(n_275),
.B2(n_286),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_255),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_225),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_257),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_220),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

OAI22x1_ASAP7_75t_L g260 ( 
.A1(n_215),
.A2(n_181),
.B1(n_162),
.B2(n_173),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_260),
.A2(n_283),
.B1(n_226),
.B2(n_231),
.Y(n_313)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_212),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_261),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_263),
.A2(n_279),
.B1(n_237),
.B2(n_244),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_225),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_265),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_191),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_270),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_239),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_267),
.B(n_277),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_223),
.Y(n_268)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_240),
.C(n_218),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_201),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_214),
.A2(n_251),
.B1(n_236),
.B2(n_229),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_190),
.B1(n_188),
.B2(n_175),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_228),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_228),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_250),
.A2(n_192),
.B1(n_163),
.B2(n_198),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_219),
.B(n_193),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_282),
.Y(n_292)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_234),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_221),
.B1(n_223),
.B2(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_246),
.Y(n_282)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_235),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_219),
.B(n_206),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_284),
.B(n_230),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_229),
.B(n_203),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_250),
.A2(n_187),
.B1(n_170),
.B2(n_168),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_290),
.A2(n_297),
.B1(n_312),
.B2(n_268),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_291),
.A2(n_304),
.B1(n_305),
.B2(n_272),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_238),
.B(n_242),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_294),
.A2(n_300),
.B(n_221),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_240),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_301),
.C(n_308),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_271),
.A2(n_230),
.B1(n_226),
.B2(n_248),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_260),
.A2(n_238),
.B(n_242),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_303),
.B(n_318),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_263),
.A2(n_238),
.B1(n_249),
.B2(n_222),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_252),
.A2(n_238),
.B1(n_249),
.B2(n_216),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_307),
.A2(n_309),
.B(n_313),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_259),
.C(n_257),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_262),
.A2(n_235),
.B(n_226),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_285),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_310),
.B(n_320),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_259),
.B(n_246),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_311),
.B(n_321),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_270),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_260),
.A2(n_254),
.B(n_274),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_319),
.B(n_252),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_267),
.B(n_231),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_216),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_279),
.B(n_234),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_282),
.C(n_258),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_286),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_323),
.Y(n_361)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_302),
.A2(n_252),
.B1(n_308),
.B2(n_319),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_325),
.A2(n_348),
.B1(n_351),
.B2(n_295),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_317),
.Y(n_326)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_326),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_301),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_340),
.C(n_352),
.Y(n_364)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_330),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_288),
.B(n_253),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_332),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_299),
.B(n_264),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_333),
.B(n_335),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_334),
.A2(n_309),
.B(n_307),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_314),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_289),
.Y(n_336)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_320),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_338),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_252),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_316),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_341),
.B(n_345),
.Y(n_378)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_289),
.Y(n_342)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_294),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_288),
.B(n_281),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_344),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_305),
.A2(n_291),
.B1(n_304),
.B2(n_321),
.Y(n_346)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_303),
.Y(n_347)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_347),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_302),
.A2(n_277),
.B1(n_276),
.B2(n_261),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_268),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_350),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_322),
.A2(n_255),
.B1(n_217),
.B2(n_224),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_311),
.B(n_217),
.C(n_255),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_353),
.A2(n_315),
.B(n_316),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_299),
.Y(n_354)
);

NAND2xp33_ASAP7_75t_R g384 ( 
.A(n_354),
.B(n_312),
.Y(n_384)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

OAI21xp33_ASAP7_75t_L g368 ( 
.A1(n_355),
.A2(n_356),
.B(n_318),
.Y(n_368)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_292),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_362),
.B(n_368),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g417 ( 
.A(n_365),
.B(n_377),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_329),
.C(n_349),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_374),
.C(n_375),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_370),
.A2(n_351),
.B(n_350),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_327),
.B(n_349),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_372),
.B(n_373),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_306),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_293),
.C(n_316),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_346),
.C(n_340),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_339),
.C(n_353),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_385),
.C(n_386),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_323),
.A2(n_295),
.B(n_293),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_380),
.A2(n_46),
.B1(n_42),
.B2(n_31),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_331),
.A2(n_312),
.B(n_12),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_382),
.A2(n_387),
.B(n_370),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_384),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_298),
.C(n_221),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_345),
.B(n_331),
.C(n_355),
.Y(n_386)
);

XOR2x2_ASAP7_75t_L g387 ( 
.A(n_323),
.B(n_221),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_330),
.Y(n_390)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_390),
.Y(n_437)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_328),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_392),
.B(n_393),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_383),
.B(n_356),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_396),
.A2(n_46),
.B(n_1),
.Y(n_436)
);

BUFx12_ASAP7_75t_L g397 ( 
.A(n_387),
.Y(n_397)
);

INVxp33_ASAP7_75t_L g439 ( 
.A(n_397),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_357),
.B(n_342),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_404),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_371),
.A2(n_348),
.B1(n_341),
.B2(n_336),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_399),
.A2(n_401),
.B1(n_378),
.B2(n_388),
.Y(n_430)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_403),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_371),
.A2(n_341),
.B1(n_324),
.B2(n_0),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_366),
.B(n_9),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_377),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_405),
.Y(n_438)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_360),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_406),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_408),
.A2(n_365),
.B(n_361),
.Y(n_421)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_359),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_409),
.A2(n_414),
.B1(n_416),
.B2(n_361),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_381),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_410),
.B(n_373),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_376),
.B(n_10),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_411),
.B(n_418),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_359),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_412),
.A2(n_378),
.B1(n_375),
.B2(n_372),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_413),
.A2(n_382),
.B1(n_31),
.B2(n_42),
.Y(n_432)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_381),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_10),
.Y(n_418)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_419),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_364),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_431),
.C(n_435),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_421),
.B(n_425),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_395),
.B(n_362),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_392),
.A2(n_388),
.B1(n_380),
.B2(n_386),
.Y(n_427)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_402),
.B(n_374),
.C(n_364),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_432),
.A2(n_391),
.B1(n_400),
.B2(n_409),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_416),
.B(n_367),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_433),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_434),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_48),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_436),
.B(n_396),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_399),
.A2(n_5),
.B1(n_13),
.B2(n_2),
.Y(n_441)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_415),
.B(n_38),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_442),
.B(n_394),
.C(n_390),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_446),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_429),
.Y(n_447)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_428),
.A2(n_407),
.B1(n_401),
.B2(n_398),
.Y(n_449)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_449),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_451),
.A2(n_460),
.B1(n_430),
.B2(n_421),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_437),
.A2(n_410),
.B1(n_405),
.B2(n_412),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_458),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_394),
.C(n_395),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_456),
.B(n_425),
.C(n_420),
.Y(n_463)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_423),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_459),
.B(n_440),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_438),
.A2(n_432),
.B1(n_434),
.B2(n_439),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_462),
.B(n_465),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_463),
.B(n_450),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_444),
.B(n_435),
.C(n_419),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_464),
.A2(n_474),
.B(n_448),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_443),
.B(n_426),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_457),
.A2(n_439),
.B(n_397),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_467),
.B(n_3),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_471),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_454),
.A2(n_408),
.B1(n_436),
.B2(n_397),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_470),
.A2(n_473),
.B1(n_475),
.B2(n_8),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_461),
.A2(n_406),
.B1(n_403),
.B2(n_424),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_442),
.Y(n_472)
);

XNOR2x1_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_476),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_461),
.A2(n_414),
.B1(n_441),
.B2(n_397),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_SL g474 ( 
.A(n_444),
.B(n_417),
.C(n_413),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_452),
.A2(n_417),
.B1(n_7),
.B2(n_3),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_456),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_448),
.C(n_453),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_481),
.B(n_486),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_478),
.B(n_457),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_482),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_466),
.B(n_451),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_484),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_485),
.B(n_491),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_453),
.C(n_445),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_490),
.C(n_472),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_477),
.Y(n_488)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_488),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_SL g489 ( 
.A1(n_467),
.A2(n_446),
.B1(n_417),
.B2(n_3),
.Y(n_489)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_489),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_38),
.C(n_5),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_478),
.B(n_4),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_491),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_470),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_499),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_500),
.A2(n_503),
.B(n_483),
.Y(n_506)
);

XNOR2x1_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_497),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_482),
.A2(n_468),
.B(n_462),
.Y(n_503)
);

OAI21x1_ASAP7_75t_SL g512 ( 
.A1(n_506),
.A2(n_498),
.B(n_12),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_496),
.C(n_504),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_508),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_496),
.A2(n_492),
.B(n_484),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_480),
.C(n_8),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_509),
.B(n_510),
.C(n_511),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_13),
.C(n_8),
.Y(n_510)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_512),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_12),
.C(n_0),
.Y(n_514)
);

OAI21xp33_ASAP7_75t_L g516 ( 
.A1(n_514),
.A2(n_12),
.B(n_0),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_516),
.B(n_513),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_518),
.B(n_515),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_517),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_520),
.A2(n_1),
.B(n_519),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_521),
.B(n_1),
.Y(n_522)
);

BUFx24_ASAP7_75t_SL g523 ( 
.A(n_522),
.Y(n_523)
);


endmodule