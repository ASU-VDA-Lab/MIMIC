module fake_netlist_5_2168_n_1786 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1786);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1786;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_42),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_66),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_146),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_111),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_95),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_122),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_4),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_22),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_61),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_39),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_54),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_10),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_14),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_137),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_67),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_68),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_49),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_82),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_62),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_76),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_80),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_169),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_34),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_57),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_84),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_33),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_79),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_53),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_132),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_52),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_98),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_157),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_161),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_13),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_9),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_63),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_110),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_168),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_2),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_60),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_87),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_21),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_20),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_112),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_134),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_143),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_59),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_21),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_151),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_118),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_23),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_14),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_154),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_59),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_36),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_10),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_119),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_116),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_16),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_23),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_43),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_165),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_45),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_71),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_1),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_96),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_64),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_107),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_35),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_24),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_162),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_24),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_38),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_106),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_141),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_55),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_58),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_50),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_160),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_48),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_155),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_1),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_130),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_4),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_75),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_129),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_17),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_52),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_42),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_17),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_124),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_51),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_101),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_50),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_97),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_6),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_105),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_26),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_103),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_35),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_30),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_51),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_77),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_90),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_86),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_99),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_150),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_94),
.Y(n_289)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_15),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_89),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_123),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_11),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_18),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_73),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_91),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_65),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_22),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_159),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_11),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_46),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_40),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_16),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_126),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_38),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_13),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_88),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_47),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_142),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_102),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_0),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_83),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_26),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_34),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_53),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_57),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_158),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_33),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_153),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_6),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_19),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_136),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_27),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_49),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_12),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_147),
.Y(n_326)
);

BUFx10_ASAP7_75t_L g327 ( 
.A(n_3),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_15),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_72),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_167),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_56),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_44),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_133),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_108),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_0),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_55),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_12),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_30),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_144),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_100),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_81),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_19),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_121),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_70),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_56),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_47),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_58),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_74),
.Y(n_348)
);

BUFx2_ASAP7_75t_SL g349 ( 
.A(n_243),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_311),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_245),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_311),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_215),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_227),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_216),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_311),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_262),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_221),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_311),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_315),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_311),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_185),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_332),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_222),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_247),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_332),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_199),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_329),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_316),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_271),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_201),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_265),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_225),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_201),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_229),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_271),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_238),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_239),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_231),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_230),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_345),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_237),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_248),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_239),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_238),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_328),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_298),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_249),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_173),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_255),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_298),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_184),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_200),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_223),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_190),
.Y(n_401)
);

INVxp33_ASAP7_75t_SL g402 ( 
.A(n_173),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_180),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_267),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_318),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_272),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_220),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_274),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_180),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_317),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_234),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_235),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_278),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_181),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_246),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_257),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_280),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_285),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_258),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_178),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_259),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_286),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_261),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_273),
.Y(n_424)
);

INVxp33_ASAP7_75t_SL g425 ( 
.A(n_181),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_282),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_318),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_283),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_287),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_183),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_288),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_294),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_183),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_299),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_302),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_320),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_174),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_366),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_366),
.B(n_223),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_357),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_357),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_363),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_367),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_363),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_350),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_350),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_367),
.B(n_276),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_400),
.B(n_192),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_370),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_391),
.B(n_238),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_357),
.B(n_262),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_370),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_374),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_357),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_377),
.B(n_276),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_374),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_L g459 ( 
.A(n_400),
.B(n_300),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_353),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_352),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_352),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_395),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_356),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_403),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_375),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_354),
.A2(n_263),
.B1(n_314),
.B2(n_250),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_375),
.B(n_284),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_356),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_382),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_382),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_400),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_359),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_359),
.Y(n_474)
);

NAND2x1p5_ASAP7_75t_L g475 ( 
.A(n_360),
.B(n_262),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_380),
.B(n_284),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_384),
.B(n_295),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_409),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_360),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_361),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_361),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_365),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_365),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_376),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_384),
.B(n_295),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_424),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_424),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_390),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_371),
.A2(n_279),
.B1(n_275),
.B2(n_270),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_355),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_376),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_390),
.A2(n_343),
.B(n_297),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_368),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_351),
.A2(n_206),
.B1(n_347),
.B2(n_346),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_398),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_393),
.B(n_297),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_399),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_399),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_393),
.B(n_343),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_407),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_397),
.B(n_194),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_407),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_411),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_397),
.B(n_195),
.Y(n_505)
);

CKINVDCx8_ASAP7_75t_R g506 ( 
.A(n_349),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_401),
.B(n_300),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_411),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_410),
.B(n_202),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_412),
.B(n_203),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_412),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_364),
.A2(n_212),
.B1(n_347),
.B2(n_346),
.Y(n_512)
);

INVx6_ASAP7_75t_L g513 ( 
.A(n_383),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_415),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_L g515 ( 
.A(n_415),
.B(n_262),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_444),
.Y(n_516)
);

OR2x6_ASAP7_75t_L g517 ( 
.A(n_513),
.B(n_349),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_441),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_457),
.B(n_262),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_444),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_441),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_444),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_506),
.B(n_391),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_444),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_506),
.B(n_379),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_479),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_457),
.B(n_291),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_457),
.B(n_476),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_506),
.B(n_386),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_479),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_461),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_446),
.Y(n_532)
);

INVx8_ASAP7_75t_L g533 ( 
.A(n_453),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_446),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_438),
.B(n_394),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_512),
.A2(n_396),
.B1(n_413),
.B2(n_404),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_447),
.Y(n_537)
);

AND2x6_ASAP7_75t_L g538 ( 
.A(n_476),
.B(n_291),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_447),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_476),
.B(n_406),
.Y(n_540)
);

INVxp33_ASAP7_75t_L g541 ( 
.A(n_467),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_465),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_461),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_509),
.A2(n_392),
.B1(n_362),
.B2(n_414),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_460),
.B(n_408),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_490),
.B(n_418),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_493),
.B(n_431),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_482),
.B(n_434),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_447),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_482),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_483),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_453),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_447),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_448),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_448),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_483),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_473),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_441),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_441),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_513),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_448),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_473),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g563 ( 
.A1(n_512),
.A2(n_358),
.B1(n_373),
.B2(n_303),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_448),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_438),
.B(n_291),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_462),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_462),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_462),
.Y(n_568)
);

INVxp33_ASAP7_75t_L g569 ( 
.A(n_467),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_473),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_473),
.Y(n_571)
);

NOR2x1p5_ASAP7_75t_L g572 ( 
.A(n_488),
.B(n_383),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_462),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_464),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_R g575 ( 
.A(n_513),
.B(n_381),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_473),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_L g577 ( 
.A(n_507),
.B(n_291),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_513),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_509),
.B(n_264),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_480),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_489),
.A2(n_269),
.B1(n_325),
.B2(n_213),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_480),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_475),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_465),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_463),
.B(n_402),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_480),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_513),
.Y(n_587)
);

INVxp33_ASAP7_75t_L g588 ( 
.A(n_478),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_502),
.B(n_505),
.C(n_485),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_507),
.A2(n_502),
.B1(n_505),
.B2(n_510),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_472),
.B(n_312),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_452),
.B(n_385),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_464),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_513),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_464),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_441),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_441),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_488),
.B(n_414),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_464),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_507),
.A2(n_430),
.B1(n_425),
.B2(n_338),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_478),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_L g602 ( 
.A1(n_452),
.A2(n_385),
.B1(n_387),
.B2(n_293),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_469),
.Y(n_603)
);

OAI22x1_ASAP7_75t_L g604 ( 
.A1(n_463),
.A2(n_427),
.B1(n_430),
.B2(n_204),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_441),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_488),
.B(n_388),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_488),
.B(n_389),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_469),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_469),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_469),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_489),
.A2(n_208),
.B1(n_204),
.B2(n_191),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_502),
.B(n_417),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_439),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_494),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_439),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_441),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_494),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_445),
.Y(n_618)
);

INVx8_ASAP7_75t_L g619 ( 
.A(n_453),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_442),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_445),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_453),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_451),
.Y(n_623)
);

AND3x2_ASAP7_75t_L g624 ( 
.A(n_477),
.B(n_290),
.C(n_433),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_442),
.Y(n_625)
);

CKINVDCx6p67_ASAP7_75t_R g626 ( 
.A(n_502),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_451),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_454),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_502),
.B(n_422),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_454),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_472),
.B(n_348),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_455),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_472),
.B(n_334),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_455),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_458),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_458),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_442),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_466),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_466),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_505),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_SL g641 ( 
.A(n_477),
.B(n_378),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_440),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_440),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_461),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_505),
.B(n_429),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_510),
.B(n_387),
.Y(n_646)
);

AND2x2_ASAP7_75t_SL g647 ( 
.A(n_515),
.B(n_218),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_461),
.B(n_474),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_442),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_440),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_510),
.B(n_369),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_510),
.B(n_416),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_510),
.B(n_405),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_440),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_477),
.A2(n_437),
.B1(n_436),
.B2(n_435),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_485),
.B(n_372),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_484),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_449),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_624),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_649),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_642),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_535),
.B(n_461),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_528),
.B(n_461),
.Y(n_663)
);

BUFx12f_ASAP7_75t_SL g664 ( 
.A(n_598),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_643),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_615),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_528),
.B(n_461),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_640),
.B(n_461),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_583),
.B(n_474),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_R g670 ( 
.A(n_641),
.B(n_174),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_649),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_584),
.B(n_598),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_526),
.B(n_474),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_526),
.B(n_474),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_633),
.A2(n_475),
.B(n_459),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_530),
.B(n_474),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_530),
.B(n_474),
.Y(n_677)
);

NOR3xp33_ASAP7_75t_L g678 ( 
.A(n_536),
.B(n_497),
.C(n_485),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_550),
.B(n_474),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_542),
.B(n_497),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_540),
.B(n_175),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_542),
.B(n_497),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_550),
.B(n_481),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_585),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_615),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_618),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_618),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_650),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_621),
.Y(n_689)
);

NOR2xp67_ASAP7_75t_L g690 ( 
.A(n_606),
.B(n_495),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_589),
.A2(n_468),
.B1(n_449),
.B2(n_475),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_590),
.B(n_481),
.Y(n_692)
);

AND2x2_ASAP7_75t_SL g693 ( 
.A(n_647),
.B(n_577),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_589),
.B(n_481),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_650),
.A2(n_468),
.B1(n_449),
.B2(n_500),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_551),
.B(n_481),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_612),
.A2(n_500),
.B1(n_211),
.B2(n_210),
.Y(n_697)
);

BUFx12f_ASAP7_75t_SL g698 ( 
.A(n_517),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_621),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_620),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_601),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_551),
.B(n_481),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_654),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_601),
.Y(n_704)
);

A2O1A1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_541),
.A2(n_500),
.B(n_492),
.C(n_511),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_588),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_548),
.B(n_175),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_620),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_656),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_579),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_556),
.B(n_481),
.Y(n_711)
);

BUFx8_ASAP7_75t_L g712 ( 
.A(n_652),
.Y(n_712)
);

NOR2xp67_ASAP7_75t_L g713 ( 
.A(n_607),
.B(n_496),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_556),
.B(n_481),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_654),
.Y(n_715)
);

OAI221xp5_ASAP7_75t_L g716 ( 
.A1(n_600),
.A2(n_514),
.B1(n_511),
.B2(n_496),
.C(n_499),
.Y(n_716)
);

INVxp67_ASAP7_75t_SL g717 ( 
.A(n_620),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_658),
.A2(n_449),
.B1(n_468),
.B2(n_481),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_658),
.B(n_449),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_613),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_613),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_569),
.A2(n_307),
.B1(n_341),
.B2(n_304),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_627),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_627),
.B(n_628),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_628),
.B(n_630),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_630),
.B(n_468),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_646),
.B(n_525),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_623),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_632),
.B(n_468),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_632),
.B(n_498),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_529),
.B(n_176),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_533),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_635),
.B(n_498),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_623),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_635),
.B(n_498),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_575),
.B(n_219),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_544),
.B(n_499),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_636),
.B(n_498),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_634),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_636),
.B(n_501),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_638),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_519),
.A2(n_527),
.B1(n_538),
.B2(n_652),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_638),
.B(n_501),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_557),
.B(n_501),
.Y(n_744)
);

NAND2x1_ASAP7_75t_L g745 ( 
.A(n_625),
.B(n_453),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_572),
.B(n_503),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_626),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_592),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_557),
.B(n_226),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_604),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_562),
.B(n_570),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_634),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_629),
.B(n_503),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_639),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_562),
.B(n_501),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_570),
.B(n_504),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_571),
.B(n_233),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_639),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_626),
.A2(n_517),
.B1(n_645),
.B2(n_653),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_576),
.B(n_242),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_576),
.B(n_504),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_523),
.B(n_514),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_L g763 ( 
.A(n_519),
.B(n_176),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_516),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_580),
.B(n_252),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_580),
.B(n_504),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_516),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_519),
.B(n_527),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_651),
.B(n_416),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_602),
.B(n_177),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_582),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_565),
.A2(n_515),
.B(n_508),
.C(n_432),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_604),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_582),
.B(n_508),
.Y(n_774)
);

AO221x1_ASAP7_75t_L g775 ( 
.A1(n_563),
.A2(n_322),
.B1(n_260),
.B2(n_266),
.C(n_289),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_586),
.B(n_292),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_586),
.B(n_296),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_545),
.B(n_177),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_572),
.A2(n_209),
.B1(n_179),
.B2(n_344),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_546),
.B(n_179),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_655),
.B(n_318),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_520),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_647),
.B(n_443),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_519),
.A2(n_492),
.B1(n_319),
.B2(n_339),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_657),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_519),
.A2(n_310),
.B1(n_309),
.B2(n_491),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_519),
.A2(n_491),
.B1(n_484),
.B2(n_256),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_611),
.A2(n_428),
.B(n_419),
.C(n_421),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_647),
.B(n_443),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_625),
.B(n_443),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_657),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_533),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_547),
.B(n_419),
.C(n_421),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_611),
.B(n_581),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_581),
.A2(n_432),
.B(n_423),
.C(n_426),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_520),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_625),
.B(n_443),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_L g798 ( 
.A(n_519),
.B(n_182),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_591),
.B(n_182),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_599),
.A2(n_436),
.B(n_423),
.C(n_426),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_552),
.B(n_188),
.Y(n_801)
);

NAND2x1_ASAP7_75t_L g802 ( 
.A(n_637),
.B(n_518),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_614),
.B(n_428),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_522),
.Y(n_804)
);

OAI221xp5_ASAP7_75t_L g805 ( 
.A1(n_599),
.A2(n_435),
.B1(n_437),
.B2(n_486),
.C(n_487),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_637),
.B(n_456),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_L g807 ( 
.A(n_527),
.B(n_538),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_527),
.A2(n_491),
.B1(n_484),
.B2(n_256),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_533),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_637),
.B(n_456),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_631),
.B(n_456),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_522),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_614),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_524),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_552),
.B(n_188),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_617),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_661),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_666),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_794),
.A2(n_538),
.B1(n_527),
.B2(n_617),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_701),
.B(n_517),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_732),
.B(n_552),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_710),
.B(n_527),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_666),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_732),
.B(n_552),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_672),
.B(n_517),
.Y(n_825)
);

CKINVDCx11_ASAP7_75t_R g826 ( 
.A(n_706),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_732),
.B(n_552),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_727),
.A2(n_517),
.B1(n_538),
.B2(n_527),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_664),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_747),
.B(n_560),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_685),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_705),
.A2(n_648),
.B(n_610),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_747),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_660),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_732),
.B(n_622),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_792),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_664),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_680),
.B(n_327),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_792),
.B(n_622),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_693),
.A2(n_560),
.B1(n_578),
.B2(n_587),
.Y(n_840)
);

BUFx12f_ASAP7_75t_L g841 ( 
.A(n_659),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_792),
.B(n_622),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_665),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_681),
.B(n_538),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_685),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_681),
.B(n_538),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_704),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_688),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_712),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_686),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_703),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_792),
.B(n_622),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_660),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_707),
.B(n_608),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_660),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_809),
.B(n_622),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_707),
.B(n_610),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_670),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_753),
.B(n_537),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_693),
.A2(n_564),
.B1(n_537),
.B2(n_539),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_660),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_686),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_682),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_715),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_687),
.Y(n_865)
);

NOR3xp33_ASAP7_75t_SL g866 ( 
.A(n_770),
.B(n_187),
.C(n_186),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_803),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_771),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_746),
.B(n_578),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_684),
.B(n_531),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_809),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_SL g872 ( 
.A1(n_813),
.A2(n_191),
.B1(n_187),
.B2(n_186),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_720),
.B(n_539),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_671),
.Y(n_874)
);

BUFx8_ASAP7_75t_L g875 ( 
.A(n_737),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_769),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_687),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_721),
.B(n_549),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_769),
.Y(n_879)
);

NAND2xp33_ASAP7_75t_SL g880 ( 
.A(n_670),
.B(n_189),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_770),
.B(n_193),
.C(n_189),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_709),
.B(n_748),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_769),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_809),
.B(n_622),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_712),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_775),
.A2(n_567),
.B1(n_549),
.B2(n_553),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_723),
.B(n_553),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_727),
.A2(n_587),
.B1(n_594),
.B2(n_210),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_671),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_712),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_781),
.B(n_327),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_692),
.A2(n_567),
.B1(n_554),
.B2(n_555),
.Y(n_892)
);

INVx5_ASAP7_75t_L g893 ( 
.A(n_809),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_690),
.A2(n_594),
.B1(n_531),
.B2(n_543),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_802),
.Y(n_895)
);

NAND3xp33_ASAP7_75t_L g896 ( 
.A(n_731),
.B(n_224),
.C(n_217),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_669),
.A2(n_619),
.B(n_533),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_746),
.B(n_486),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_713),
.A2(n_644),
.B1(n_543),
.B2(n_531),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_689),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_741),
.B(n_554),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_663),
.A2(n_619),
.B(n_533),
.Y(n_902)
);

BUFx12f_ASAP7_75t_L g903 ( 
.A(n_746),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_724),
.B(n_555),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_762),
.B(n_487),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_689),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_816),
.B(n_208),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_699),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_678),
.B(n_470),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_750),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_662),
.B(n_531),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_793),
.B(n_470),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_667),
.A2(n_619),
.B(n_644),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_725),
.B(n_561),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_759),
.B(n_543),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_700),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_799),
.B(n_561),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_799),
.B(n_564),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_728),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_754),
.B(n_471),
.Y(n_920)
);

AND2x2_ASAP7_75t_SL g921 ( 
.A(n_731),
.B(n_644),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_758),
.B(n_471),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_788),
.A2(n_212),
.B(n_324),
.C(n_325),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_778),
.B(n_327),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_700),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_717),
.B(n_566),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_728),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_734),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_773),
.B(n_543),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_783),
.B(n_644),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_734),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_692),
.A2(n_694),
.B1(n_752),
.B2(n_739),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_788),
.A2(n_568),
.B(n_573),
.C(n_609),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_789),
.B(n_518),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_778),
.B(n_568),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_739),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_708),
.B(n_518),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_691),
.A2(n_209),
.B1(n_196),
.B2(n_197),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_752),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_726),
.B(n_573),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_729),
.B(n_574),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_795),
.B(n_619),
.Y(n_942)
);

AND3x1_ASAP7_75t_L g943 ( 
.A(n_795),
.B(n_324),
.C(n_331),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_694),
.B(n_521),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_751),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_736),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_811),
.A2(n_619),
.B(n_616),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_695),
.B(n_593),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_764),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_764),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_767),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_742),
.B(n_521),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_736),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_SL g954 ( 
.A(n_745),
.B(n_193),
.Y(n_954)
);

NAND3xp33_ASAP7_75t_L g955 ( 
.A(n_780),
.B(n_313),
.C(n_228),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_780),
.B(n_595),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_730),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_675),
.B(n_521),
.Y(n_958)
);

CKINVDCx8_ASAP7_75t_R g959 ( 
.A(n_722),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_719),
.Y(n_960)
);

NOR2x2_ASAP7_75t_L g961 ( 
.A(n_697),
.B(n_256),
.Y(n_961)
);

OR2x6_ASAP7_75t_L g962 ( 
.A(n_719),
.B(n_595),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_779),
.B(n_716),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_767),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_698),
.B(n_603),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_782),
.Y(n_966)
);

OAI22xp33_ASAP7_75t_L g967 ( 
.A1(n_805),
.A2(n_331),
.B1(n_213),
.B2(n_335),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_782),
.Y(n_968)
);

AND2x6_ASAP7_75t_L g969 ( 
.A(n_698),
.B(n_603),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_733),
.B(n_609),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_705),
.B(n_749),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_735),
.B(n_558),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_SL g973 ( 
.A1(n_768),
.A2(n_807),
.B1(n_763),
.B2(n_798),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_757),
.Y(n_974)
);

AND2x2_ASAP7_75t_SL g975 ( 
.A(n_768),
.B(n_484),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_757),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_796),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_738),
.B(n_558),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_796),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_740),
.B(n_558),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_743),
.A2(n_335),
.B1(n_336),
.B2(n_342),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_804),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_804),
.B(n_559),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_673),
.B(n_559),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_812),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_812),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_760),
.Y(n_987)
);

BUFx4f_ASAP7_75t_L g988 ( 
.A(n_785),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_814),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_674),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_676),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_814),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_677),
.B(n_559),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_668),
.A2(n_616),
.B(n_605),
.Y(n_994)
);

NAND3xp33_ASAP7_75t_L g995 ( 
.A(n_760),
.B(n_306),
.C(n_232),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_765),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_791),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_679),
.B(n_596),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_683),
.B(n_596),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_696),
.B(n_596),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_817),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_945),
.B(n_859),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_867),
.B(n_801),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_SL g1004 ( 
.A(n_881),
.B(n_800),
.C(n_772),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_905),
.B(n_702),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_825),
.B(n_959),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_905),
.B(n_711),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_863),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_847),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_963),
.A2(n_924),
.B(n_953),
.C(n_946),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_871),
.A2(n_790),
.B(n_810),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_L g1012 ( 
.A(n_882),
.B(n_808),
.C(n_787),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_950),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_871),
.A2(n_806),
.B(n_797),
.Y(n_1014)
);

INVxp67_ASAP7_75t_L g1015 ( 
.A(n_863),
.Y(n_1015)
);

AO21x1_ASAP7_75t_L g1016 ( 
.A1(n_915),
.A2(n_765),
.B(n_776),
.Y(n_1016)
);

OA22x2_ASAP7_75t_L g1017 ( 
.A1(n_872),
.A2(n_336),
.B1(n_342),
.B2(n_251),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_882),
.B(n_988),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_L g1019 ( 
.A(n_836),
.B(n_714),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_843),
.Y(n_1020)
);

INVxp33_ASAP7_75t_SL g1021 ( 
.A(n_837),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_883),
.B(n_801),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_838),
.B(n_800),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_921),
.A2(n_784),
.B1(n_718),
.B2(n_786),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_848),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_950),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_935),
.B(n_744),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_891),
.B(n_776),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_907),
.B(n_815),
.Y(n_1029)
);

OAI22x1_ASAP7_75t_L g1030 ( 
.A1(n_876),
.A2(n_268),
.B1(n_236),
.B2(n_240),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_879),
.B(n_815),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_935),
.B(n_755),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_826),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_910),
.B(n_777),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_SL g1035 ( 
.A(n_955),
.B(n_896),
.C(n_866),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_870),
.B(n_756),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_R g1037 ( 
.A(n_858),
.B(n_761),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_851),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_864),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_929),
.B(n_766),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_837),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_L g1042 ( 
.A(n_866),
.B(n_880),
.C(n_981),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_988),
.B(n_774),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_829),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_908),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_929),
.B(n_597),
.Y(n_1046)
);

AOI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_938),
.A2(n_277),
.B(n_241),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_982),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_921),
.B(n_197),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_957),
.B(n_597),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_836),
.Y(n_1051)
);

OA22x2_ASAP7_75t_L g1052 ( 
.A1(n_961),
.A2(n_301),
.B1(n_323),
.B2(n_321),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_981),
.B(n_898),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_987),
.B(n_244),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_974),
.A2(n_605),
.B(n_330),
.C(n_326),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_927),
.Y(n_1056)
);

INVx6_ASAP7_75t_L g1057 ( 
.A(n_875),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_995),
.B(n_198),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_971),
.A2(n_909),
.B1(n_960),
.B2(n_957),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_868),
.B(n_524),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_987),
.B(n_253),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_952),
.A2(n_534),
.B(n_532),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_875),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_928),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_931),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_893),
.A2(n_911),
.B(n_897),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_982),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_898),
.B(n_491),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_833),
.B(n_254),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_819),
.A2(n_198),
.B1(n_205),
.B2(n_344),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_854),
.B(n_450),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_893),
.B(n_205),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_911),
.A2(n_326),
.B(n_340),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_819),
.A2(n_207),
.B1(n_340),
.B2(n_333),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_902),
.A2(n_333),
.B(n_330),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_996),
.B(n_281),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_857),
.B(n_207),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_913),
.A2(n_930),
.B(n_958),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_996),
.B(n_305),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_833),
.B(n_308),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_976),
.A2(n_211),
.B(n_214),
.C(n_5),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_834),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_958),
.A2(n_453),
.B(n_85),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_985),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_948),
.A2(n_453),
.B1(n_3),
.B2(n_5),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_939),
.Y(n_1086)
);

INVxp67_ASAP7_75t_SL g1087 ( 
.A(n_874),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_990),
.B(n_2),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_990),
.B(n_7),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_991),
.B(n_7),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_934),
.A2(n_453),
.B(n_92),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_834),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_844),
.A2(n_846),
.B(n_822),
.C(n_956),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_940),
.A2(n_78),
.B(n_163),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_R g1095 ( 
.A(n_885),
.B(n_69),
.Y(n_1095)
);

O2A1O1Ixp5_ASAP7_75t_L g1096 ( 
.A1(n_917),
.A2(n_93),
.B(n_152),
.C(n_149),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_967),
.A2(n_8),
.B1(n_25),
.B2(n_27),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_SL g1098 ( 
.A(n_923),
.B(n_25),
.C(n_28),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_991),
.B(n_28),
.Y(n_1099)
);

OR2x6_ASAP7_75t_L g1100 ( 
.A(n_890),
.B(n_104),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_841),
.B(n_29),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_985),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_923),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_L g1104 ( 
.A(n_967),
.B(n_888),
.C(n_849),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_903),
.B(n_31),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_874),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_918),
.A2(n_32),
.B(n_36),
.C(n_37),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_997),
.B(n_37),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_941),
.A2(n_904),
.B(n_914),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_969),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_890),
.B(n_115),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_889),
.B(n_39),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_989),
.Y(n_1113)
);

NOR3xp33_ASAP7_75t_SL g1114 ( 
.A(n_954),
.B(n_965),
.C(n_840),
.Y(n_1114)
);

AOI221x1_ASAP7_75t_L g1115 ( 
.A1(n_832),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.C(n_44),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_947),
.A2(n_125),
.B(n_148),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_869),
.B(n_120),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_869),
.B(n_117),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_932),
.A2(n_127),
.B1(n_145),
.B2(n_140),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_932),
.A2(n_109),
.B1(n_138),
.B2(n_135),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_828),
.A2(n_41),
.B(n_45),
.C(n_46),
.Y(n_1121)
);

O2A1O1Ixp5_ASAP7_75t_L g1122 ( 
.A1(n_934),
.A2(n_114),
.B(n_131),
.C(n_166),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_853),
.Y(n_1123)
);

CKINVDCx10_ASAP7_75t_R g1124 ( 
.A(n_820),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_933),
.A2(n_994),
.B(n_993),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_975),
.A2(n_48),
.B1(n_54),
.B2(n_973),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_989),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_903),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_912),
.B(n_920),
.Y(n_1129)
);

AO22x1_ASAP7_75t_L g1130 ( 
.A1(n_969),
.A2(n_830),
.B1(n_912),
.B2(n_853),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_969),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_943),
.Y(n_1132)
);

AOI222xp33_ASAP7_75t_L g1133 ( 
.A1(n_920),
.A2(n_922),
.B1(n_830),
.B2(n_944),
.C1(n_966),
.C2(n_977),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_972),
.A2(n_978),
.B(n_980),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_SL g1135 ( 
.A1(n_886),
.A2(n_999),
.B(n_984),
.C(n_855),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_SL g1136 ( 
.A1(n_944),
.A2(n_937),
.B(n_993),
.C(n_821),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_969),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_992),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1066),
.A2(n_1000),
.B(n_998),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_1016),
.A2(n_999),
.A3(n_984),
.B(n_970),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1001),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_SL g1142 ( 
.A1(n_1024),
.A2(n_820),
.B(n_942),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1109),
.A2(n_926),
.B(n_820),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_1129),
.B(n_855),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1044),
.Y(n_1145)
);

AOI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1097),
.A2(n_1047),
.B1(n_1107),
.B2(n_1103),
.C(n_1042),
.Y(n_1146)
);

AOI211x1_ASAP7_75t_L g1147 ( 
.A1(n_1126),
.A2(n_901),
.B(n_878),
.C(n_873),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_SL g1148 ( 
.A1(n_1010),
.A2(n_942),
.B(n_899),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_1093),
.A2(n_886),
.B(n_860),
.Y(n_1149)
);

AOI211x1_ASAP7_75t_L g1150 ( 
.A1(n_1020),
.A2(n_1025),
.B(n_1039),
.C(n_1038),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1027),
.A2(n_827),
.B(n_835),
.Y(n_1151)
);

BUFx4f_ASAP7_75t_SL g1152 ( 
.A(n_1033),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1018),
.A2(n_887),
.B(n_937),
.C(n_925),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1053),
.B(n_861),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1026),
.Y(n_1155)
);

OAI22x1_ASAP7_75t_L g1156 ( 
.A1(n_1132),
.A2(n_861),
.B1(n_823),
.B2(n_936),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1011),
.A2(n_892),
.B(n_983),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1029),
.A2(n_916),
.B(n_894),
.C(n_818),
.Y(n_1158)
);

NAND3x1_ASAP7_75t_L g1159 ( 
.A(n_1101),
.B(n_916),
.C(n_968),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_1057),
.B(n_962),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_SL g1161 ( 
.A1(n_1059),
.A2(n_823),
.B(n_936),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1032),
.A2(n_824),
.B(n_856),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1009),
.Y(n_1163)
);

BUFx12f_ASAP7_75t_L g1164 ( 
.A(n_1057),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1002),
.B(n_862),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1036),
.A2(n_900),
.B(n_831),
.Y(n_1166)
);

OA21x2_ASAP7_75t_L g1167 ( 
.A1(n_1096),
.A2(n_845),
.B(n_831),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1006),
.A2(n_969),
.B1(n_962),
.B2(n_906),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1135),
.A2(n_824),
.B(n_835),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1008),
.B(n_900),
.Y(n_1170)
);

INVx3_ASAP7_75t_SL g1171 ( 
.A(n_1128),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1014),
.A2(n_862),
.B(n_919),
.Y(n_1172)
);

BUFx12f_ASAP7_75t_L g1173 ( 
.A(n_1063),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1115),
.A2(n_949),
.A3(n_951),
.B(n_845),
.Y(n_1174)
);

AOI221x1_ASAP7_75t_L g1175 ( 
.A1(n_1104),
.A2(n_949),
.B1(n_951),
.B2(n_850),
.C(n_919),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1028),
.B(n_865),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_1008),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1062),
.A2(n_906),
.B(n_877),
.Y(n_1178)
);

OR2x6_ASAP7_75t_L g1179 ( 
.A(n_1130),
.B(n_962),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1037),
.B(n_968),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1031),
.A2(n_877),
.B(n_850),
.C(n_865),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1059),
.B(n_1040),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1116),
.A2(n_992),
.B(n_986),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1005),
.B(n_986),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1136),
.A2(n_839),
.B(n_842),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1071),
.A2(n_1019),
.B(n_1046),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1004),
.A2(n_979),
.B(n_964),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1050),
.A2(n_1083),
.B(n_1060),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1003),
.B(n_895),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1007),
.B(n_1023),
.Y(n_1190)
);

OAI21xp33_ASAP7_75t_L g1191 ( 
.A1(n_1054),
.A2(n_839),
.B(n_842),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1077),
.B(n_895),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1091),
.A2(n_852),
.B(n_856),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_SL g1194 ( 
.A1(n_1097),
.A2(n_1085),
.B(n_1103),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_SL g1195 ( 
.A1(n_1121),
.A2(n_852),
.B(n_884),
.C(n_895),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1043),
.A2(n_884),
.B(n_895),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1087),
.B(n_1045),
.Y(n_1197)
);

AOI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1049),
.A2(n_1075),
.B(n_1112),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1087),
.B(n_1056),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_1051),
.Y(n_1200)
);

BUFx4_ASAP7_75t_SL g1201 ( 
.A(n_1100),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_SL g1202 ( 
.A1(n_1131),
.A2(n_1120),
.B(n_1119),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1203)
);

OAI21xp33_ASAP7_75t_L g1204 ( 
.A1(n_1061),
.A2(n_1076),
.B(n_1079),
.Y(n_1204)
);

OAI22x1_ASAP7_75t_L g1205 ( 
.A1(n_1132),
.A2(n_1022),
.B1(n_1108),
.B2(n_1015),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1122),
.A2(n_1067),
.B(n_1138),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1048),
.A2(n_1084),
.B(n_1127),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1102),
.A2(n_1113),
.B(n_1094),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1086),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1004),
.A2(n_1114),
.B(n_1012),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1082),
.A2(n_1123),
.B(n_1092),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1069),
.B(n_1015),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1131),
.A2(n_1137),
.B(n_1110),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1133),
.A2(n_1117),
.B(n_1118),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1106),
.B(n_1068),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1041),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1100),
.B(n_1111),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_SL g1218 ( 
.A1(n_1110),
.A2(n_1137),
.B(n_1051),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1072),
.A2(n_1089),
.B(n_1090),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1095),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1106),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1082),
.A2(n_1123),
.B(n_1092),
.Y(n_1222)
);

O2A1O1Ixp5_ASAP7_75t_L g1223 ( 
.A1(n_1088),
.A2(n_1099),
.B(n_1055),
.C(n_1073),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1104),
.B(n_1108),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1100),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1034),
.B(n_1080),
.Y(n_1226)
);

AOI21xp33_ASAP7_75t_L g1227 ( 
.A1(n_1107),
.A2(n_1085),
.B(n_1074),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1051),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1051),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1035),
.A2(n_1058),
.B(n_1070),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1110),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1114),
.B(n_1137),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1110),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1081),
.A2(n_1111),
.B(n_1030),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1017),
.A2(n_1105),
.B(n_1052),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1098),
.B(n_1021),
.Y(n_1236)
);

BUFx12f_ASAP7_75t_L g1237 ( 
.A(n_1111),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1124),
.A2(n_1109),
.B(n_893),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1013),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1110),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1016),
.A2(n_1078),
.A3(n_1093),
.B(n_1115),
.Y(n_1241)
);

NOR2xp67_ASAP7_75t_L g1242 ( 
.A(n_1035),
.B(n_867),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1093),
.A2(n_1109),
.B(n_1134),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1093),
.A2(n_1109),
.B(n_1134),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1002),
.B(n_945),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1110),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1051),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1093),
.A2(n_1109),
.B(n_1134),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1010),
.A2(n_684),
.B(n_1018),
.C(n_452),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1002),
.B(n_945),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1066),
.A2(n_1125),
.B(n_1078),
.Y(n_1251)
);

AOI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1066),
.A2(n_915),
.B(n_1078),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1051),
.Y(n_1253)
);

AOI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1066),
.A2(n_915),
.B(n_1078),
.Y(n_1254)
);

INVx4_ASAP7_75t_L g1255 ( 
.A(n_1051),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1002),
.B(n_945),
.Y(n_1256)
);

AO32x2_ASAP7_75t_L g1257 ( 
.A1(n_1126),
.A2(n_1120),
.A3(n_1119),
.B1(n_1074),
.B2(n_1070),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1002),
.B(n_945),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1110),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1002),
.B(n_945),
.Y(n_1260)
);

OAI21xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1085),
.A2(n_1002),
.B(n_693),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1059),
.A2(n_1085),
.B1(n_1097),
.B2(n_1002),
.Y(n_1262)
);

NOR2x1_ASAP7_75t_SL g1263 ( 
.A(n_1131),
.B(n_820),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1042),
.B(n_881),
.C(n_924),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1002),
.B(n_945),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1002),
.B(n_945),
.Y(n_1266)
);

OAI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1194),
.A2(n_1224),
.B1(n_1262),
.B2(n_1265),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1204),
.A2(n_1219),
.B(n_1223),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1252),
.A2(n_1254),
.B(n_1251),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1212),
.B(n_1176),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1245),
.B(n_1250),
.Y(n_1271)
);

BUFx8_ASAP7_75t_L g1272 ( 
.A(n_1164),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1228),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1207),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1154),
.B(n_1144),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1190),
.B(n_1224),
.Y(n_1276)
);

AO21x2_ASAP7_75t_L g1277 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1244),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1226),
.A2(n_1227),
.B(n_1249),
.C(n_1210),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1155),
.Y(n_1279)
);

NAND2x1p5_ASAP7_75t_L g1280 ( 
.A(n_1177),
.B(n_1217),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1146),
.B(n_1214),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1264),
.A2(n_1146),
.B(n_1210),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1194),
.A2(n_1261),
.B(n_1227),
.C(n_1262),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1239),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1163),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1143),
.A2(n_1202),
.B(n_1186),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1256),
.B(n_1258),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1160),
.B(n_1233),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1139),
.A2(n_1172),
.B(n_1157),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1216),
.Y(n_1290)
);

AOI22x1_ASAP7_75t_L g1291 ( 
.A1(n_1205),
.A2(n_1238),
.B1(n_1234),
.B2(n_1156),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1228),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1188),
.A2(n_1183),
.B(n_1208),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1190),
.B(n_1182),
.Y(n_1294)
);

NAND2x1p5_ASAP7_75t_L g1295 ( 
.A(n_1177),
.B(n_1217),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1256),
.B(n_1258),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1145),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1230),
.A2(n_1192),
.B(n_1158),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1203),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1228),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1220),
.A2(n_1237),
.B1(n_1236),
.B2(n_1225),
.Y(n_1301)
);

BUFx12f_ASAP7_75t_L g1302 ( 
.A(n_1173),
.Y(n_1302)
);

AOI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1260),
.A2(n_1265),
.B1(n_1266),
.B2(n_1236),
.C(n_1182),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1203),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1178),
.A2(n_1206),
.B(n_1185),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1167),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1175),
.A2(n_1169),
.A3(n_1193),
.B(n_1181),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1167),
.Y(n_1308)
);

NAND2x1p5_ASAP7_75t_L g1309 ( 
.A(n_1233),
.B(n_1189),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1187),
.A2(n_1162),
.B(n_1193),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1148),
.A2(n_1142),
.B(n_1161),
.Y(n_1311)
);

NAND2x1p5_ASAP7_75t_L g1312 ( 
.A(n_1211),
.B(n_1222),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1151),
.A2(n_1196),
.A3(n_1232),
.B(n_1263),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1209),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1260),
.B(n_1266),
.Y(n_1315)
);

AO21x2_ASAP7_75t_L g1316 ( 
.A1(n_1187),
.A2(n_1198),
.B(n_1166),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1150),
.Y(n_1317)
);

INVx5_ASAP7_75t_L g1318 ( 
.A(n_1247),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1242),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1191),
.A2(n_1153),
.B(n_1196),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1170),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1168),
.A2(n_1159),
.B(n_1232),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1215),
.B(n_1165),
.Y(n_1323)
);

BUFx12f_ASAP7_75t_L g1324 ( 
.A(n_1247),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1221),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1197),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1149),
.A2(n_1199),
.B(n_1184),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1165),
.A2(n_1241),
.B(n_1235),
.Y(n_1328)
);

OAI221xp5_ASAP7_75t_L g1329 ( 
.A1(n_1171),
.A2(n_1160),
.B1(n_1180),
.B2(n_1195),
.C(n_1179),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1213),
.A2(n_1218),
.B(n_1246),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1229),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1240),
.A2(n_1259),
.B(n_1246),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1241),
.A2(n_1140),
.B(n_1179),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1174),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1247),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1174),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1253),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1140),
.A2(n_1179),
.B(n_1147),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1253),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1174),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1231),
.B(n_1200),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1253),
.Y(n_1342)
);

CKINVDCx11_ASAP7_75t_R g1343 ( 
.A(n_1152),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1140),
.A2(n_1257),
.B(n_1231),
.Y(n_1344)
);

OR2x6_ASAP7_75t_L g1345 ( 
.A(n_1231),
.B(n_1200),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1257),
.A2(n_1255),
.B(n_1201),
.Y(n_1346)
);

AO221x2_ASAP7_75t_L g1347 ( 
.A1(n_1257),
.A2(n_1255),
.B1(n_1194),
.B2(n_1205),
.C(n_1224),
.Y(n_1347)
);

O2A1O1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1204),
.A2(n_1224),
.B(n_1226),
.C(n_1010),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_SL g1349 ( 
.A1(n_1263),
.A2(n_1214),
.B(n_1234),
.Y(n_1349)
);

OR2x6_ASAP7_75t_L g1350 ( 
.A(n_1179),
.B(n_1142),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1207),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1216),
.Y(n_1352)
);

OAI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1194),
.A2(n_1224),
.B1(n_1115),
.B2(n_1262),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1177),
.B(n_1131),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_SL g1355 ( 
.A1(n_1224),
.A2(n_1121),
.B(n_1227),
.C(n_1232),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1207),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1233),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1141),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1207),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1204),
.A2(n_1219),
.B(n_1010),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1204),
.B(n_684),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1244),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1204),
.B(n_684),
.Y(n_1363)
);

OR2x6_ASAP7_75t_L g1364 ( 
.A(n_1179),
.B(n_1142),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1212),
.B(n_672),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1141),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1154),
.B(n_1160),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1141),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1141),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1141),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1212),
.B(n_672),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1204),
.A2(n_1219),
.B(n_1010),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_SL g1373 ( 
.A1(n_1224),
.A2(n_1121),
.B(n_1227),
.C(n_1232),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1163),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1204),
.A2(n_1224),
.B1(n_959),
.B2(n_1266),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1245),
.B(n_1250),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1163),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1163),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1207),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_1152),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1204),
.A2(n_1219),
.B(n_1010),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1207),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1177),
.B(n_1131),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1281),
.A2(n_1375),
.B(n_1282),
.C(n_1363),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1315),
.B(n_1326),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1361),
.B(n_1363),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1270),
.B(n_1275),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1365),
.B(n_1371),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1315),
.A2(n_1287),
.B1(n_1376),
.B2(n_1296),
.Y(n_1389)
);

INVx5_ASAP7_75t_L g1390 ( 
.A(n_1350),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1325),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1276),
.B(n_1303),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1281),
.A2(n_1283),
.B1(n_1361),
.B2(n_1353),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1380),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1326),
.B(n_1267),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1321),
.B(n_1347),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1348),
.A2(n_1278),
.B(n_1319),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1283),
.A2(n_1353),
.B1(n_1267),
.B2(n_1304),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1360),
.A2(n_1381),
.B(n_1372),
.C(n_1355),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1355),
.A2(n_1373),
.B(n_1268),
.C(n_1329),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1323),
.B(n_1299),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1347),
.B(n_1280),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1347),
.B(n_1294),
.Y(n_1403)
);

OAI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1286),
.A2(n_1291),
.B1(n_1298),
.B2(n_1322),
.C(n_1301),
.Y(n_1404)
);

AOI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1373),
.A2(n_1320),
.B1(n_1294),
.B2(n_1349),
.C(n_1285),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1374),
.A2(n_1378),
.B(n_1290),
.C(n_1309),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1280),
.B(n_1295),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1309),
.A2(n_1368),
.B(n_1314),
.C(n_1370),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1305),
.A2(n_1289),
.B(n_1269),
.Y(n_1409)
);

NOR2xp67_ASAP7_75t_L g1410 ( 
.A(n_1279),
.B(n_1284),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1358),
.B(n_1366),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1369),
.A2(n_1377),
.B(n_1297),
.C(n_1383),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1352),
.B(n_1377),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1331),
.B(n_1277),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1330),
.B(n_1346),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1328),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1277),
.B(n_1362),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1380),
.Y(n_1418)
);

NOR2xp67_ASAP7_75t_L g1419 ( 
.A(n_1302),
.B(n_1357),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1341),
.B(n_1350),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1354),
.A2(n_1383),
.B(n_1364),
.C(n_1350),
.Y(n_1421)
);

NOR2x1_ASAP7_75t_L g1422 ( 
.A(n_1357),
.B(n_1345),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1362),
.A2(n_1364),
.B(n_1345),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1324),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1346),
.B(n_1335),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1327),
.Y(n_1426)
);

O2A1O1Ixp5_ASAP7_75t_L g1427 ( 
.A1(n_1334),
.A2(n_1336),
.B(n_1340),
.C(n_1382),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1337),
.B(n_1342),
.Y(n_1428)
);

AOI21x1_ASAP7_75t_SL g1429 ( 
.A1(n_1272),
.A2(n_1338),
.B(n_1313),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1364),
.A2(n_1344),
.B1(n_1318),
.B2(n_1334),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1339),
.B(n_1344),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1344),
.B(n_1273),
.Y(n_1432)
);

AND2x2_ASAP7_75t_SL g1433 ( 
.A(n_1310),
.B(n_1300),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1318),
.A2(n_1345),
.B1(n_1302),
.B2(n_1324),
.Y(n_1434)
);

O2A1O1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1311),
.A2(n_1382),
.B(n_1379),
.C(n_1359),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1313),
.B(n_1333),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1343),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1273),
.A2(n_1292),
.B(n_1300),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1318),
.A2(n_1292),
.B1(n_1343),
.B2(n_1312),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1292),
.B(n_1332),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1313),
.B(n_1316),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1274),
.A2(n_1356),
.B(n_1351),
.C(n_1312),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1318),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1351),
.A2(n_1308),
.B1(n_1306),
.B2(n_1307),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1306),
.A2(n_1308),
.B1(n_1307),
.B2(n_1313),
.Y(n_1445)
);

OA22x2_ASAP7_75t_L g1446 ( 
.A1(n_1293),
.A2(n_1282),
.B1(n_1115),
.B2(n_1194),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1343),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1288),
.B(n_1367),
.Y(n_1448)
);

AND2x6_ASAP7_75t_L g1449 ( 
.A(n_1317),
.B(n_1232),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1268),
.A2(n_1305),
.B(n_1289),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1315),
.B(n_1271),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1315),
.A2(n_1097),
.B1(n_1194),
.B2(n_1085),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1315),
.B(n_1326),
.Y(n_1453)
);

O2A1O1Ixp5_ASAP7_75t_L g1454 ( 
.A1(n_1281),
.A2(n_1282),
.B(n_1227),
.C(n_1353),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1315),
.B(n_1326),
.Y(n_1455)
);

BUFx4f_ASAP7_75t_L g1456 ( 
.A(n_1302),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1276),
.B(n_1321),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1276),
.B(n_1321),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1325),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1343),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1315),
.A2(n_1097),
.B1(n_1194),
.B2(n_1085),
.Y(n_1461)
);

AOI221xp5_ASAP7_75t_L g1462 ( 
.A1(n_1281),
.A2(n_1204),
.B1(n_1282),
.B2(n_770),
.C(n_1375),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1315),
.A2(n_1097),
.B1(n_1194),
.B2(n_1085),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1270),
.B(n_1275),
.Y(n_1464)
);

O2A1O1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1281),
.A2(n_1204),
.B(n_1224),
.C(n_1375),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1414),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1440),
.B(n_1390),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1416),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1417),
.B(n_1431),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1433),
.B(n_1426),
.Y(n_1470)
);

INVx1_ASAP7_75t_SL g1471 ( 
.A(n_1459),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1415),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_1459),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1389),
.B(n_1385),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1389),
.B(n_1385),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1457),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1427),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1453),
.B(n_1455),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1445),
.B(n_1432),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1409),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1415),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1435),
.A2(n_1445),
.B(n_1429),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1396),
.B(n_1403),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1453),
.B(n_1455),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1391),
.Y(n_1485)
);

AOI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1393),
.A2(n_1398),
.B(n_1444),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1462),
.A2(n_1386),
.B1(n_1393),
.B2(n_1463),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1450),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1450),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1436),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1441),
.B(n_1402),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1451),
.B(n_1395),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1425),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1454),
.A2(n_1399),
.B(n_1384),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1411),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1430),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1442),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1423),
.B(n_1421),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1410),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1465),
.A2(n_1397),
.B(n_1400),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1390),
.Y(n_1501)
);

NOR2x1_ASAP7_75t_L g1502 ( 
.A(n_1408),
.B(n_1412),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1446),
.B(n_1398),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1437),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1446),
.B(n_1395),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1420),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1449),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1405),
.B(n_1448),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1404),
.A2(n_1392),
.B(n_1463),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1449),
.Y(n_1510)
);

NAND2x1_ASAP7_75t_L g1511 ( 
.A(n_1498),
.B(n_1422),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1471),
.Y(n_1512)
);

INVxp67_ASAP7_75t_L g1513 ( 
.A(n_1502),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1487),
.B(n_1452),
.C(n_1461),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1468),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1466),
.B(n_1458),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1468),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1472),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1469),
.B(n_1413),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1500),
.A2(n_1452),
.B1(n_1461),
.B2(n_1388),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1469),
.B(n_1401),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1466),
.B(n_1406),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1474),
.B(n_1407),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1479),
.B(n_1464),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1490),
.Y(n_1525)
);

INVxp67_ASAP7_75t_SL g1526 ( 
.A(n_1477),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1474),
.B(n_1428),
.Y(n_1527)
);

OAI221xp5_ASAP7_75t_L g1528 ( 
.A1(n_1500),
.A2(n_1456),
.B1(n_1439),
.B2(n_1434),
.C(n_1419),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1498),
.Y(n_1529)
);

OR2x6_ASAP7_75t_L g1530 ( 
.A(n_1498),
.B(n_1434),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1481),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1475),
.B(n_1387),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1480),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1470),
.B(n_1491),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1467),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1475),
.B(n_1493),
.Y(n_1536)
);

INVxp67_ASAP7_75t_SL g1537 ( 
.A(n_1513),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1532),
.B(n_1523),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1533),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1533),
.Y(n_1540)
);

OAI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1514),
.A2(n_1494),
.B1(n_1509),
.B2(n_1498),
.Y(n_1541)
);

AO21x2_ASAP7_75t_L g1542 ( 
.A1(n_1526),
.A2(n_1488),
.B(n_1489),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1514),
.A2(n_1494),
.B1(n_1509),
.B2(n_1502),
.Y(n_1543)
);

OAI221xp5_ASAP7_75t_L g1544 ( 
.A1(n_1513),
.A2(n_1509),
.B1(n_1498),
.B2(n_1492),
.C(n_1503),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1534),
.B(n_1491),
.Y(n_1545)
);

OAI33xp33_ASAP7_75t_L g1546 ( 
.A1(n_1522),
.A2(n_1492),
.A3(n_1485),
.B1(n_1493),
.B2(n_1483),
.B3(n_1495),
.Y(n_1546)
);

NAND4xp25_ASAP7_75t_SL g1547 ( 
.A(n_1520),
.B(n_1503),
.C(n_1505),
.D(n_1483),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1520),
.A2(n_1509),
.B1(n_1503),
.B2(n_1486),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1535),
.B(n_1472),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1534),
.B(n_1470),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1515),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1525),
.Y(n_1552)
);

OAI211xp5_ASAP7_75t_L g1553 ( 
.A1(n_1522),
.A2(n_1509),
.B(n_1486),
.C(n_1496),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_1519),
.Y(n_1554)
);

AOI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1536),
.A2(n_1505),
.B1(n_1476),
.B2(n_1485),
.C(n_1478),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1531),
.Y(n_1556)
);

OAI211xp5_ASAP7_75t_L g1557 ( 
.A1(n_1536),
.A2(n_1496),
.B(n_1505),
.C(n_1478),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1519),
.B(n_1476),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1531),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1530),
.B(n_1498),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1531),
.Y(n_1561)
);

BUFx2_ASAP7_75t_L g1562 ( 
.A(n_1535),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1530),
.A2(n_1508),
.B1(n_1507),
.B2(n_1506),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1532),
.A2(n_1508),
.B1(n_1484),
.B2(n_1507),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1515),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1524),
.B(n_1470),
.Y(n_1566)
);

AOI211xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1528),
.A2(n_1508),
.B(n_1438),
.C(n_1510),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1518),
.B(n_1472),
.Y(n_1568)
);

OAI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1528),
.A2(n_1530),
.B1(n_1507),
.B2(n_1511),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1527),
.B(n_1471),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1517),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1527),
.B(n_1473),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1523),
.A2(n_1516),
.B1(n_1526),
.B2(n_1484),
.C(n_1495),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_L g1574 ( 
.A(n_1511),
.B(n_1497),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1512),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1551),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1551),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1565),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1542),
.Y(n_1579)
);

CKINVDCx16_ASAP7_75t_R g1580 ( 
.A(n_1543),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1542),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1552),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1574),
.B(n_1529),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1565),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1575),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1574),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1571),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1537),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1556),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1568),
.B(n_1529),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1571),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1561),
.Y(n_1592)
);

NAND3xp33_ASAP7_75t_L g1593 ( 
.A(n_1543),
.B(n_1529),
.C(n_1499),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1538),
.B(n_1512),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1560),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1542),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1555),
.B(n_1524),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1554),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1539),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1573),
.B(n_1521),
.Y(n_1600)
);

INVx4_ASAP7_75t_SL g1601 ( 
.A(n_1560),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1558),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1561),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1560),
.B(n_1530),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1568),
.B(n_1560),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_SL g1606 ( 
.A1(n_1541),
.A2(n_1530),
.B(n_1501),
.Y(n_1606)
);

INVx4_ASAP7_75t_SL g1607 ( 
.A(n_1560),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1580),
.B(n_1562),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1576),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1580),
.B(n_1540),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1600),
.B(n_1570),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1586),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1576),
.Y(n_1613)
);

NAND2x1p5_ASAP7_75t_L g1614 ( 
.A(n_1586),
.B(n_1482),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_SL g1615 ( 
.A1(n_1589),
.A2(n_1548),
.B(n_1559),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1592),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1597),
.B(n_1570),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1596),
.Y(n_1618)
);

INVxp67_ASAP7_75t_SL g1619 ( 
.A(n_1596),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1596),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1601),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1577),
.B(n_1578),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1605),
.B(n_1562),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1598),
.B(n_1572),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1582),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1602),
.B(n_1588),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1579),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1585),
.B(n_1546),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1605),
.B(n_1549),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1577),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1579),
.Y(n_1631)
);

AOI222xp33_ASAP7_75t_SL g1632 ( 
.A1(n_1588),
.A2(n_1548),
.B1(n_1564),
.B2(n_1473),
.C1(n_1547),
.C2(n_1553),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1578),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1592),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1601),
.B(n_1549),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1605),
.B(n_1549),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1603),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1601),
.B(n_1550),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1593),
.B(n_1569),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1584),
.B(n_1557),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1587),
.B(n_1564),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1601),
.B(n_1550),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1581),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1587),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1591),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1601),
.B(n_1566),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1607),
.B(n_1545),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1622),
.Y(n_1648)
);

AO21x1_ASAP7_75t_L g1649 ( 
.A1(n_1628),
.A2(n_1583),
.B(n_1595),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1622),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1622),
.Y(n_1651)
);

OAI21xp33_ASAP7_75t_L g1652 ( 
.A1(n_1628),
.A2(n_1606),
.B(n_1547),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1625),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1609),
.Y(n_1654)
);

NAND2x2_ASAP7_75t_L g1655 ( 
.A(n_1616),
.B(n_1394),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1616),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1616),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1608),
.B(n_1590),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1626),
.B(n_1594),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1626),
.B(n_1558),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1609),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1613),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1616),
.B(n_1607),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1624),
.B(n_1519),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1624),
.B(n_1603),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1634),
.Y(n_1666)
);

INVxp67_ASAP7_75t_SL g1667 ( 
.A(n_1637),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1613),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1608),
.B(n_1590),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1630),
.Y(n_1670)
);

INVxp67_ASAP7_75t_SL g1671 ( 
.A(n_1637),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1611),
.B(n_1589),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1639),
.A2(n_1544),
.B1(n_1606),
.B2(n_1563),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1611),
.B(n_1599),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1637),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1617),
.B(n_1521),
.Y(n_1676)
);

NOR2xp67_ASAP7_75t_SL g1677 ( 
.A(n_1621),
.B(n_1447),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1617),
.B(n_1521),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1630),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1637),
.B(n_1607),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1633),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1608),
.B(n_1590),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1653),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1658),
.B(n_1621),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1653),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1669),
.B(n_1621),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1666),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1682),
.B(n_1646),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1666),
.B(n_1625),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1667),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1663),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1667),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1671),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1663),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1671),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1680),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1648),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1660),
.B(n_1640),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1675),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1657),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1650),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1680),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1652),
.A2(n_1639),
.B1(n_1595),
.B2(n_1604),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1656),
.B(n_1635),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1672),
.B(n_1640),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1651),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1656),
.B(n_1634),
.Y(n_1707)
);

AOI222xp33_ASAP7_75t_L g1708 ( 
.A1(n_1673),
.A2(n_1641),
.B1(n_1632),
.B2(n_1615),
.C1(n_1607),
.C2(n_1612),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1708),
.A2(n_1673),
.B(n_1610),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1690),
.Y(n_1710)
);

AOI21xp33_ASAP7_75t_L g1711 ( 
.A1(n_1687),
.A2(n_1649),
.B(n_1665),
.Y(n_1711)
);

OAI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1703),
.A2(n_1655),
.B1(n_1659),
.B2(n_1672),
.C(n_1677),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1698),
.A2(n_1610),
.B1(n_1635),
.B2(n_1595),
.Y(n_1713)
);

NOR2xp67_ASAP7_75t_SL g1714 ( 
.A(n_1696),
.B(n_1447),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1688),
.A2(n_1595),
.B1(n_1635),
.B2(n_1604),
.Y(n_1715)
);

AOI332xp33_ASAP7_75t_L g1716 ( 
.A1(n_1683),
.A2(n_1661),
.A3(n_1679),
.B1(n_1654),
.B2(n_1670),
.B3(n_1668),
.C1(n_1662),
.C2(n_1681),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1684),
.B(n_1646),
.Y(n_1717)
);

NOR2x1_ASAP7_75t_L g1718 ( 
.A(n_1690),
.B(n_1612),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1684),
.A2(n_1632),
.B1(n_1635),
.B2(n_1646),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1685),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1698),
.A2(n_1610),
.B1(n_1635),
.B2(n_1604),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1685),
.Y(n_1722)
);

OAI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1689),
.A2(n_1567),
.B1(n_1641),
.B2(n_1604),
.Y(n_1723)
);

AOI211xp5_ASAP7_75t_L g1724 ( 
.A1(n_1694),
.A2(n_1612),
.B(n_1647),
.C(n_1642),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1699),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1705),
.A2(n_1604),
.B1(n_1638),
.B2(n_1642),
.Y(n_1726)
);

OAI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1705),
.A2(n_1567),
.B1(n_1678),
.B2(n_1676),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1702),
.B(n_1674),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1717),
.B(n_1686),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1725),
.B(n_1702),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1710),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1720),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1725),
.B(n_1691),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1718),
.B(n_1699),
.Y(n_1734)
);

INVx2_ASAP7_75t_SL g1735 ( 
.A(n_1722),
.Y(n_1735)
);

NOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1709),
.B(n_1685),
.Y(n_1736)
);

INVxp67_ASAP7_75t_L g1737 ( 
.A(n_1714),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1728),
.B(n_1692),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1712),
.B(n_1691),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1724),
.B(n_1686),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1736),
.A2(n_1719),
.B1(n_1709),
.B2(n_1727),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1734),
.Y(n_1742)
);

NOR2x1p5_ASAP7_75t_L g1743 ( 
.A(n_1730),
.B(n_1696),
.Y(n_1743)
);

AOI322xp5_ASAP7_75t_L g1744 ( 
.A1(n_1739),
.A2(n_1711),
.A3(n_1740),
.B1(n_1723),
.B2(n_1731),
.C1(n_1734),
.C2(n_1738),
.Y(n_1744)
);

OAI21xp33_ASAP7_75t_L g1745 ( 
.A1(n_1729),
.A2(n_1715),
.B(n_1707),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1737),
.A2(n_1713),
.B(n_1721),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1738),
.A2(n_1683),
.B(n_1692),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1733),
.B(n_1693),
.Y(n_1748)
);

OAI211xp5_ASAP7_75t_L g1749 ( 
.A1(n_1735),
.A2(n_1716),
.B(n_1693),
.C(n_1695),
.Y(n_1749)
);

OAI211xp5_ASAP7_75t_L g1750 ( 
.A1(n_1732),
.A2(n_1695),
.B(n_1696),
.C(n_1699),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_SL g1751 ( 
.A1(n_1740),
.A2(n_1726),
.B1(n_1696),
.B2(n_1688),
.Y(n_1751)
);

NOR2x1_ASAP7_75t_L g1752 ( 
.A(n_1742),
.B(n_1700),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1748),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1750),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1741),
.A2(n_1704),
.B1(n_1700),
.B2(n_1701),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1744),
.A2(n_1704),
.B(n_1701),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1743),
.Y(n_1757)
);

AOI222xp33_ASAP7_75t_L g1758 ( 
.A1(n_1749),
.A2(n_1706),
.B1(n_1697),
.B2(n_1700),
.C1(n_1704),
.C2(n_1615),
.Y(n_1758)
);

XOR2xp5_ASAP7_75t_L g1759 ( 
.A(n_1755),
.B(n_1751),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1752),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1754),
.A2(n_1756),
.B1(n_1745),
.B2(n_1746),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1757),
.B(n_1747),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1753),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1758),
.Y(n_1764)
);

NOR3xp33_ASAP7_75t_L g1765 ( 
.A(n_1757),
.B(n_1706),
.C(n_1697),
.Y(n_1765)
);

OAI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1764),
.A2(n_1704),
.B1(n_1674),
.B2(n_1664),
.Y(n_1766)
);

AOI221x1_ASAP7_75t_SL g1767 ( 
.A1(n_1762),
.A2(n_1618),
.B1(n_1620),
.B2(n_1631),
.C(n_1643),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1760),
.Y(n_1768)
);

O2A1O1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1761),
.A2(n_1615),
.B(n_1614),
.C(n_1619),
.Y(n_1769)
);

NOR2x1_ASAP7_75t_L g1770 ( 
.A(n_1763),
.B(n_1447),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_1770),
.Y(n_1771)
);

NAND4xp75_ASAP7_75t_L g1772 ( 
.A(n_1768),
.B(n_1759),
.C(n_1765),
.D(n_1456),
.Y(n_1772)
);

AOI322xp5_ASAP7_75t_L g1773 ( 
.A1(n_1766),
.A2(n_1767),
.A3(n_1619),
.B1(n_1769),
.B2(n_1618),
.C1(n_1620),
.C2(n_1627),
.Y(n_1773)
);

AND2x2_ASAP7_75t_SL g1774 ( 
.A(n_1772),
.B(n_1460),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1774),
.Y(n_1775)
);

AOI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1771),
.B1(n_1773),
.B2(n_1620),
.C(n_1618),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1775),
.B(n_1418),
.Y(n_1777)
);

AO221x1_ASAP7_75t_L g1778 ( 
.A1(n_1776),
.A2(n_1631),
.B1(n_1627),
.B2(n_1643),
.C(n_1633),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1777),
.Y(n_1779)
);

OAI21xp5_ASAP7_75t_SL g1780 ( 
.A1(n_1779),
.A2(n_1647),
.B(n_1642),
.Y(n_1780)
);

OAI22x1_ASAP7_75t_SL g1781 ( 
.A1(n_1780),
.A2(n_1504),
.B1(n_1778),
.B2(n_1443),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1781),
.A2(n_1643),
.B1(n_1631),
.B2(n_1627),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1782),
.B(n_1647),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1783),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1784),
.A2(n_1623),
.B1(n_1636),
.B2(n_1629),
.Y(n_1785)
);

AOI211xp5_ASAP7_75t_L g1786 ( 
.A1(n_1785),
.A2(n_1424),
.B(n_1645),
.C(n_1644),
.Y(n_1786)
);


endmodule