module real_jpeg_6663_n_17 (n_108, n_8, n_0, n_111, n_2, n_10, n_114, n_9, n_12, n_107, n_6, n_106, n_11, n_14, n_110, n_112, n_7, n_3, n_5, n_4, n_109, n_115, n_1, n_16, n_15, n_13, n_113, n_17);

input n_108;
input n_8;
input n_0;
input n_111;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_107;
input n_6;
input n_106;
input n_11;
input n_14;
input n_110;
input n_112;
input n_7;
input n_3;
input n_5;
input n_4;
input n_109;
input n_115;
input n_1;
input n_16;
input n_15;
input n_13;
input n_113;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_0),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_1),
.B(n_33),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_2),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_2),
.B(n_93),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_3),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_3),
.B(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_5),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_5),
.B(n_80),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_7),
.B(n_44),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_9),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_9),
.B(n_30),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_11),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_11),
.B(n_38),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_12),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_14),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_16),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_16),
.B(n_55),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_26),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_31),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_66),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_22),
.B(n_89),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_49),
.B(n_97),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR4xp25_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.C(n_37),
.D(n_43),
.Y(n_28)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_37),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21x1_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_92),
.B(n_96),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_87),
.B(n_91),
.Y(n_51)
);

AO221x1_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_63),
.B1(n_84),
.B2(n_85),
.C(n_86),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_68),
.B(n_83),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_67),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_79),
.B(n_82),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_74),
.B(n_78),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_90),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

A2O1A1O1Ixp25_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B(n_102),
.C(n_103),
.D(n_104),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_106),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_107),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_108),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_109),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_110),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_111),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_112),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_113),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_114),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_115),
.Y(n_94)
);


endmodule