module fake_netlist_1_12561_n_22 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_22);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_22;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_5), .B(n_7), .Y(n_10) );
OA22x2_ASAP7_75t_L g11 ( .A1(n_3), .A2(n_6), .B1(n_1), .B2(n_4), .Y(n_11) );
INVx5_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
BUFx8_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
AOI21xp5_ASAP7_75t_L g15 ( .A1(n_9), .A2(n_0), .B(n_1), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_15), .B(n_12), .Y(n_16) );
OR2x2_ASAP7_75t_L g17 ( .A(n_14), .B(n_12), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_16), .B(n_12), .Y(n_18) );
O2A1O1Ixp5_ASAP7_75t_SL g19 ( .A1(n_18), .A2(n_10), .B(n_11), .C(n_16), .Y(n_19) );
AOI211x1_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_10), .B(n_11), .C(n_3), .Y(n_20) );
AOI21x1_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_17), .B(n_2), .Y(n_21) );
AOI211xp5_ASAP7_75t_SL g22 ( .A1(n_21), .A2(n_6), .B(n_0), .C(n_2), .Y(n_22) );
endmodule