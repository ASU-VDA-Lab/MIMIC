module real_jpeg_24271_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_150;
wire n_41;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_74;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_1),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_1),
.A2(n_26),
.B1(n_59),
.B2(n_60),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_1),
.A2(n_26),
.B1(n_69),
.B2(n_70),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_4),
.A2(n_10),
.B1(n_28),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_122),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_122),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_4),
.A2(n_69),
.B1(n_70),
.B2(n_122),
.Y(n_242)
);

INVx8_ASAP7_75t_SL g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_6),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_6),
.A2(n_46),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_6),
.B(n_33),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g217 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_110),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_6),
.B(n_70),
.C(n_82),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_6),
.B(n_58),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_6),
.A2(n_67),
.B1(n_236),
.B2(n_242),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_7),
.A2(n_64),
.B1(n_69),
.B2(n_70),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_7),
.A2(n_59),
.B1(n_60),
.B2(n_64),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_52),
.B1(n_69),
.B2(n_70),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_8),
.A2(n_28),
.B1(n_30),
.B2(n_52),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_8),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_44),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_11),
.A2(n_44),
.B1(n_59),
.B2(n_60),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_11),
.A2(n_44),
.B1(n_69),
.B2(n_70),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_12),
.A2(n_69),
.B1(n_70),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_12),
.A2(n_59),
.B1(n_60),
.B2(n_75),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_14),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_14),
.A2(n_69),
.B1(n_70),
.B2(n_86),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_86),
.Y(n_144)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_15),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_150),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_149),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_20),
.B(n_123),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.C(n_105),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_21),
.B(n_92),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_65),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_48),
.B2(n_49),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_24),
.B(n_48),
.C(n_65),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_33),
.B2(n_43),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_25),
.A2(n_31),
.B1(n_33),
.B2(n_121),
.Y(n_120)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_30),
.B(n_110),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_30),
.B(n_35),
.C(n_37),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_31),
.A2(n_43),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_31),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_40),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_32),
.B(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_32),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_161)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_35),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_34),
.A2(n_38),
.B(n_109),
.C(n_111),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g192 ( 
.A(n_34),
.B(n_110),
.CON(n_192),
.SN(n_192)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_35),
.A2(n_57),
.A3(n_60),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_62),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_51),
.B(n_58),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_53),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_53),
.A2(n_118),
.B1(n_143),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_53),
.A2(n_143),
.B1(n_160),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_54),
.B(n_63),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_54),
.A2(n_58),
.B1(n_183),
.B2(n_192),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

AO22x1_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_56),
.B(n_59),
.Y(n_193)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_58),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_60),
.B1(n_82),
.B2(n_84),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_60),
.B(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_80),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_66),
.B(n_80),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_73),
.B(n_76),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_67),
.A2(n_131),
.B(n_133),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_67),
.A2(n_76),
.B(n_133),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_67),
.A2(n_95),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_67),
.A2(n_233),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_77),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_71),
.B1(n_74),
.B2(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_68),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_70),
.B1(n_82),
.B2(n_84),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_69),
.B(n_247),
.Y(n_246)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_85),
.B(n_87),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_91),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_81),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_81),
.B(n_110),
.Y(n_240)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_103),
.B(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_88),
.A2(n_128),
.B(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_88),
.A2(n_102),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_88),
.A2(n_198),
.B(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_88),
.A2(n_102),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_88),
.A2(n_102),
.B1(n_197),
.B2(n_218),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_100),
.B2(n_104),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_104),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_97),
.A2(n_99),
.B(n_115),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_97),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_97),
.B(n_110),
.Y(n_247)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_100),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_105),
.A2(n_106),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_116),
.C(n_120),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_107),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_108),
.A2(n_112),
.B1(n_113),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_109),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_121),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_148),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_134),
.B1(n_146),
.B2(n_147),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_141),
.B2(n_142),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B(n_145),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_184),
.B(n_262),
.C(n_267),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_171),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_171),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_168),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_166),
.B2(n_167),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_154),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_154),
.B(n_167),
.C(n_168),
.Y(n_263)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_174),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_161),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.C(n_177),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_172),
.B(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_175),
.B(n_177),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.C(n_181),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_203),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_257),
.B(n_261),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_212),
.B(n_256),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_199),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_189),
.B(n_199),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.C(n_196),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_195),
.B(n_196),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_207),
.C(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_211),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_251),
.B(n_255),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_229),
.B(n_250),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_221),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_215),
.B(n_221),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_219),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_227),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_226),
.C(n_227),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_228),
.Y(n_234)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_238),
.B(n_249),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_237),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_237),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_244),
.B(n_248),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_241),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_258),
.B(n_259),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);


endmodule