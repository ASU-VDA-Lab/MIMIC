module real_jpeg_19829_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_255;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx13_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_1),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_1),
.A2(n_36),
.B1(n_67),
.B2(n_72),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_1),
.A2(n_36),
.B1(n_54),
.B2(n_55),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_1),
.A2(n_36),
.B1(n_39),
.B2(n_44),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_32),
.B1(n_54),
.B2(n_55),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_2),
.A2(n_32),
.B1(n_39),
.B2(n_44),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_3),
.A2(n_67),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_3),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_73),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_3),
.A2(n_28),
.B1(n_31),
.B2(n_73),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_3),
.A2(n_39),
.B1(n_44),
.B2(n_73),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_4),
.A2(n_67),
.B1(n_72),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_4),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_134),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_4),
.A2(n_39),
.B1(n_44),
.B2(n_134),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_4),
.A2(n_28),
.B1(n_31),
.B2(n_134),
.Y(n_191)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_66),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_7),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_7),
.A2(n_26),
.B(n_124),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_7),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_9),
.A2(n_67),
.B1(n_72),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_9),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_106),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_9),
.A2(n_28),
.B1(n_31),
.B2(n_106),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_9),
.A2(n_39),
.B1(n_44),
.B2(n_106),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_10),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_10),
.A2(n_14),
.B(n_28),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_10),
.A2(n_39),
.B1(n_44),
.B2(n_121),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_10),
.A2(n_27),
.B1(n_191),
.B2(n_192),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_10),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_10),
.B(n_54),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_10),
.A2(n_54),
.B(n_218),
.Y(n_222)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_12),
.A2(n_39),
.B1(n_44),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_12),
.A2(n_28),
.B1(n_31),
.B2(n_47),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_13),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_13),
.A2(n_45),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_13),
.A2(n_28),
.B1(n_31),
.B2(n_45),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_14),
.A2(n_39),
.B(n_40),
.C(n_41),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_39),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_14),
.A2(n_28),
.B1(n_31),
.B2(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_15),
.Y(n_39)
);

HAxp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_137),
.CON(n_16),
.SN(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_19),
.B(n_108),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_77),
.B2(n_78),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_24),
.B(n_37),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_27),
.A2(n_29),
.B(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_27),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_27),
.A2(n_96),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_27),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_27),
.A2(n_177),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_27),
.A2(n_33),
.B(n_179),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_29),
.B(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_29),
.B(n_121),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_31),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_34),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_35),
.A2(n_98),
.B(n_175),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_41),
.B1(n_43),
.B2(n_46),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_38),
.A2(n_46),
.B(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_38),
.A2(n_83),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_38),
.A2(n_41),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_38),
.A2(n_41),
.B1(n_187),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_38),
.A2(n_41),
.B1(n_209),
.B2(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_38),
.A2(n_225),
.B(n_241),
.Y(n_240)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

AOI32xp33_ASAP7_75t_L g217 ( 
.A1(n_39),
.A2(n_52),
.A3(n_55),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_41),
.A2(n_43),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_41),
.B(n_121),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_42),
.A2(n_44),
.B(n_121),
.C(n_183),
.Y(n_182)
);

NAND2xp33_ASAP7_75t_SL g219 ( 
.A(n_44),
.B(n_51),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_62),
.B1(n_63),
.B2(n_76),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_56),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_51),
.B(n_54),
.C(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_61),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_50),
.B(n_101),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_50),
.A2(n_58),
.B1(n_128),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_50),
.A2(n_58),
.B1(n_150),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_50),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_50),
.A2(n_58),
.B1(n_163),
.B2(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_54),
.Y(n_59)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_66),
.Y(n_119)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_55),
.A2(n_69),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_57),
.A2(n_127),
.B(n_129),
.Y(n_126)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_71),
.B(n_74),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_64),
.A2(n_71),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_64),
.A2(n_105),
.B1(n_107),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_65),
.A2(n_70),
.B1(n_120),
.B2(n_133),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_69),
.C(n_70),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

HAxp5_ASAP7_75t_SL g120 ( 
.A(n_67),
.B(n_121),
.CON(n_120),
.SN(n_120)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_86),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_85),
.B(n_147),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_99),
.C(n_103),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_89),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_107),
.B(n_121),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_115),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_109),
.A2(n_113),
.B1(n_114),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_109),
.Y(n_255)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_115),
.A2(n_116),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_126),
.C(n_130),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_122),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_130),
.B1(n_131),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_126),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_167),
.B(n_250),
.C(n_256),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_156),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_139),
.B(n_156),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_152),
.B2(n_155),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_142),
.B(n_143),
.C(n_155),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_151),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_161),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_157),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_165),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_162),
.B(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_164),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_249),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_243),
.B(n_248),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_230),
.B(n_242),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_212),
.B(n_229),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_200),
.B(n_211),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_188),
.B(n_199),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_180),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_180),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_182),
.B(n_184),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_194),
.B(n_198),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_193),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_201),
.B(n_202),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_210),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_208),
.C(n_210),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_214),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_220),
.B1(n_227),
.B2(n_228),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_221),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_226),
.C(n_227),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_231),
.B(n_232),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_238),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_239),
.C(n_240),
.Y(n_244)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_252),
.Y(n_256)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);


endmodule