module fake_jpeg_15851_n_173 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_23),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_5),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_1),
.Y(n_74)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_5),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_81),
.Y(n_96)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_85),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_91),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_64),
.C(n_72),
.Y(n_91)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_95),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_56),
.B1(n_51),
.B2(n_66),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_76),
.B1(n_74),
.B2(n_73),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_61),
.B1(n_67),
.B2(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_59),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_65),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_123),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_113),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_115),
.Y(n_127)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_124),
.B1(n_69),
.B2(n_70),
.Y(n_128)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_120),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_72),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_121),
.B(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_64),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_68),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_49),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_129),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_52),
.B1(n_57),
.B2(n_55),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_59),
.B1(n_70),
.B2(n_53),
.Y(n_130)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_75),
.B1(n_60),
.B2(n_62),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_126),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_141),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_143),
.Y(n_145)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_140),
.A2(n_134),
.B(n_138),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_149),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_131),
.B1(n_122),
.B2(n_132),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_116),
.B1(n_130),
.B2(n_129),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_137),
.B1(n_121),
.B2(n_108),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_103),
.B(n_133),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_146),
.A2(n_142),
.B1(n_137),
.B2(n_132),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_145),
.B1(n_147),
.B2(n_105),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_152),
.B(n_153),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_150),
.B(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_155),
.B(n_151),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_104),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_158),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_154),
.B1(n_28),
.B2(n_31),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_75),
.C(n_20),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_19),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_22),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_17),
.C(n_46),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_16),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_33),
.B(n_45),
.Y(n_166)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_15),
.B(n_43),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_11),
.B(n_41),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_9),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_38),
.B(n_37),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_36),
.A3(n_35),
.B1(n_34),
.B2(n_2),
.C1(n_3),
.C2(n_4),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g173 ( 
.A(n_172),
.Y(n_173)
);


endmodule