module fake_aes_5730_n_470 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_470);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_470;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g69 ( .A(n_52), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_22), .Y(n_70) );
CKINVDCx16_ASAP7_75t_R g71 ( .A(n_23), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_43), .Y(n_72) );
INVxp67_ASAP7_75t_L g73 ( .A(n_47), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_38), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_51), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_33), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_60), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_30), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_32), .Y(n_79) );
INVxp67_ASAP7_75t_L g80 ( .A(n_48), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_29), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_7), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_6), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_42), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_59), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_37), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_39), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_58), .Y(n_88) );
BUFx10_ASAP7_75t_L g89 ( .A(n_53), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_26), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_13), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_64), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_9), .Y(n_93) );
NOR2xp33_ASAP7_75t_L g94 ( .A(n_65), .B(n_61), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_5), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_7), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_68), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_25), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_54), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_4), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_20), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_35), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_71), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_78), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_82), .B(n_0), .Y(n_105) );
OA21x2_ASAP7_75t_L g106 ( .A1(n_72), .A2(n_0), .B(n_1), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_72), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_95), .Y(n_108) );
CKINVDCx8_ASAP7_75t_R g109 ( .A(n_95), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_89), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_74), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_74), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_78), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_102), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_89), .B(n_1), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_75), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_89), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_96), .B(n_2), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_102), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_96), .B(n_2), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_75), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_73), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_80), .Y(n_123) );
AND2x4_ASAP7_75t_L g124 ( .A(n_76), .B(n_3), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_76), .Y(n_125) );
BUFx2_ASAP7_75t_L g126 ( .A(n_108), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_110), .B(n_91), .Y(n_127) );
AO22x2_ASAP7_75t_L g128 ( .A1(n_124), .A2(n_101), .B1(n_77), .B2(n_88), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_116), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_116), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_110), .B(n_87), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_116), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_116), .Y(n_133) );
OAI22xp33_ASAP7_75t_L g134 ( .A1(n_109), .A2(n_83), .B1(n_100), .B2(n_93), .Y(n_134) );
AND2x6_ASAP7_75t_L g135 ( .A(n_124), .B(n_101), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_116), .Y(n_136) );
INVx8_ASAP7_75t_L g137 ( .A(n_110), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_110), .B(n_86), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_110), .B(n_77), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_116), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_122), .B(n_99), .Y(n_142) );
OR2x2_ASAP7_75t_SL g143 ( .A(n_108), .B(n_88), .Y(n_143) );
INVx4_ASAP7_75t_L g144 ( .A(n_124), .Y(n_144) );
AO21x2_ASAP7_75t_L g145 ( .A1(n_105), .A2(n_98), .B(n_97), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_116), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_124), .B(n_69), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_125), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_124), .Y(n_149) );
INVxp67_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_125), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_129), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_149), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_150), .B(n_123), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_139), .B(n_115), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_139), .B(n_115), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_127), .B(n_118), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_149), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_139), .B(n_114), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_139), .B(n_119), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_144), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_129), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_128), .A2(n_120), .B1(n_118), .B2(n_112), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_127), .B(n_118), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_126), .B(n_109), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_143), .A2(n_109), .B1(n_117), .B2(n_113), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_144), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_147), .B(n_103), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_126), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_128), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_147), .A2(n_121), .B(n_112), .C(n_107), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_129), .Y(n_179) );
XOR2xp5_ASAP7_75t_L g180 ( .A(n_128), .B(n_113), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_129), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_137), .Y(n_182) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_147), .B(n_106), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_133), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_137), .B(n_120), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_164), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
INVxp67_ASAP7_75t_SL g188 ( .A(n_176), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_168), .A2(n_128), .B1(n_135), .B2(n_147), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_159), .B(n_135), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_159), .B(n_145), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_155), .A2(n_137), .B(n_131), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_159), .B(n_145), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_168), .A2(n_135), .B1(n_145), .B2(n_134), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_155), .A2(n_137), .B(n_138), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_160), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_182), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_159), .B(n_104), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_170), .B(n_135), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_180), .A2(n_143), .B1(n_107), .B2(n_111), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_161), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_160), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_170), .B(n_135), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_175), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_185), .A2(n_137), .B(n_140), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_169), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_170), .B(n_120), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_182), .Y(n_211) );
NOR2xp67_ASAP7_75t_L g212 ( .A(n_154), .B(n_121), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_154), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_154), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
INVx1_ASAP7_75t_SL g218 ( .A(n_171), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_210), .B(n_170), .Y(n_219) );
OAI221xp5_ASAP7_75t_L g220 ( .A1(n_203), .A2(n_172), .B1(n_156), .B2(n_180), .C(n_163), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_209), .Y(n_221) );
AOI221xp5_ASAP7_75t_L g222 ( .A1(n_203), .A2(n_171), .B1(n_142), .B2(n_162), .C(n_174), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_209), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_213), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_210), .B(n_157), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g226 ( .A1(n_207), .A2(n_117), .B1(n_164), .B2(n_158), .Y(n_226) );
INVx6_ASAP7_75t_L g227 ( .A(n_186), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_192), .B(n_183), .Y(n_228) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_193), .A2(n_111), .B(n_107), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_218), .B(n_177), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_205), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_218), .A2(n_135), .B1(n_173), .B2(n_164), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_189), .A2(n_173), .B1(n_183), .B2(n_105), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_198), .A2(n_208), .B(n_199), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_201), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_189), .A2(n_183), .B1(n_173), .B2(n_121), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_199), .A2(n_173), .B(n_184), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_201), .B(n_121), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_192), .A2(n_121), .B1(n_106), .B2(n_111), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g240 ( .A1(n_188), .A2(n_106), .B1(n_84), .B2(n_111), .Y(n_240) );
CKINVDCx14_ASAP7_75t_R g241 ( .A(n_194), .Y(n_241) );
AOI22xp33_ASAP7_75t_SL g242 ( .A1(n_194), .A2(n_106), .B1(n_107), .B2(n_81), .Y(n_242) );
NAND2x1p5_ASAP7_75t_L g243 ( .A(n_186), .B(n_106), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_225), .B(n_213), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_228), .B(n_196), .Y(n_245) );
OAI211xp5_ASAP7_75t_L g246 ( .A1(n_226), .A2(n_196), .B(n_202), .C(n_212), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_231), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_231), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_228), .B(n_205), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_241), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_220), .A2(n_205), .B1(n_202), .B2(n_191), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_229), .A2(n_234), .B(n_243), .Y(n_252) );
OAI22xp5_ASAP7_75t_SL g253 ( .A1(n_241), .A2(n_235), .B1(n_242), .B2(n_238), .Y(n_253) );
AOI22xp5_ASAP7_75t_SL g254 ( .A1(n_236), .A2(n_106), .B1(n_200), .B2(n_211), .Y(n_254) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_229), .A2(n_212), .B(n_92), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_222), .A2(n_190), .B1(n_206), .B2(n_195), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_221), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_225), .B(n_187), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_219), .B(n_215), .Y(n_259) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_233), .A2(n_200), .B1(n_211), .B2(n_197), .Y(n_260) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_243), .A2(n_187), .B(n_191), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_223), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_224), .B(n_187), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_230), .A2(n_197), .B1(n_191), .B2(n_204), .Y(n_264) );
OAI211xp5_ASAP7_75t_L g265 ( .A1(n_246), .A2(n_239), .B(n_240), .C(n_232), .Y(n_265) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_252), .A2(n_237), .B(n_70), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_248), .Y(n_267) );
NOR4xp25_ASAP7_75t_SL g268 ( .A(n_248), .B(n_90), .C(n_85), .D(n_79), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_247), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_249), .B(n_243), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_253), .A2(n_227), .B1(n_125), .B2(n_197), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_257), .Y(n_272) );
AOI33xp33_ASAP7_75t_L g273 ( .A1(n_251), .A2(n_141), .A3(n_130), .B1(n_136), .B2(n_140), .B3(n_151), .Y(n_273) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_252), .A2(n_261), .B(n_264), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_249), .B(n_204), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_261), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_247), .Y(n_277) );
OAI211xp5_ASAP7_75t_L g278 ( .A1(n_246), .A2(n_94), .B(n_215), .C(n_216), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_261), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_252), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_245), .B(n_214), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_253), .A2(n_227), .B1(n_125), .B2(n_204), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_249), .B(n_214), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_257), .B(n_214), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_245), .A2(n_227), .B1(n_125), .B2(n_217), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_247), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_272), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g288 ( .A1(n_271), .A2(n_259), .B1(n_251), .B2(n_260), .C(n_244), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_270), .B(n_245), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_270), .B(n_257), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_277), .Y(n_291) );
OAI31xp33_ASAP7_75t_L g292 ( .A1(n_278), .A2(n_260), .A3(n_250), .B(n_258), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_270), .B(n_262), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_275), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_275), .B(n_258), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_277), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_269), .B(n_262), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_276), .B(n_255), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_277), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_272), .B(n_250), .Y(n_300) );
AOI221x1_ASAP7_75t_L g301 ( .A1(n_284), .A2(n_262), .B1(n_263), .B2(n_244), .C(n_254), .Y(n_301) );
INVxp67_ASAP7_75t_L g302 ( .A(n_275), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_267), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_267), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_286), .B(n_258), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_286), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_286), .B(n_263), .Y(n_307) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_276), .B(n_254), .Y(n_308) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_271), .B(n_264), .C(n_125), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_284), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_276), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_279), .Y(n_312) );
AOI32xp33_ASAP7_75t_L g313 ( .A1(n_282), .A2(n_256), .A3(n_4), .B1(n_5), .B2(n_6), .Y(n_313) );
CKINVDCx16_ASAP7_75t_R g314 ( .A(n_281), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_279), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_281), .B(n_255), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_314), .B(n_281), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_290), .B(n_279), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_291), .Y(n_319) );
OR2x6_ASAP7_75t_L g320 ( .A(n_308), .B(n_280), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_290), .B(n_280), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_314), .B(n_283), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_294), .B(n_282), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_300), .B(n_285), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_300), .B(n_302), .Y(n_325) );
NOR3xp33_ASAP7_75t_SL g326 ( .A(n_292), .B(n_278), .C(n_265), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_293), .B(n_280), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_292), .A2(n_285), .B1(n_255), .B2(n_266), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_303), .B(n_265), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_297), .Y(n_330) );
CKINVDCx16_ASAP7_75t_R g331 ( .A(n_293), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_289), .B(n_266), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_297), .B(n_273), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_288), .A2(n_255), .B1(n_227), .B2(n_266), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_289), .B(n_266), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_291), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_303), .B(n_304), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_304), .B(n_305), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_287), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_287), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_310), .Y(n_341) );
AND2x4_ASAP7_75t_SL g342 ( .A(n_307), .B(n_217), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_295), .B(n_274), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_307), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_296), .B(n_274), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_316), .B(n_268), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_316), .B(n_3), .Y(n_347) );
AOI33xp33_ASAP7_75t_L g348 ( .A1(n_311), .A2(n_268), .A3(n_9), .B1(n_10), .B2(n_11), .B3(n_12), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_309), .A2(n_125), .B1(n_216), .B2(n_217), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_299), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_309), .B(n_8), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_299), .Y(n_352) );
NAND2xp33_ASAP7_75t_R g353 ( .A(n_312), .B(n_315), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_299), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_312), .B(n_8), .Y(n_355) );
NAND2xp33_ASAP7_75t_SL g356 ( .A(n_315), .B(n_186), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_331), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_344), .Y(n_358) );
OAI322xp33_ASAP7_75t_L g359 ( .A1(n_347), .A2(n_311), .A3(n_308), .B1(n_125), .B2(n_315), .C1(n_306), .C2(n_313), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_318), .B(n_298), .Y(n_360) );
AOI22xp33_ASAP7_75t_SL g361 ( .A1(n_347), .A2(n_298), .B1(n_315), .B2(n_306), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g362 ( .A1(n_348), .A2(n_313), .B(n_298), .C(n_306), .Y(n_362) );
AOI21xp33_ASAP7_75t_L g363 ( .A1(n_329), .A2(n_298), .B(n_11), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_321), .B(n_10), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_339), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_351), .A2(n_301), .B1(n_186), .B2(n_195), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_340), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_341), .Y(n_368) );
INVxp67_ASAP7_75t_SL g369 ( .A(n_336), .Y(n_369) );
AOI21xp33_ASAP7_75t_L g370 ( .A1(n_346), .A2(n_12), .B(n_13), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_337), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_351), .A2(n_195), .B1(n_132), .B2(n_141), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_326), .A2(n_130), .B1(n_136), .B2(n_146), .C(n_151), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_319), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_342), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_337), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_325), .Y(n_377) );
XNOR2xp5_ASAP7_75t_L g378 ( .A(n_322), .B(n_14), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_321), .B(n_14), .Y(n_379) );
NOR4xp75_ASAP7_75t_L g380 ( .A(n_355), .B(n_15), .C(n_16), .D(n_17), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_324), .A2(n_333), .B1(n_323), .B2(n_328), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_356), .A2(n_166), .B(n_181), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_338), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_330), .B(n_15), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_327), .B(n_16), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_319), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_332), .B(n_17), .Y(n_387) );
INVx1_ASAP7_75t_SL g388 ( .A(n_317), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_350), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_328), .A2(n_132), .B1(n_133), .B2(n_148), .Y(n_390) );
OAI33xp33_ASAP7_75t_L g391 ( .A1(n_343), .A2(n_148), .A3(n_19), .B1(n_21), .B2(n_24), .B3(n_27), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_352), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_354), .Y(n_393) );
NAND2x1_ASAP7_75t_L g394 ( .A(n_320), .B(n_132), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_335), .B(n_18), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_349), .A2(n_132), .B1(n_31), .B2(n_34), .Y(n_396) );
NOR3xp33_ASAP7_75t_L g397 ( .A(n_348), .B(n_28), .C(n_36), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_357), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_365), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_378), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_368), .B(n_334), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_367), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_381), .B(n_345), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_394), .Y(n_404) );
OAI32xp33_ASAP7_75t_L g405 ( .A1(n_358), .A2(n_353), .A3(n_356), .B1(n_349), .B2(n_345), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_388), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_371), .B(n_320), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_368), .Y(n_408) );
XOR2x2_ASAP7_75t_L g409 ( .A(n_380), .B(n_353), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_376), .B(n_40), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_369), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_383), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_377), .B(n_41), .Y(n_413) );
INVx2_ASAP7_75t_SL g414 ( .A(n_375), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_360), .B(n_44), .Y(n_415) );
NAND4xp25_ASAP7_75t_SL g416 ( .A(n_397), .B(n_45), .C(n_46), .D(n_49), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_369), .B(n_50), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_374), .Y(n_418) );
NOR3xp33_ASAP7_75t_SL g419 ( .A(n_359), .B(n_55), .C(n_56), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_392), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_364), .B(n_57), .Y(n_421) );
NOR3xp33_ASAP7_75t_SL g422 ( .A(n_363), .B(n_62), .C(n_63), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_393), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_379), .B(n_66), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_384), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_389), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_387), .B(n_67), .Y(n_427) );
NAND2xp33_ASAP7_75t_L g428 ( .A(n_362), .B(n_152), .Y(n_428) );
INVxp67_ASAP7_75t_L g429 ( .A(n_408), .Y(n_429) );
OAI221xp5_ASAP7_75t_SL g430 ( .A1(n_406), .A2(n_385), .B1(n_361), .B2(n_362), .C(n_390), .Y(n_430) );
NAND4xp75_ASAP7_75t_L g431 ( .A(n_419), .B(n_370), .C(n_382), .D(n_395), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g432 ( .A(n_428), .B(n_419), .C(n_401), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_403), .B(n_361), .Y(n_433) );
XOR2xp5_ASAP7_75t_L g434 ( .A(n_398), .B(n_372), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_404), .B(n_386), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_401), .A2(n_391), .B1(n_366), .B2(n_373), .C(n_396), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_409), .A2(n_152), .B1(n_166), .B2(n_167), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_426), .Y(n_438) );
OAI21xp33_ASAP7_75t_SL g439 ( .A1(n_404), .A2(n_167), .B(n_178), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_420), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_405), .A2(n_167), .B1(n_178), .B2(n_179), .C(n_181), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_423), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_418), .Y(n_443) );
XNOR2xp5_ASAP7_75t_L g444 ( .A(n_400), .B(n_178), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_399), .Y(n_445) );
NOR2xp33_ASAP7_75t_R g446 ( .A(n_444), .B(n_400), .Y(n_446) );
OAI211xp5_ASAP7_75t_L g447 ( .A1(n_430), .A2(n_411), .B(n_414), .C(n_407), .Y(n_447) );
NAND4xp25_ASAP7_75t_L g448 ( .A(n_432), .B(n_424), .C(n_421), .D(n_427), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_434), .Y(n_449) );
OAI21xp33_ASAP7_75t_SL g450 ( .A1(n_429), .A2(n_418), .B(n_425), .Y(n_450) );
AOI221xp5_ASAP7_75t_SL g451 ( .A1(n_433), .A2(n_402), .B1(n_413), .B2(n_415), .C(n_417), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_431), .A2(n_416), .B1(n_422), .B2(n_410), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_436), .A2(n_179), .B1(n_181), .B2(n_441), .Y(n_453) );
AOI322xp5_ASAP7_75t_L g454 ( .A1(n_440), .A2(n_445), .A3(n_442), .B1(n_438), .B2(n_435), .C1(n_439), .C2(n_437), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_443), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_430), .A2(n_433), .B1(n_429), .B2(n_401), .C(n_412), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_443), .Y(n_457) );
OAI22xp33_ASAP7_75t_L g458 ( .A1(n_432), .A2(n_331), .B1(n_357), .B2(n_433), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_456), .A2(n_447), .B1(n_458), .B2(n_449), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_446), .Y(n_460) );
NAND5xp2_ASAP7_75t_L g461 ( .A(n_453), .B(n_452), .C(n_451), .D(n_454), .E(n_455), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_457), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_460), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_462), .Y(n_464) );
XNOR2xp5_ASAP7_75t_L g465 ( .A(n_459), .B(n_448), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_464), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_463), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_466), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_468), .A2(n_467), .B1(n_465), .B2(n_450), .Y(n_469) );
NAND2x2_ASAP7_75t_L g470 ( .A(n_469), .B(n_461), .Y(n_470) );
endmodule