module fake_jpeg_24068_n_257 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_39),
.CON(n_55),
.SN(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_45),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_2),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_3),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_35),
.Y(n_53)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_51),
.B1(n_68),
.B2(n_17),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_34),
.B1(n_23),
.B2(n_33),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_65),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_34),
.B1(n_31),
.B2(n_23),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_36),
.B1(n_42),
.B2(n_23),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_31),
.B1(n_22),
.B2(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_19),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_73),
.B(n_76),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_47),
.B(n_25),
.Y(n_76)
);

AOI32xp33_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_42),
.A3(n_45),
.B1(n_36),
.B2(n_46),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_79),
.A2(n_88),
.B1(n_106),
.B2(n_105),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_35),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_45),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_46),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_103),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_21),
.B1(n_18),
.B2(n_72),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_50),
.B(n_27),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_32),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_69),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_58),
.B(n_17),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_26),
.B1(n_20),
.B2(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_58),
.B(n_29),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_105),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_36),
.B1(n_18),
.B2(n_29),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_26),
.B1(n_20),
.B2(n_32),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_3),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_67),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_72),
.A2(n_36),
.B1(n_28),
.B2(n_21),
.Y(n_106)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_111),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_131),
.B1(n_101),
.B2(n_94),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_110),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_85),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_52),
.B1(n_48),
.B2(n_64),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_95),
.B1(n_78),
.B2(n_75),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_132),
.B1(n_83),
.B2(n_77),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_15),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_121),
.Y(n_142)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_32),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_4),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_126),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_67),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_103),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_32),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_43),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_32),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_129),
.B(n_104),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_135),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_109),
.B1(n_122),
.B2(n_129),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_141),
.B1(n_150),
.B2(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_90),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_148),
.C(n_153),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_159),
.Y(n_166)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_152),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_92),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_99),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_99),
.B1(n_104),
.B2(n_78),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_103),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_92),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_43),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_119),
.C(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_75),
.Y(n_160)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_135),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_162),
.B(n_150),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_172),
.C(n_173),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_124),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_174),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_116),
.Y(n_171)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_124),
.C(n_114),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_119),
.C(n_128),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_158),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_133),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_147),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_116),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_128),
.B1(n_116),
.B2(n_132),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_183),
.A3(n_149),
.B1(n_146),
.B2(n_142),
.C1(n_144),
.C2(n_134),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_117),
.C(n_43),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_141),
.C(n_134),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_136),
.A2(n_102),
.B1(n_82),
.B2(n_108),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_177),
.B1(n_171),
.B2(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_182),
.B1(n_161),
.B2(n_163),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_188),
.A2(n_201),
.B(n_202),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_179),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_196),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_140),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_195),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_173),
.C(n_169),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_164),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_149),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_198),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_180),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_175),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_199),
.B(n_5),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_63),
.A3(n_61),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_149),
.B(n_157),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_154),
.B(n_26),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_206),
.C(n_216),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_174),
.C(n_170),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_212),
.B1(n_214),
.B2(n_185),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_181),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_211),
.B(n_202),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_102),
.B1(n_77),
.B2(n_93),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_187),
.A2(n_192),
.B1(n_195),
.B2(n_191),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_213),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_49),
.B1(n_26),
.B2(n_20),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_4),
.C(n_5),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_5),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_222),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_194),
.B1(n_186),
.B2(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_220),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_208),
.A2(n_198),
.B(n_186),
.Y(n_220)
);

FAx1_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_190),
.CI(n_213),
.CON(n_221),
.SN(n_221)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_227),
.B(n_216),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_201),
.B1(n_193),
.B2(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

INVx11_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_197),
.B(n_7),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_6),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_229),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_210),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_232),
.C(n_238),
.Y(n_244)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_204),
.C(n_209),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_9),
.C(n_10),
.Y(n_238)
);

AOI31xp67_ASAP7_75t_SL g240 ( 
.A1(n_231),
.A2(n_227),
.A3(n_221),
.B(n_223),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_242),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_221),
.B(n_223),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_241),
.A2(n_243),
.B(n_237),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_228),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_10),
.B(n_11),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_233),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_248),
.B(n_249),
.Y(n_250)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_244),
.B(n_232),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_234),
.C(n_235),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_234),
.B(n_238),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_10),
.C(n_11),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_247),
.A2(n_230),
.B(n_235),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_11),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_253),
.B(n_254),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_250),
.B(n_13),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_14),
.Y(n_257)
);


endmodule