module fake_jpeg_15737_n_12 (n_3, n_2, n_1, n_0, n_4, n_12);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_12;

wire n_11;
wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

INVx5_ASAP7_75t_L g5 ( 
.A(n_4),
.Y(n_5)
);

BUFx12_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

OAI21xp33_ASAP7_75t_L g7 ( 
.A1(n_6),
.A2(n_0),
.B(n_1),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_8),
.B(n_6),
.Y(n_9)
);

OAI21xp33_ASAP7_75t_L g10 ( 
.A1(n_9),
.A2(n_8),
.B(n_0),
.Y(n_10)
);

AOI322xp5_ASAP7_75t_L g11 ( 
.A1(n_10),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_0),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_2),
.C(n_5),
.Y(n_12)
);


endmodule