module fake_jpeg_9566_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_31),
.Y(n_39)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_32),
.Y(n_48)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_38),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_26),
.C(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.C(n_26),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_28),
.B1(n_19),
.B2(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_24),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_19),
.B1(n_17),
.B2(n_26),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_19),
.B1(n_17),
.B2(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_15),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_53),
.B1(n_62),
.B2(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_51),
.B(n_54),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_30),
.B(n_31),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_48),
.B(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_38),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_61),
.Y(n_64)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_28),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_16),
.B1(n_33),
.B2(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_46),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_25),
.B(n_36),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_71),
.B1(n_36),
.B2(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_70),
.Y(n_82)
);

INVxp67_ASAP7_75t_SL g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_41),
.B1(n_29),
.B2(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_74),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_25),
.B1(n_16),
.B2(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_76),
.Y(n_81)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_60),
.B(n_20),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_87),
.B(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_85),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_59),
.B1(n_13),
.B2(n_14),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_49),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_1),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_68),
.C(n_70),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_90),
.C(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_91),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_0),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_87),
.B1(n_89),
.B2(n_82),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_100),
.C(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_71),
.C(n_78),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_23),
.A3(n_21),
.B1(n_16),
.B2(n_9),
.C1(n_12),
.C2(n_11),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_102),
.B(n_1),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_104),
.B1(n_102),
.B2(n_95),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_108),
.C(n_110),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_86),
.C(n_83),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_23),
.B1(n_21),
.B2(n_3),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_12),
.B1(n_3),
.B2(n_4),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_109),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_105),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_121),
.C(n_114),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

OAI21x1_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_110),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_2),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_127),
.C(n_128),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_125),
.B(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_2),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_129),
.A2(n_5),
.B(n_6),
.Y(n_133)
);

NOR2xp67_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_122),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_133),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_132),
.B(n_126),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_135),
.Y(n_137)
);


endmodule