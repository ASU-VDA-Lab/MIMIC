module fake_jpeg_19758_n_174 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_36),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_13),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_43),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_31),
.B1(n_16),
.B2(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_48),
.A2(n_62),
.B1(n_1),
.B2(n_2),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_57),
.B1(n_60),
.B2(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_68),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_18),
.B1(n_29),
.B2(n_27),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_18),
.B1(n_27),
.B2(n_23),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_16),
.B1(n_30),
.B2(n_20),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_21),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_77),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_41),
.B1(n_21),
.B2(n_34),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_78),
.B1(n_86),
.B2(n_56),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_79),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_82),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_35),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_20),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_28),
.B1(n_24),
.B2(n_21),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_28),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_17),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_34),
.C(n_35),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_88),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_65),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_54),
.A2(n_34),
.B1(n_17),
.B2(n_2),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_17),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_0),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_51),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_51),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_101),
.Y(n_113)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_74),
.B1(n_90),
.B2(n_91),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_96),
.B1(n_102),
.B2(n_83),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_58),
.B1(n_54),
.B2(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_66),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_58),
.B1(n_67),
.B2(n_56),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_107),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_117),
.Y(n_126)
);

AOI22x1_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_84),
.B1(n_79),
.B2(n_89),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_121),
.B(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_122),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_81),
.C(n_80),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_120),
.C(n_97),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_92),
.C(n_101),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_92),
.B(n_102),
.C(n_109),
.D(n_97),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_89),
.B(n_86),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_98),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_114),
.A2(n_94),
.B1(n_108),
.B2(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_120),
.B(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_132),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_138),
.B1(n_125),
.B2(n_111),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_100),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_117),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_100),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_104),
.A3(n_70),
.B1(n_77),
.B2(n_108),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_121),
.B(n_125),
.C(n_124),
.D(n_114),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_108),
.B1(n_73),
.B2(n_65),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_131),
.C(n_119),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_128),
.B1(n_137),
.B2(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_112),
.B1(n_114),
.B2(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_133),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_151),
.B1(n_156),
.B2(n_144),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_153),
.A2(n_155),
.B(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_148),
.B(n_71),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_146),
.B(n_140),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_70),
.A3(n_14),
.B1(n_11),
.B2(n_65),
.C1(n_8),
.C2(n_2),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_139),
.C(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_158),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_160),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_169),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_SL g168 ( 
.A(n_166),
.B(n_153),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_164),
.B(n_11),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g169 ( 
.A1(n_163),
.A2(n_156),
.B(n_158),
.C(n_161),
.D(n_6),
.Y(n_169)
);

AOI31xp33_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_14),
.A3(n_8),
.B(n_10),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_170),
.B(n_10),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_10),
.Y(n_174)
);


endmodule