module real_jpeg_16999_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_4),
.B(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_4),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_4),
.B(n_60),
.Y(n_59)
);

AND2x4_ASAP7_75t_SL g63 ( 
.A(n_4),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_4),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_4),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_4),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_4),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_5),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_5),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_7),
.Y(n_159)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_7),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_8),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_47),
.Y(n_46)
);

AND2x4_ASAP7_75t_SL g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_8),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_8),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_8),
.B(n_28),
.Y(n_104)
);

NAND2x1p5_ASAP7_75t_L g124 ( 
.A(n_8),
.B(n_125),
.Y(n_124)
);

NAND2x1_ASAP7_75t_L g167 ( 
.A(n_8),
.B(n_168),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_9),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_10),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_10),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_10),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_10),
.B(n_196),
.Y(n_195)
);

BUFx8_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_11),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_180),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_144),
.B(n_179),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_113),
.B(n_143),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_85),
.B(n_112),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_50),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_18),
.B(n_50),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_35),
.C(n_43),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_23),
.B1(n_33),
.B2(n_34),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_20),
.A2(n_33),
.B1(n_132),
.B2(n_136),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_20),
.A2(n_95),
.B(n_104),
.C(n_133),
.Y(n_151)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_24),
.A2(n_25),
.B1(n_119),
.B2(n_128),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_29),
.C(n_33),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_41),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_26),
.B(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_30),
.B(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_32),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_35),
.A2(n_43),
.B1(n_44),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_35),
.A2(n_36),
.B(n_39),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_39),
.A2(n_40),
.B1(n_54),
.B2(n_55),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_39),
.A2(n_40),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_55),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_46),
.B(n_91),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_47),
.Y(n_172)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_69),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_70),
.C(n_84),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_62),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_53),
.A2(n_101),
.B(n_105),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_53),
.A2(n_63),
.B(n_68),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_63),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_88),
.B(n_90),
.C(n_95),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_88),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_63),
.A2(n_67),
.B1(n_88),
.B2(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_66),
.B(n_119),
.C(n_124),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_83),
.B2(n_84),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_82),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_72),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_72),
.B(n_76),
.C(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_78),
.Y(n_176)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_79),
.A2(n_140),
.B1(n_155),
.B2(n_161),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_99),
.B(n_111),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_96),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_88),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_88),
.B(n_103),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_88),
.B(n_104),
.C(n_167),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_88),
.A2(n_109),
.B1(n_193),
.B2(n_199),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_91),
.A2(n_93),
.B1(n_156),
.B2(n_160),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_91),
.B(n_140),
.C(n_156),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_107),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_106),
.B(n_110),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_103),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_104),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_115),
.Y(n_143)
);

XOR2x2_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_130),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_129),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_129),
.C(n_130),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_123),
.B1(n_124),
.B2(n_128),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

OR2x6_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_138),
.C(n_142),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_146),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_162),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_149),
.C(n_162),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_154),
.C(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_178),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_164),
.B(n_170),
.C(n_178),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_169),
.Y(n_164)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_173),
.B(n_177),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_173),
.Y(n_177)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_219),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_184),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_202),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_200),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_192),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_218),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_214),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);


endmodule