module fake_netlist_5_2359_n_70 (n_8, n_10, n_4, n_5, n_7, n_0, n_12, n_9, n_14, n_2, n_16, n_13, n_3, n_11, n_17, n_15, n_6, n_1, n_70);

input n_8;
input n_10;
input n_4;
input n_5;
input n_7;
input n_0;
input n_12;
input n_9;
input n_14;
input n_2;
input n_16;
input n_13;
input n_3;
input n_11;
input n_17;
input n_15;
input n_6;
input n_1;

output n_70;

wire n_54;
wire n_29;
wire n_43;
wire n_47;
wire n_58;
wire n_67;
wire n_69;
wire n_36;
wire n_25;
wire n_53;
wire n_18;
wire n_27;
wire n_42;
wire n_64;
wire n_22;
wire n_45;
wire n_24;
wire n_46;
wire n_28;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_38;
wire n_61;
wire n_68;
wire n_35;
wire n_32;
wire n_41;
wire n_65;
wire n_56;
wire n_51;
wire n_63;
wire n_19;
wire n_57;
wire n_37;
wire n_59;
wire n_26;
wire n_30;
wire n_33;
wire n_55;
wire n_48;
wire n_31;
wire n_23;
wire n_50;
wire n_66;
wire n_49;
wire n_52;
wire n_60;
wire n_20;
wire n_39;

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_3),
.Y(n_18)
);

OA21x2_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_7),
.B(n_10),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_4),
.B1(n_1),
.B2(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_5),
.B(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2x1_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_21),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_20),
.B(n_30),
.Y(n_37)
);

OAI21x1_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_22),
.B(n_19),
.Y(n_38)
);

AOI21x1_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_18),
.B(n_23),
.Y(n_39)
);

OAI21x1_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_19),
.B(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2x1_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_19),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_37),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_49),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_48),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_50),
.B1(n_44),
.B2(n_31),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_54),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_55),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_22),
.B(n_26),
.C(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_63),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

OAI21x1_ASAP7_75t_SL g67 ( 
.A1(n_64),
.A2(n_60),
.B(n_28),
.Y(n_67)
);

AOI221xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_29),
.B1(n_27),
.B2(n_58),
.C(n_60),
.Y(n_68)
);

XNOR2x1_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_66),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g70 ( 
.A(n_69),
.Y(n_70)
);


endmodule