module fake_jpeg_24360_n_206 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_15),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_33),
.Y(n_55)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_27),
.B1(n_26),
.B2(n_21),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_51),
.B1(n_25),
.B2(n_18),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_27),
.B1(n_21),
.B2(n_22),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_27),
.B1(n_21),
.B2(n_22),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_15),
.C(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_23),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_61),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_36),
.B1(n_32),
.B2(n_34),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_18),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_22),
.B1(n_20),
.B2(n_14),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_69),
.B1(n_18),
.B2(n_14),
.Y(n_80)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_44),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_81),
.Y(n_92)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_76),
.Y(n_100)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_55),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_53),
.B1(n_50),
.B2(n_45),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_58),
.B1(n_46),
.B2(n_43),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_36),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_60),
.C(n_24),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_14),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_107),
.B1(n_88),
.B2(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_74),
.B(n_57),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_101),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_62),
.B(n_36),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_91),
.B(n_83),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_105),
.C(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_62),
.C(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_78),
.B(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_43),
.C(n_41),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_94),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_86),
.C(n_78),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_92),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_86),
.B(n_85),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_116),
.B(n_121),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_114),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_77),
.B(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_17),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_97),
.B(n_109),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_124),
.B1(n_126),
.B2(n_125),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_83),
.B1(n_87),
.B2(n_43),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_41),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_87),
.B1(n_46),
.B2(n_41),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_128),
.A2(n_123),
.B1(n_116),
.B2(n_127),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_75),
.Y(n_130)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_105),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_137),
.C(n_142),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_139),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_144),
.B1(n_17),
.B2(n_16),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_136),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_112),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_24),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_143),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_24),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_24),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_17),
.B1(n_24),
.B2(n_13),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_121),
.A3(n_111),
.B1(n_137),
.B2(n_131),
.C1(n_113),
.C2(n_142),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_16),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_138),
.A2(n_124),
.B(n_119),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_R g163 ( 
.A(n_146),
.B(n_16),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_151),
.A2(n_154),
.B1(n_155),
.B2(n_158),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_0),
.B(n_1),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_134),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_149),
.A2(n_141),
.B(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_162),
.Y(n_173)
);

AO21x1_ASAP7_75t_SL g160 ( 
.A1(n_156),
.A2(n_16),
.B(n_3),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_150),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_16),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_168),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_148),
.B(n_11),
.Y(n_162)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_11),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_157),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_155),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_1),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_10),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_174),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_179),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_157),
.C(n_151),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_168),
.C(n_170),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_173),
.A2(n_161),
.B1(n_152),
.B2(n_6),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_184),
.B(n_175),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_171),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_6),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_188),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_172),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_190),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_187),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_181),
.A2(n_7),
.B(n_8),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_194),
.B(n_185),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_SL g195 ( 
.A(n_193),
.B(n_183),
.Y(n_195)
);

OAI21x1_ASAP7_75t_SL g201 ( 
.A1(n_195),
.A2(n_7),
.B(n_8),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_197),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_189),
.B(n_191),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_198),
.A2(n_199),
.B(n_7),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_SL g205 ( 
.A(n_204),
.B(n_202),
.C(n_203),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_SL g206 ( 
.A(n_205),
.B(n_8),
.Y(n_206)
);


endmodule