module fake_ariane_2007_n_1751 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1751);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1751;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_263;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_114),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_64),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_35),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_11),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_25),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_25),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_117),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_10),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_81),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

BUFx8_ASAP7_75t_SL g172 ( 
.A(n_150),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_48),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_127),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_17),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_126),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_141),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_17),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_53),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_46),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_93),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_145),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_129),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_155),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_132),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_49),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_121),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_72),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_54),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_120),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_21),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_75),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_62),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_66),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_74),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_77),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_29),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_37),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_88),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_103),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_105),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_3),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_57),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_148),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_29),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_106),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_19),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_34),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_31),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_28),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_69),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_99),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_45),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_86),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_10),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_13),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_20),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_115),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_133),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_65),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_2),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_123),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_112),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_104),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_21),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_3),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_142),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_109),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_34),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_71),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_9),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_18),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_92),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_134),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_90),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_55),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_84),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_78),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_48),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_50),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_52),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_41),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_42),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_91),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_139),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_76),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_0),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_18),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_50),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_96),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_54),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_124),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_47),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_102),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_119),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_144),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_45),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_38),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_70),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_67),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_94),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_131),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_108),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_116),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_46),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_107),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_60),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_137),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_49),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_130),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_16),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_27),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_153),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_39),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_38),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_89),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_110),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_101),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_37),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_51),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_61),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_51),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_63),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_16),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_27),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_5),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_32),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_151),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_2),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_55),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_138),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_95),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_125),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_32),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_85),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_211),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_172),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_196),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_297),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_187),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_266),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_211),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_211),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_266),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_192),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_211),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_187),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_212),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_211),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_211),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_207),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_220),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_165),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_212),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_211),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_162),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_211),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_161),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_298),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_249),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_254),
.B(n_0),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_167),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_211),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_173),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_278),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_156),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_156),
.B(n_1),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_192),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_170),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_170),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_171),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_171),
.B(n_1),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_198),
.B(n_4),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_198),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_199),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_283),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_199),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_175),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_203),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_203),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_178),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_R g351 ( 
.A(n_157),
.B(n_98),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_190),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_276),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_254),
.B(n_4),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_218),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_218),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_223),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_206),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_223),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_209),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_276),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_227),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_276),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_276),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_168),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_214),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_301),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_217),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_301),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_219),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_227),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_228),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_256),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_228),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_221),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_301),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_229),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_224),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_319),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_316),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_305),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_319),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_305),
.Y(n_384)
);

AND2x2_ASAP7_75t_SL g385 ( 
.A(n_341),
.B(n_191),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_311),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_335),
.B(n_229),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_335),
.B(n_256),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_338),
.B(n_239),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_365),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_318),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_310),
.B(n_239),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_324),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_326),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_338),
.B(n_260),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_339),
.B(n_260),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_326),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_309),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_339),
.B(n_268),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_340),
.B(n_243),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_340),
.B(n_243),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_343),
.B(n_301),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_337),
.B(n_314),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_344),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_346),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_348),
.B(n_251),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_348),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_349),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_317),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_349),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_355),
.B(n_162),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_355),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_356),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_356),
.B(n_357),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_357),
.B(n_251),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_359),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_359),
.B(n_180),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_323),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_362),
.B(n_252),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_371),
.B(n_252),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_371),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_313),
.B(n_263),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_372),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_372),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_374),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_337),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_377),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_377),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_341),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_336),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_373),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_325),
.B(n_263),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_396),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_361),
.Y(n_452)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_410),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_428),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

OR2x6_ASAP7_75t_L g457 ( 
.A(n_415),
.B(n_373),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_396),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_396),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_385),
.B(n_342),
.C(n_351),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_327),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_415),
.B(n_331),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_383),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_383),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_416),
.B(n_307),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_333),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_381),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_415),
.B(n_347),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_447),
.B(n_350),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_381),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_391),
.Y(n_472)
);

BUFx4f_ASAP7_75t_L g473 ( 
.A(n_447),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_428),
.Y(n_474)
);

OR2x6_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_330),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_352),
.Y(n_476)
);

BUFx6f_ASAP7_75t_SL g477 ( 
.A(n_385),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_380),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_403),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_360),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_447),
.B(n_366),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_450),
.B(n_330),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_428),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_380),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_447),
.B(n_368),
.Y(n_486)
);

INVxp33_ASAP7_75t_SL g487 ( 
.A(n_424),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_428),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_445),
.B(n_370),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_385),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_391),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_428),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_385),
.A2(n_322),
.B1(n_328),
.B2(n_354),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_428),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_449),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_438),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_449),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_438),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_391),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_438),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_399),
.A2(n_354),
.B1(n_376),
.B2(n_353),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_426),
.B(n_432),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_398),
.Y(n_503)
);

NAND3xp33_ASAP7_75t_L g504 ( 
.A(n_445),
.B(n_193),
.C(n_264),
.Y(n_504)
);

OAI22xp33_ASAP7_75t_L g505 ( 
.A1(n_434),
.A2(n_164),
.B1(n_245),
.B2(n_179),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_399),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_403),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_398),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_438),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_391),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_408),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_417),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_410),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_398),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_444),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_449),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_391),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_398),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_417),
.Y(n_521)
);

AND2x2_ASAP7_75t_SL g522 ( 
.A(n_426),
.B(n_191),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_391),
.Y(n_523)
);

BUFx4f_ASAP7_75t_L g524 ( 
.A(n_402),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_402),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_416),
.B(n_375),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_417),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_434),
.B(n_378),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_429),
.B(n_215),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_429),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_429),
.B(n_216),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_420),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_391),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_L g535 ( 
.A(n_414),
.B(n_418),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_402),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_420),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_391),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_420),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_390),
.B(n_201),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_420),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_390),
.B(n_201),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_402),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_402),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_440),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_392),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_408),
.B(n_306),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_426),
.B(n_432),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_419),
.B(n_422),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_426),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_433),
.B(n_363),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_440),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_440),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_410),
.Y(n_554)
);

INVx5_ASAP7_75t_L g555 ( 
.A(n_410),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_392),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_440),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_392),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_433),
.B(n_364),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_392),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_392),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_402),
.Y(n_562)
);

AOI21x1_ASAP7_75t_L g563 ( 
.A1(n_382),
.A2(n_267),
.B(n_264),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_433),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_426),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_390),
.B(n_201),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_392),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_424),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_446),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_439),
.B(n_270),
.C(n_267),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_444),
.A2(n_329),
.B1(n_320),
.B2(n_345),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_416),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_446),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_432),
.B(n_180),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_439),
.A2(n_369),
.B1(n_367),
.B2(n_200),
.Y(n_575)
);

AND2x2_ASAP7_75t_SL g576 ( 
.A(n_432),
.B(n_204),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_402),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_392),
.Y(n_578)
);

INVxp33_ASAP7_75t_L g579 ( 
.A(n_406),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_L g580 ( 
.A(n_422),
.B(n_158),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_423),
.B(n_270),
.Y(n_581)
);

BUFx10_ASAP7_75t_L g582 ( 
.A(n_432),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_423),
.B(n_271),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_446),
.Y(n_584)
);

AOI21x1_ASAP7_75t_L g585 ( 
.A1(n_382),
.A2(n_386),
.B(n_384),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_425),
.B(n_308),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_425),
.B(n_435),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_406),
.B(n_201),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_406),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_402),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_405),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_392),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_446),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_405),
.Y(n_594)
);

AO21x2_ASAP7_75t_L g595 ( 
.A1(n_387),
.A2(n_272),
.B(n_271),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_506),
.B(n_384),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_522),
.A2(n_405),
.B1(n_427),
.B2(n_431),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_496),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_461),
.B(n_435),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_564),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_476),
.B(n_522),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_522),
.B(n_441),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_496),
.Y(n_603)
);

INVx8_ASAP7_75t_L g604 ( 
.A(n_457),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_576),
.B(n_441),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_507),
.Y(n_606)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_571),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_576),
.B(n_386),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_500),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_576),
.B(n_442),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_495),
.B(n_442),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_495),
.B(n_443),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_506),
.B(n_443),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_506),
.B(n_388),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_582),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_582),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_582),
.B(n_388),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_582),
.B(n_389),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_460),
.A2(n_490),
.B1(n_477),
.B2(n_457),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_500),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_497),
.B(n_518),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_508),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_512),
.B(n_405),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_497),
.B(n_518),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_512),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_471),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_508),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_502),
.B(n_427),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_L g629 ( 
.A(n_550),
.B(n_389),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_471),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_510),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_550),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_506),
.B(n_528),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_565),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_565),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_477),
.A2(n_405),
.B1(n_431),
.B2(n_436),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_514),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_472),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_462),
.B(n_393),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_502),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_514),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_463),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_502),
.B(n_431),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_548),
.B(n_394),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_468),
.B(n_394),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_520),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_463),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_579),
.B(n_397),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_548),
.B(n_397),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_548),
.B(n_400),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_548),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_572),
.B(n_321),
.Y(n_652)
);

NAND3xp33_ASAP7_75t_L g653 ( 
.A(n_460),
.B(n_401),
.C(n_400),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_586),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_472),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_549),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_530),
.B(n_401),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_572),
.B(n_334),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_472),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_526),
.B(n_387),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_575),
.A2(n_273),
.B1(n_303),
.B2(n_299),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_530),
.B(n_404),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_540),
.B(n_404),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_540),
.B(n_407),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_542),
.B(n_407),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_594),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_542),
.B(n_409),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_566),
.B(n_409),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_566),
.B(n_412),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_564),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_588),
.B(n_395),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_480),
.B(n_489),
.Y(n_672)
);

OAI21xp33_ASAP7_75t_L g673 ( 
.A1(n_493),
.A2(n_411),
.B(n_395),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_490),
.B(n_412),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_473),
.B(n_379),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_526),
.B(n_411),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_457),
.B(n_413),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_472),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_464),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_591),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_588),
.B(n_413),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_457),
.B(n_437),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_467),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_473),
.A2(n_535),
.B(n_452),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_464),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_477),
.A2(n_437),
.B1(n_436),
.B2(n_430),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_529),
.B(n_421),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_591),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_457),
.B(n_430),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_451),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_469),
.B(n_379),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_472),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_479),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_513),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_532),
.B(n_379),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_465),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_568),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_R g698 ( 
.A(n_466),
.B(n_231),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_517),
.B(n_200),
.Y(n_699)
);

BUFx12f_ASAP7_75t_L g700 ( 
.A(n_465),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_574),
.B(n_213),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_521),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_481),
.B(n_379),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_475),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_451),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_574),
.B(n_379),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_574),
.B(n_379),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_475),
.A2(n_272),
.B1(n_275),
.B2(n_292),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_473),
.B(n_275),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_574),
.B(n_213),
.Y(n_710)
);

NOR2xp67_ASAP7_75t_L g711 ( 
.A(n_570),
.B(n_292),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_521),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_SL g713 ( 
.A(n_487),
.B(n_232),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_486),
.B(n_237),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_520),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_475),
.B(n_226),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_556),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_498),
.B(n_204),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_498),
.B(n_269),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_475),
.B(n_226),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_498),
.B(n_269),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_475),
.B(n_235),
.Y(n_722)
);

BUFx6f_ASAP7_75t_SL g723 ( 
.A(n_482),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_589),
.B(n_238),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_498),
.B(n_242),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_527),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_482),
.A2(n_194),
.B1(n_304),
.B2(n_302),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_520),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_482),
.B(n_235),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_482),
.A2(n_188),
.B1(n_300),
.B2(n_205),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_482),
.B(n_246),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_556),
.Y(n_732)
);

INVxp33_ASAP7_75t_L g733 ( 
.A(n_551),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_458),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_570),
.A2(n_184),
.B1(n_189),
.B2(n_202),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_527),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_504),
.Y(n_737)
);

INVx8_ASAP7_75t_L g738 ( 
.A(n_503),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_556),
.B(n_290),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_531),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_556),
.B(n_290),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_504),
.B(n_247),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_531),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_559),
.B(n_246),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_595),
.A2(n_261),
.B1(n_296),
.B2(n_295),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_533),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_581),
.A2(n_261),
.B1(n_296),
.B2(n_295),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_503),
.B(n_509),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_533),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_503),
.B(n_248),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_509),
.B(n_253),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_509),
.B(n_587),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_547),
.B(n_258),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_654),
.A2(n_580),
.B(n_583),
.C(n_539),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_684),
.A2(n_524),
.B(n_516),
.Y(n_755)
);

OAI21xp5_ASAP7_75t_L g756 ( 
.A1(n_653),
.A2(n_585),
.B(n_524),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_675),
.A2(n_524),
.B(n_516),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_671),
.B(n_501),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_681),
.B(n_516),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_675),
.A2(n_544),
.B(n_525),
.Y(n_760)
);

AO21x1_ASAP7_75t_L g761 ( 
.A1(n_672),
.A2(n_563),
.B(n_539),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_615),
.Y(n_762)
);

NAND2x1p5_ASAP7_75t_L g763 ( 
.A(n_615),
.B(n_537),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_SL g764 ( 
.A1(n_633),
.A2(n_541),
.B(n_593),
.C(n_537),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_599),
.B(n_595),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_672),
.A2(n_544),
.B(n_525),
.Y(n_766)
);

OAI21xp5_ASAP7_75t_L g767 ( 
.A1(n_748),
.A2(n_585),
.B(n_545),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_SL g768 ( 
.A(n_713),
.B(n_670),
.C(n_600),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_601),
.B(n_615),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_606),
.Y(n_770)
);

OAI21xp33_ASAP7_75t_L g771 ( 
.A1(n_654),
.A2(n_277),
.B(n_255),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_660),
.A2(n_552),
.B(n_593),
.C(n_541),
.Y(n_772)
);

AO21x1_ASAP7_75t_L g773 ( 
.A1(n_596),
.A2(n_563),
.B(n_552),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_596),
.A2(n_573),
.B1(n_553),
.B2(n_545),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_614),
.A2(n_573),
.B1(n_553),
.B2(n_569),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_689),
.B(n_595),
.Y(n_776)
);

AO21x1_ASAP7_75t_L g777 ( 
.A1(n_614),
.A2(n_569),
.B(n_557),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_676),
.A2(n_557),
.B(n_584),
.C(n_505),
.Y(n_778)
);

NOR2xp67_ASAP7_75t_L g779 ( 
.A(n_626),
.B(n_630),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_615),
.B(n_616),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_690),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_697),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_616),
.B(n_556),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_598),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_687),
.B(n_590),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_629),
.A2(n_499),
.B(n_491),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_705),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_689),
.B(n_584),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_648),
.B(n_459),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_648),
.B(n_470),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_706),
.A2(n_511),
.B(n_491),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_656),
.B(n_470),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_652),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_603),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_673),
.A2(n_265),
.B(n_289),
.C(n_291),
.Y(n_795)
);

BUFx2_ASAP7_75t_SL g796 ( 
.A(n_723),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_663),
.B(n_478),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_625),
.B(n_637),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_737),
.B(n_590),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_707),
.A2(n_523),
.B(n_511),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_664),
.B(n_478),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_665),
.B(n_484),
.Y(n_802)
);

O2A1O1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_667),
.A2(n_258),
.B(n_265),
.C(n_289),
.Y(n_803)
);

INVx5_ASAP7_75t_L g804 ( 
.A(n_604),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_668),
.B(n_484),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_609),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_715),
.A2(n_546),
.B(n_519),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_737),
.B(n_590),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_715),
.A2(n_546),
.B(n_519),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_602),
.B(n_592),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_669),
.B(n_485),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_682),
.B(n_485),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_617),
.A2(n_561),
.B(n_534),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_604),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_695),
.A2(n_534),
.B(n_523),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_682),
.B(n_590),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_617),
.A2(n_538),
.B(n_578),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_618),
.A2(n_538),
.B(n_578),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_734),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_618),
.A2(n_561),
.B(n_558),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_640),
.B(n_536),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_639),
.B(n_536),
.Y(n_822)
);

AO21x1_ASAP7_75t_L g823 ( 
.A1(n_691),
.A2(n_492),
.B(n_483),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_733),
.B(n_536),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_605),
.B(n_610),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_718),
.A2(n_567),
.B(n_560),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_639),
.B(n_543),
.Y(n_827)
);

BUFx12f_ASAP7_75t_L g828 ( 
.A(n_700),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_645),
.B(n_543),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_658),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_645),
.B(n_543),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_632),
.B(n_592),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_718),
.A2(n_558),
.B(n_567),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_701),
.B(n_562),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_719),
.A2(n_560),
.B(n_577),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_634),
.B(n_592),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_701),
.B(n_562),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_604),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_651),
.B(n_562),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_680),
.B(n_688),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_738),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_710),
.B(n_577),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_644),
.A2(n_650),
.B(n_649),
.C(n_628),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_691),
.A2(n_455),
.B(n_454),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_710),
.B(n_577),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_642),
.Y(n_846)
);

AOI21xp33_ASAP7_75t_L g847 ( 
.A1(n_714),
.A2(n_455),
.B(n_494),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_711),
.A2(n_291),
.B(n_494),
.C(n_492),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_719),
.A2(n_483),
.B(n_454),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_725),
.B(n_592),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_635),
.B(n_592),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_721),
.A2(n_488),
.B(n_474),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_641),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_725),
.B(n_456),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_647),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_738),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_703),
.A2(n_674),
.B(n_721),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_613),
.A2(n_488),
.B(n_474),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_696),
.B(n_280),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_619),
.B(n_453),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_752),
.A2(n_554),
.B(n_515),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_738),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_714),
.A2(n_281),
.B(n_294),
.C(n_293),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_677),
.B(n_284),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_623),
.B(n_288),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_611),
.A2(n_555),
.B(n_554),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_679),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_724),
.B(n_716),
.Y(n_868)
);

NOR2x1_ASAP7_75t_R g869 ( 
.A(n_683),
.B(n_159),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_724),
.B(n_720),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_612),
.A2(n_554),
.B(n_515),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_722),
.B(n_160),
.Y(n_872)
);

BUFx4f_ASAP7_75t_L g873 ( 
.A(n_677),
.Y(n_873)
);

INVx11_ASAP7_75t_L g874 ( 
.A(n_693),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_703),
.A2(n_410),
.B(n_554),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_729),
.B(n_166),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_608),
.A2(n_709),
.B(n_662),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_620),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_608),
.A2(n_554),
.B(n_515),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_638),
.B(n_453),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_685),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_677),
.A2(n_234),
.B1(n_169),
.B2(n_174),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_666),
.B(n_7),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_728),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_731),
.B(n_176),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_709),
.A2(n_555),
.B(n_515),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_621),
.B(n_177),
.Y(n_887)
);

INVx8_ASAP7_75t_L g888 ( 
.A(n_723),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_622),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_674),
.A2(n_410),
.B(n_515),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_643),
.A2(n_163),
.B1(n_274),
.B2(n_210),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_L g892 ( 
.A(n_638),
.B(n_410),
.Y(n_892)
);

OAI22xp33_ASAP7_75t_L g893 ( 
.A1(n_708),
.A2(n_163),
.B1(n_186),
.B2(n_195),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_638),
.B(n_453),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_699),
.B(n_195),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_745),
.A2(n_197),
.B1(n_274),
.B2(n_410),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_627),
.Y(n_897)
);

NOR3xp33_ASAP7_75t_L g898 ( 
.A(n_661),
.B(n_257),
.C(n_250),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_657),
.A2(n_453),
.B(n_555),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_624),
.B(n_181),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_686),
.B(n_182),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_686),
.B(n_183),
.Y(n_902)
);

AO21x1_ASAP7_75t_L g903 ( 
.A1(n_739),
.A2(n_168),
.B(n_268),
.Y(n_903)
);

NAND2x1_ASAP7_75t_L g904 ( 
.A(n_728),
.B(n_268),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_646),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_631),
.A2(n_555),
.B(n_453),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_597),
.B(n_185),
.Y(n_907)
);

NAND3xp33_ASAP7_75t_SL g908 ( 
.A(n_698),
.B(n_236),
.C(n_233),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_694),
.Y(n_909)
);

INVx3_ASAP7_75t_SL g910 ( 
.A(n_753),
.Y(n_910)
);

AO21x1_ASAP7_75t_L g911 ( 
.A1(n_739),
.A2(n_168),
.B(n_268),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_597),
.B(n_225),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_702),
.A2(n_555),
.B(n_287),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_712),
.A2(n_740),
.B(n_736),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_726),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_704),
.B(n_7),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_638),
.B(n_168),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_753),
.B(n_8),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_743),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_750),
.B(n_286),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_746),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_636),
.A2(n_646),
.B1(n_749),
.B2(n_750),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_751),
.B(n_285),
.Y(n_923)
);

AOI33xp33_ASAP7_75t_L g924 ( 
.A1(n_747),
.A2(n_8),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.B3(n_14),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_751),
.A2(n_732),
.B(n_678),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_636),
.B(n_12),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_655),
.A2(n_732),
.B(n_717),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_655),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_655),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_659),
.Y(n_930)
);

BUFx5_ASAP7_75t_L g931 ( 
.A(n_659),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_SL g932 ( 
.A(n_828),
.B(n_838),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_850),
.A2(n_732),
.B(n_678),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_798),
.B(n_607),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_868),
.A2(n_730),
.B(n_727),
.C(n_745),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_788),
.B(n_659),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_784),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_870),
.A2(n_732),
.B1(n_692),
.B2(n_717),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_919),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_793),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_922),
.B(n_659),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_854),
.A2(n_678),
.B(n_717),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_926),
.A2(n_735),
.B1(n_742),
.B2(n_744),
.Y(n_943)
);

INVx3_ASAP7_75t_SL g944 ( 
.A(n_782),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_925),
.A2(n_741),
.B(n_692),
.Y(n_945)
);

BUFx8_ASAP7_75t_SL g946 ( 
.A(n_918),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_910),
.B(n_758),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_840),
.B(n_698),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_921),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_910),
.B(n_15),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_759),
.A2(n_692),
.B1(n_282),
.B2(n_279),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_770),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_767),
.A2(n_168),
.B(n_268),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_853),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_863),
.A2(n_15),
.B(n_19),
.C(n_22),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_853),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_856),
.Y(n_957)
);

O2A1O1Ixp5_ASAP7_75t_L g958 ( 
.A1(n_777),
.A2(n_168),
.B(n_23),
.C(n_24),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_863),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_856),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_840),
.B(n_26),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_865),
.B(n_26),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_794),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_804),
.B(n_268),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_L g965 ( 
.A1(n_823),
.A2(n_761),
.B(n_773),
.C(n_756),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_830),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_766),
.A2(n_262),
.B(n_259),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_765),
.A2(n_244),
.B(n_241),
.Y(n_968)
);

CKINVDCx8_ASAP7_75t_R g969 ( 
.A(n_796),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_843),
.A2(n_240),
.B(n_230),
.C(n_222),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_785),
.B(n_28),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_781),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_785),
.B(n_30),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_869),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_755),
.A2(n_208),
.B(n_113),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_825),
.B(n_30),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_877),
.A2(n_799),
.B(n_808),
.C(n_916),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_895),
.B(n_31),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_SL g979 ( 
.A(n_768),
.B(n_33),
.C(n_35),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_774),
.A2(n_97),
.B(n_152),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_838),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_776),
.B(n_168),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_825),
.B(n_33),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_814),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_775),
.A2(n_80),
.B(n_149),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_824),
.B(n_36),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_929),
.B(n_168),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_929),
.B(n_168),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_898),
.A2(n_771),
.B(n_859),
.C(n_754),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_888),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_806),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_799),
.B(n_39),
.Y(n_992)
);

OAI22x1_ASAP7_75t_L g993 ( 
.A1(n_864),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_804),
.B(n_43),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_878),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_889),
.Y(n_996)
);

OR2x6_ASAP7_75t_SL g997 ( 
.A(n_901),
.B(n_43),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_807),
.A2(n_59),
.B(n_140),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_834),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_787),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_814),
.Y(n_1001)
);

AO22x1_ASAP7_75t_L g1002 ( 
.A1(n_898),
.A2(n_44),
.B1(n_47),
.B2(n_52),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_920),
.A2(n_44),
.B1(n_56),
.B2(n_57),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_808),
.A2(n_56),
.B(n_58),
.C(n_68),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_824),
.B(n_58),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_883),
.B(n_73),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_809),
.A2(n_79),
.B(n_136),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_797),
.A2(n_143),
.B(n_801),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_883),
.B(n_909),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_802),
.A2(n_811),
.B(n_805),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_927),
.A2(n_757),
.B(n_822),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_916),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_897),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_804),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_859),
.B(n_864),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_874),
.Y(n_1016)
);

BUFx12f_ASAP7_75t_L g1017 ( 
.A(n_804),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_915),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_779),
.B(n_873),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_837),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_827),
.A2(n_829),
.B(n_831),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_862),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_873),
.Y(n_1023)
);

AO221x2_ASAP7_75t_L g1024 ( 
.A1(n_893),
.A2(n_924),
.B1(n_923),
.B2(n_857),
.C(n_891),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_929),
.Y(n_1025)
);

OAI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_882),
.A2(n_789),
.B1(n_790),
.B2(n_893),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_819),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_760),
.A2(n_813),
.B(n_818),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_778),
.B(n_792),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_862),
.B(n_821),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_842),
.A2(n_845),
.B1(n_839),
.B2(n_907),
.Y(n_1031)
);

AO21x2_ASAP7_75t_L g1032 ( 
.A1(n_847),
.A2(n_844),
.B(n_815),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_929),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_803),
.A2(n_772),
.B(n_764),
.C(n_887),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_888),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_821),
.B(n_795),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_795),
.A2(n_914),
.B(n_839),
.C(n_924),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_912),
.A2(n_900),
.B1(n_884),
.B2(n_816),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_812),
.B(n_872),
.Y(n_1039)
);

AND2x2_ASAP7_75t_SL g1040 ( 
.A(n_896),
.B(n_902),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_817),
.A2(n_820),
.B(n_764),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_876),
.B(n_885),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_888),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_884),
.A2(n_763),
.B1(n_905),
.B2(n_762),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_846),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_762),
.B(n_905),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_930),
.B(n_931),
.Y(n_1047)
);

INVx5_ASAP7_75t_L g1048 ( 
.A(n_930),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_930),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_763),
.A2(n_841),
.B1(n_930),
.B2(n_928),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_855),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_769),
.Y(n_1052)
);

AND2x2_ASAP7_75t_SL g1053 ( 
.A(n_896),
.B(n_892),
.Y(n_1053)
);

O2A1O1Ixp5_ASAP7_75t_L g1054 ( 
.A1(n_917),
.A2(n_851),
.B(n_836),
.C(n_832),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_769),
.B(n_810),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_867),
.B(n_881),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_931),
.B(n_913),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_SL g1058 ( 
.A1(n_904),
.A2(n_841),
.B1(n_908),
.B2(n_890),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_848),
.B(n_810),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_931),
.B(n_780),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_791),
.A2(n_800),
.B(n_833),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_880),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_880),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_894),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_780),
.B(n_832),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_836),
.B(n_851),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_848),
.A2(n_858),
.B(n_786),
.C(n_852),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_931),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_860),
.A2(n_783),
.B1(n_917),
.B2(n_903),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_931),
.B(n_783),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_931),
.Y(n_1071)
);

AO32x2_ASAP7_75t_L g1072 ( 
.A1(n_911),
.A2(n_860),
.A3(n_826),
.B1(n_849),
.B2(n_835),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_894),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_879),
.B(n_875),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_899),
.B(n_866),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1015),
.B(n_1012),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1015),
.B(n_871),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_969),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_1016),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_989),
.A2(n_906),
.B(n_886),
.C(n_861),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_934),
.B(n_954),
.Y(n_1081)
);

INVx5_ASAP7_75t_L g1082 ( 
.A(n_1014),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_954),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1021),
.A2(n_1010),
.B(n_977),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_1041),
.A2(n_1011),
.B(n_1028),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_SL g1086 ( 
.A1(n_1029),
.A2(n_1006),
.B(n_935),
.Y(n_1086)
);

O2A1O1Ixp5_ASAP7_75t_L g1087 ( 
.A1(n_1057),
.A2(n_965),
.B(n_941),
.C(n_1026),
.Y(n_1087)
);

AOI31xp67_ASAP7_75t_L g1088 ( 
.A1(n_1075),
.A2(n_941),
.A3(n_1057),
.B(n_936),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1039),
.B(n_1009),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_953),
.A2(n_945),
.B(n_1061),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_937),
.Y(n_1091)
);

INVx3_ASAP7_75t_SL g1092 ( 
.A(n_944),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_965),
.A2(n_1037),
.B(n_983),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_942),
.A2(n_1074),
.B(n_933),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1012),
.A2(n_961),
.B(n_948),
.C(n_1026),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_SL g1096 ( 
.A1(n_992),
.A2(n_1004),
.B(n_971),
.C(n_973),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_940),
.B(n_956),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_SL g1098 ( 
.A1(n_970),
.A2(n_1042),
.B(n_1070),
.C(n_1047),
.Y(n_1098)
);

AOI221x1_ASAP7_75t_L g1099 ( 
.A1(n_993),
.A2(n_1003),
.B1(n_1005),
.B2(n_986),
.C(n_976),
.Y(n_1099)
);

BUFx12f_ASAP7_75t_L g1100 ( 
.A(n_974),
.Y(n_1100)
);

AND2x6_ASAP7_75t_L g1101 ( 
.A(n_994),
.B(n_1059),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_947),
.B(n_994),
.Y(n_1102)
);

OAI22x1_ASAP7_75t_L g1103 ( 
.A1(n_947),
.A2(n_943),
.B1(n_983),
.B2(n_976),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1008),
.A2(n_1067),
.B(n_938),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_956),
.B(n_949),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_SL g1106 ( 
.A1(n_1031),
.A2(n_1038),
.B(n_1036),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_963),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_975),
.A2(n_985),
.B(n_980),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_1030),
.B(n_1035),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_966),
.B(n_952),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_990),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_991),
.B(n_995),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_996),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_986),
.A2(n_1005),
.B1(n_1053),
.B2(n_978),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_984),
.Y(n_1116)
);

INVx3_ASAP7_75t_SL g1117 ( 
.A(n_944),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1034),
.A2(n_959),
.B(n_955),
.C(n_958),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1013),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1020),
.B(n_999),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_1001),
.B(n_946),
.Y(n_1121)
);

O2A1O1Ixp5_ASAP7_75t_SL g1122 ( 
.A1(n_982),
.A2(n_987),
.B(n_988),
.C(n_936),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1018),
.B(n_1023),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_958),
.A2(n_962),
.B(n_979),
.C(n_950),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1043),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_1055),
.A2(n_1065),
.B(n_1053),
.C(n_1066),
.Y(n_1126)
);

AOI221x1_ASAP7_75t_L g1127 ( 
.A1(n_1055),
.A2(n_1066),
.B1(n_998),
.B2(n_1007),
.C(n_1065),
.Y(n_1127)
);

INVx3_ASAP7_75t_SL g1128 ( 
.A(n_1035),
.Y(n_1128)
);

CKINVDCx6p67_ASAP7_75t_R g1129 ( 
.A(n_997),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1049),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_979),
.B(n_1019),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1024),
.A2(n_1040),
.B1(n_1002),
.B2(n_932),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1045),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1070),
.A2(n_1047),
.B(n_1060),
.Y(n_1134)
);

NOR2x1_ASAP7_75t_L g1135 ( 
.A(n_1022),
.B(n_981),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1054),
.A2(n_982),
.B(n_1068),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1054),
.A2(n_1040),
.B(n_968),
.C(n_1052),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1049),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1024),
.B(n_1052),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_1056),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_1017),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1032),
.A2(n_1071),
.B(n_1044),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1048),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1025),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1032),
.A2(n_1058),
.B(n_1068),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_981),
.B(n_1048),
.Y(n_1146)
);

AO32x2_ASAP7_75t_L g1147 ( 
.A1(n_1050),
.A2(n_1024),
.A3(n_951),
.B1(n_1072),
.B2(n_1069),
.Y(n_1147)
);

OAI22x1_ASAP7_75t_L g1148 ( 
.A1(n_1073),
.A2(n_1051),
.B1(n_1027),
.B2(n_1000),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_972),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1062),
.B(n_1064),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1062),
.B(n_1064),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1048),
.B(n_1064),
.Y(n_1152)
);

INVxp67_ASAP7_75t_L g1153 ( 
.A(n_1046),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1048),
.A2(n_967),
.B(n_1033),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1062),
.B(n_1064),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_957),
.B(n_960),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_957),
.A2(n_960),
.B1(n_964),
.B2(n_1062),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1063),
.A2(n_1025),
.B1(n_1033),
.B2(n_1072),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1063),
.B(n_1025),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1072),
.A2(n_1063),
.B(n_1033),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1063),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1021),
.A2(n_850),
.B(n_854),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_965),
.A2(n_977),
.B(n_601),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1015),
.A2(n_601),
.B(n_989),
.C(n_654),
.Y(n_1164)
);

CKINVDCx11_ASAP7_75t_R g1165 ( 
.A(n_969),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_1021),
.A2(n_823),
.A3(n_777),
.B(n_773),
.Y(n_1166)
);

O2A1O1Ixp5_ASAP7_75t_SL g1167 ( 
.A1(n_982),
.A2(n_988),
.B(n_987),
.C(n_936),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_977),
.A2(n_633),
.B(n_601),
.C(n_1006),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1041),
.A2(n_1011),
.B(n_1028),
.Y(n_1169)
);

AO21x1_ASAP7_75t_L g1170 ( 
.A1(n_1026),
.A2(n_1006),
.B(n_1015),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1015),
.A2(n_607),
.B1(n_586),
.B2(n_926),
.Y(n_1171)
);

BUFx12f_ASAP7_75t_L g1172 ( 
.A(n_1016),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_940),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1041),
.A2(n_1011),
.B(n_1028),
.Y(n_1174)
);

AOI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1041),
.A2(n_1011),
.B(n_1075),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1021),
.A2(n_850),
.B(n_854),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1015),
.A2(n_601),
.B(n_989),
.C(n_654),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1015),
.A2(n_601),
.B(n_989),
.C(n_654),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1021),
.A2(n_850),
.B(n_854),
.Y(n_1179)
);

AOI221x1_ASAP7_75t_L g1180 ( 
.A1(n_1015),
.A2(n_993),
.B1(n_1004),
.B2(n_1003),
.C(n_935),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_937),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1021),
.A2(n_850),
.B(n_854),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1021),
.A2(n_850),
.B(n_854),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_940),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_937),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1015),
.A2(n_601),
.B1(n_961),
.B2(n_926),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1021),
.A2(n_850),
.B(n_854),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1021),
.A2(n_823),
.A3(n_777),
.B(n_773),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1015),
.B(n_948),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1041),
.A2(n_1011),
.B(n_1028),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1015),
.A2(n_654),
.B1(n_601),
.B2(n_1026),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1041),
.A2(n_1011),
.B(n_1028),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1029),
.B(n_825),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1041),
.A2(n_1011),
.B(n_1028),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1015),
.A2(n_601),
.B1(n_961),
.B2(n_926),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_990),
.Y(n_1196)
);

AOI31xp67_ASAP7_75t_L g1197 ( 
.A1(n_1075),
.A2(n_941),
.A3(n_1057),
.B(n_936),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1041),
.A2(n_1011),
.B(n_1028),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_939),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1021),
.A2(n_850),
.B(n_854),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1021),
.A2(n_823),
.A3(n_777),
.B(n_773),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1015),
.A2(n_607),
.B1(n_586),
.B2(n_926),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1015),
.B(n_948),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1021),
.A2(n_850),
.B(n_854),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1015),
.A2(n_601),
.B(n_989),
.C(n_654),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1021),
.A2(n_823),
.A3(n_777),
.B(n_773),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1021),
.A2(n_850),
.B(n_854),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_940),
.B(n_572),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1015),
.A2(n_654),
.B(n_601),
.C(n_461),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1021),
.A2(n_850),
.B(n_854),
.Y(n_1210)
);

AO21x2_ASAP7_75t_L g1211 ( 
.A1(n_982),
.A2(n_1061),
.B(n_1032),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1015),
.B(n_654),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1021),
.A2(n_850),
.B(n_854),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1041),
.A2(n_1011),
.B(n_1028),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_965),
.A2(n_977),
.B(n_601),
.Y(n_1215)
);

NOR4xp25_ASAP7_75t_L g1216 ( 
.A(n_955),
.B(n_924),
.C(n_959),
.D(n_1026),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_1021),
.A2(n_823),
.A3(n_777),
.B(n_773),
.Y(n_1217)
);

BUFx2_ASAP7_75t_R g1218 ( 
.A(n_969),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1029),
.B(n_825),
.Y(n_1219)
);

AO21x2_ASAP7_75t_L g1220 ( 
.A1(n_982),
.A2(n_1061),
.B(n_1032),
.Y(n_1220)
);

CKINVDCx16_ASAP7_75t_R g1221 ( 
.A(n_1078),
.Y(n_1221)
);

CKINVDCx11_ASAP7_75t_R g1222 ( 
.A(n_1165),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1113),
.Y(n_1223)
);

OAI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1132),
.A2(n_1191),
.B1(n_1115),
.B2(n_1212),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1218),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1076),
.B(n_1089),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1171),
.A2(n_1202),
.B1(n_1115),
.B2(n_1186),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1101),
.Y(n_1228)
);

INVx4_ASAP7_75t_SL g1229 ( 
.A(n_1101),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1109),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1091),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1097),
.B(n_1083),
.Y(n_1232)
);

CKINVDCx11_ASAP7_75t_R g1233 ( 
.A(n_1092),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1109),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1211),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1089),
.B(n_1189),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1186),
.A2(n_1195),
.B1(n_1103),
.B2(n_1170),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1107),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1203),
.B(n_1120),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1114),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1211),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1117),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1164),
.A2(n_1205),
.B1(n_1177),
.B2(n_1178),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1195),
.A2(n_1129),
.B1(n_1093),
.B2(n_1101),
.Y(n_1244)
);

INVxp67_ASAP7_75t_SL g1245 ( 
.A(n_1105),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1119),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1093),
.A2(n_1101),
.B1(n_1081),
.B2(n_1139),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1220),
.Y(n_1248)
);

AOI22x1_ASAP7_75t_SL g1249 ( 
.A1(n_1173),
.A2(n_1116),
.B1(n_1181),
.B2(n_1185),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1220),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_SL g1251 ( 
.A1(n_1099),
.A2(n_1180),
.B(n_1209),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1161),
.B(n_1150),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1139),
.A2(n_1131),
.B1(n_1140),
.B2(n_1163),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1133),
.Y(n_1254)
);

CKINVDCx6p67_ASAP7_75t_R g1255 ( 
.A(n_1082),
.Y(n_1255)
);

BUFx10_ASAP7_75t_L g1256 ( 
.A(n_1121),
.Y(n_1256)
);

BUFx12f_ASAP7_75t_L g1257 ( 
.A(n_1100),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1079),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1172),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1173),
.B(n_1193),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1163),
.A2(n_1215),
.B1(n_1219),
.B2(n_1193),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1184),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1126),
.A2(n_1118),
.B1(n_1086),
.B2(n_1095),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1219),
.B(n_1111),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1116),
.B(n_1208),
.Y(n_1265)
);

CKINVDCx11_ASAP7_75t_R g1266 ( 
.A(n_1128),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1123),
.Y(n_1267)
);

CKINVDCx6p67_ASAP7_75t_R g1268 ( 
.A(n_1082),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1215),
.A2(n_1102),
.B1(n_1199),
.B2(n_1149),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1148),
.A2(n_1153),
.B1(n_1216),
.B2(n_1077),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1125),
.Y(n_1271)
);

INVx5_ASAP7_75t_L g1272 ( 
.A(n_1143),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1110),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1216),
.A2(n_1084),
.B1(n_1155),
.B2(n_1130),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1138),
.A2(n_1104),
.B1(n_1150),
.B2(n_1151),
.Y(n_1275)
);

CKINVDCx6p67_ASAP7_75t_R g1276 ( 
.A(n_1146),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_1141),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1146),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1124),
.A2(n_1106),
.B1(n_1137),
.B2(n_1108),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1143),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1160),
.Y(n_1281)
);

INVx6_ASAP7_75t_L g1282 ( 
.A(n_1156),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1151),
.A2(n_1145),
.B1(n_1179),
.B2(n_1213),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1162),
.A2(n_1210),
.B1(n_1187),
.B2(n_1200),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1176),
.A2(n_1183),
.B1(n_1182),
.B2(n_1204),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1157),
.Y(n_1286)
);

BUFx8_ASAP7_75t_L g1287 ( 
.A(n_1112),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1207),
.A2(n_1142),
.B1(n_1159),
.B2(n_1158),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1196),
.B(n_1135),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_SL g1290 ( 
.A1(n_1147),
.A2(n_1096),
.B1(n_1087),
.B2(n_1144),
.Y(n_1290)
);

BUFx12f_ASAP7_75t_L g1291 ( 
.A(n_1152),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1136),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1158),
.A2(n_1134),
.B1(n_1147),
.B2(n_1154),
.Y(n_1293)
);

BUFx12f_ASAP7_75t_L g1294 ( 
.A(n_1098),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1090),
.A2(n_1094),
.B1(n_1127),
.B2(n_1168),
.Y(n_1295)
);

INVx6_ASAP7_75t_L g1296 ( 
.A(n_1088),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1085),
.A2(n_1190),
.B1(n_1192),
.B2(n_1214),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1175),
.A2(n_1122),
.B1(n_1167),
.B2(n_1197),
.Y(n_1298)
);

CKINVDCx11_ASAP7_75t_R g1299 ( 
.A(n_1166),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1169),
.A2(n_1194),
.B1(n_1198),
.B2(n_1174),
.Y(n_1300)
);

BUFx12f_ASAP7_75t_L g1301 ( 
.A(n_1166),
.Y(n_1301)
);

INVx8_ASAP7_75t_L g1302 ( 
.A(n_1080),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1188),
.A2(n_1201),
.B1(n_1206),
.B2(n_1217),
.Y(n_1303)
);

CKINVDCx11_ASAP7_75t_R g1304 ( 
.A(n_1188),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1201),
.A2(n_1202),
.B1(n_1171),
.B2(n_1115),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1201),
.A2(n_1202),
.B1(n_1171),
.B2(n_1115),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1206),
.A2(n_1132),
.B1(n_1191),
.B2(n_1015),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1217),
.B(n_1212),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1097),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1113),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1165),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1115),
.A2(n_1015),
.B1(n_571),
.B2(n_1186),
.Y(n_1312)
);

INVx5_ASAP7_75t_L g1313 ( 
.A(n_1101),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1113),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1165),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1115),
.A2(n_1015),
.B1(n_713),
.B2(n_600),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1171),
.A2(n_1202),
.B1(n_1115),
.B2(n_926),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1113),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1171),
.A2(n_1202),
.B1(n_1115),
.B2(n_926),
.Y(n_1319)
);

BUFx8_ASAP7_75t_L g1320 ( 
.A(n_1125),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1171),
.A2(n_1202),
.B1(n_1115),
.B2(n_926),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1113),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1113),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1165),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_SL g1325 ( 
.A1(n_1115),
.A2(n_1015),
.B1(n_571),
.B2(n_1186),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1208),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1146),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1171),
.A2(n_1202),
.B1(n_1115),
.B2(n_926),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1081),
.B(n_1076),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1109),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1212),
.A2(n_1015),
.B1(n_1191),
.B2(n_601),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1109),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1132),
.A2(n_1191),
.B1(n_1015),
.B2(n_1115),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1083),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1101),
.Y(n_1335)
);

BUFx8_ASAP7_75t_L g1336 ( 
.A(n_1079),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1165),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_1165),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1146),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1113),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1115),
.A2(n_1015),
.B1(n_571),
.B2(n_1186),
.Y(n_1341)
);

BUFx2_ASAP7_75t_R g1342 ( 
.A(n_1092),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1113),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1296),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1316),
.A2(n_1312),
.B1(n_1325),
.B2(n_1341),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1273),
.Y(n_1346)
);

INVxp67_ASAP7_75t_SL g1347 ( 
.A(n_1334),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1297),
.A2(n_1300),
.B(n_1285),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1308),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1226),
.B(n_1329),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1297),
.A2(n_1300),
.B(n_1285),
.Y(n_1351)
);

AO21x1_ASAP7_75t_SL g1352 ( 
.A1(n_1237),
.A2(n_1227),
.B(n_1244),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1284),
.A2(n_1295),
.B(n_1283),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1284),
.A2(n_1295),
.B(n_1279),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1231),
.B(n_1238),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1296),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1283),
.A2(n_1292),
.B(n_1248),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1263),
.A2(n_1333),
.B(n_1243),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1232),
.B(n_1309),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1240),
.B(n_1246),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1282),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1292),
.A2(n_1250),
.B(n_1235),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1282),
.Y(n_1363)
);

BUFx8_ASAP7_75t_SL g1364 ( 
.A(n_1337),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1261),
.B(n_1237),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1302),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1303),
.B(n_1245),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1221),
.B(n_1271),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1254),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1267),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1264),
.B(n_1260),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1278),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1265),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1241),
.A2(n_1250),
.B(n_1248),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1261),
.B(n_1247),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1302),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1262),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1301),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1288),
.A2(n_1281),
.B(n_1293),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1301),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1331),
.A2(n_1251),
.B(n_1224),
.Y(n_1381)
);

INVxp67_ASAP7_75t_SL g1382 ( 
.A(n_1307),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1239),
.B(n_1236),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1223),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1310),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1313),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1298),
.A2(n_1227),
.B(n_1244),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1314),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1318),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1322),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1305),
.A2(n_1306),
.B(n_1270),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1323),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1252),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1340),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1343),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1313),
.B(n_1229),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1247),
.B(n_1253),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1288),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1253),
.B(n_1306),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1305),
.B(n_1304),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1299),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1275),
.A2(n_1274),
.B(n_1270),
.Y(n_1402)
);

INVxp67_ASAP7_75t_SL g1403 ( 
.A(n_1274),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1290),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1269),
.A2(n_1327),
.B(n_1339),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1269),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1342),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1294),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1317),
.B(n_1319),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1369),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1359),
.B(n_1326),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1359),
.B(n_1256),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1347),
.B(n_1319),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1370),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1348),
.A2(n_1351),
.B(n_1354),
.Y(n_1415)
);

A2O1A1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1345),
.A2(n_1317),
.B(n_1321),
.C(n_1328),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1349),
.B(n_1294),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1358),
.A2(n_1228),
.B1(n_1335),
.B2(n_1328),
.Y(n_1418)
);

AND2x6_ASAP7_75t_L g1419 ( 
.A(n_1396),
.B(n_1335),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1372),
.B(n_1256),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1372),
.B(n_1225),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1381),
.A2(n_1289),
.B(n_1272),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1369),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1348),
.A2(n_1351),
.B(n_1354),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1382),
.A2(n_1403),
.B1(n_1365),
.B2(n_1391),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1355),
.B(n_1360),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1346),
.B(n_1324),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1373),
.B(n_1330),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1355),
.B(n_1332),
.Y(n_1429)
);

INVx4_ASAP7_75t_L g1430 ( 
.A(n_1408),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1379),
.A2(n_1249),
.B(n_1286),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1349),
.B(n_1280),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1397),
.A2(n_1399),
.B(n_1387),
.C(n_1365),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1398),
.B(n_1280),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1399),
.A2(n_1330),
.B(n_1230),
.C(n_1332),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1375),
.A2(n_1234),
.B(n_1258),
.C(n_1277),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1375),
.A2(n_1258),
.B(n_1259),
.C(n_1242),
.Y(n_1437)
);

AO32x2_ASAP7_75t_L g1438 ( 
.A1(n_1393),
.A2(n_1324),
.A3(n_1320),
.B1(n_1255),
.B2(n_1268),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1384),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_1364),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_SL g1441 ( 
.A(n_1396),
.B(n_1276),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_SL g1442 ( 
.A1(n_1407),
.A2(n_1377),
.B(n_1368),
.C(n_1383),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1400),
.A2(n_1336),
.B(n_1291),
.C(n_1311),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1357),
.A2(n_1320),
.B(n_1287),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1398),
.B(n_1287),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1400),
.A2(n_1336),
.B(n_1311),
.C(n_1257),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1409),
.A2(n_1257),
.B1(n_1287),
.B2(n_1233),
.Y(n_1447)
);

INVx4_ASAP7_75t_L g1448 ( 
.A(n_1408),
.Y(n_1448)
);

OAI211xp5_ASAP7_75t_L g1449 ( 
.A1(n_1402),
.A2(n_1266),
.B(n_1338),
.C(n_1315),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1350),
.B(n_1222),
.Y(n_1450)
);

NOR2x1_ASAP7_75t_SL g1451 ( 
.A(n_1352),
.B(n_1336),
.Y(n_1451)
);

A2O1A1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1404),
.A2(n_1409),
.B(n_1406),
.C(n_1401),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1402),
.A2(n_1404),
.B1(n_1376),
.B2(n_1366),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1402),
.A2(n_1353),
.B(n_1406),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1361),
.B(n_1363),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1378),
.B(n_1380),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1384),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1361),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1371),
.B(n_1363),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1395),
.B(n_1402),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1362),
.A2(n_1374),
.B(n_1405),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1366),
.A2(n_1376),
.B1(n_1352),
.B2(n_1367),
.Y(n_1462)
);

A2O1A1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1401),
.A2(n_1367),
.B(n_1366),
.C(n_1376),
.Y(n_1463)
);

OAI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1353),
.A2(n_1392),
.B1(n_1390),
.B2(n_1394),
.C(n_1389),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1385),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1378),
.B(n_1380),
.Y(n_1466)
);

OR2x6_ASAP7_75t_L g1467 ( 
.A(n_1396),
.B(n_1386),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1467),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1426),
.B(n_1353),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1460),
.B(n_1388),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1410),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1416),
.A2(n_1353),
.B(n_1441),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1461),
.Y(n_1473)
);

NOR2xp67_ASAP7_75t_L g1474 ( 
.A(n_1464),
.B(n_1376),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1439),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1444),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1423),
.Y(n_1477)
);

NAND2xp33_ASAP7_75t_R g1478 ( 
.A(n_1431),
.B(n_1396),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1457),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1415),
.B(n_1344),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1460),
.B(n_1388),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1465),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1415),
.B(n_1356),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1424),
.B(n_1356),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1461),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1414),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1458),
.B(n_1392),
.Y(n_1487)
);

BUFx8_ASAP7_75t_L g1488 ( 
.A(n_1438),
.Y(n_1488)
);

NOR2x1_ASAP7_75t_L g1489 ( 
.A(n_1449),
.B(n_1463),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1464),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1444),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1458),
.B(n_1459),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_1434),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1454),
.B(n_1390),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1419),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1434),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1453),
.B(n_1394),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1433),
.A2(n_1425),
.B1(n_1413),
.B2(n_1449),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1473),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1469),
.B(n_1412),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1471),
.Y(n_1501)
);

OAI21xp33_ASAP7_75t_L g1502 ( 
.A1(n_1489),
.A2(n_1425),
.B(n_1452),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1469),
.B(n_1420),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1481),
.B(n_1411),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1498),
.A2(n_1453),
.B1(n_1418),
.B2(n_1462),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1473),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1471),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1473),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1471),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1492),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1477),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1473),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1477),
.Y(n_1513)
);

AOI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1485),
.A2(n_1447),
.B(n_1445),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1477),
.Y(n_1515)
);

AND2x2_ASAP7_75t_SL g1516 ( 
.A(n_1490),
.B(n_1431),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1469),
.B(n_1455),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1479),
.Y(n_1518)
);

NAND3xp33_ASAP7_75t_L g1519 ( 
.A(n_1490),
.B(n_1437),
.C(n_1442),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1475),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1486),
.B(n_1421),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1481),
.B(n_1428),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1493),
.B(n_1417),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1485),
.Y(n_1524)
);

NAND3xp33_ASAP7_75t_L g1525 ( 
.A(n_1490),
.B(n_1445),
.C(n_1417),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1486),
.B(n_1429),
.Y(n_1526)
);

INVx1_ASAP7_75t_SL g1527 ( 
.A(n_1492),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1481),
.B(n_1432),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1494),
.B(n_1432),
.Y(n_1529)
);

INVx4_ASAP7_75t_L g1530 ( 
.A(n_1495),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1475),
.Y(n_1531)
);

AOI221x1_ASAP7_75t_L g1532 ( 
.A1(n_1498),
.A2(n_1447),
.B1(n_1446),
.B2(n_1462),
.C(n_1422),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1468),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1493),
.B(n_1430),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1487),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1496),
.B(n_1430),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1488),
.A2(n_1451),
.B1(n_1422),
.B2(n_1441),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1468),
.B(n_1448),
.Y(n_1538)
);

OAI221xp5_ASAP7_75t_SL g1539 ( 
.A1(n_1472),
.A2(n_1436),
.B1(n_1443),
.B2(n_1450),
.C(n_1435),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1503),
.B(n_1476),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1499),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1501),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1501),
.B(n_1497),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1530),
.B(n_1495),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1529),
.B(n_1470),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1503),
.B(n_1476),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1507),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1507),
.B(n_1497),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1530),
.B(n_1495),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1500),
.B(n_1476),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1500),
.B(n_1480),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1506),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1530),
.B(n_1480),
.Y(n_1553)
);

INVxp67_ASAP7_75t_SL g1554 ( 
.A(n_1506),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1509),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1509),
.B(n_1470),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1530),
.B(n_1495),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1511),
.B(n_1482),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1511),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1513),
.B(n_1482),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1508),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1514),
.B(n_1480),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1514),
.B(n_1483),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1508),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1521),
.B(n_1483),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1513),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1512),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1515),
.B(n_1494),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1515),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1529),
.B(n_1528),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1521),
.B(n_1483),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1526),
.B(n_1520),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1517),
.B(n_1484),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1512),
.Y(n_1574)
);

NAND4xp25_ASAP7_75t_L g1575 ( 
.A(n_1532),
.B(n_1489),
.C(n_1427),
.D(n_1472),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1518),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1544),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1547),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1544),
.A2(n_1505),
.B1(n_1502),
.B2(n_1519),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1575),
.B(n_1510),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1575),
.B(n_1440),
.Y(n_1581)
);

INVxp67_ASAP7_75t_SL g1582 ( 
.A(n_1547),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1542),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1544),
.B(n_1538),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1544),
.B(n_1502),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1570),
.B(n_1504),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1541),
.Y(n_1587)
);

NOR2xp67_ASAP7_75t_SL g1588 ( 
.A(n_1562),
.B(n_1519),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1572),
.B(n_1527),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_1543),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1544),
.B(n_1525),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1544),
.B(n_1538),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1549),
.B(n_1526),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1572),
.B(n_1535),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1572),
.B(n_1525),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1542),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1541),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1542),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1555),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1555),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1570),
.B(n_1504),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1555),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1570),
.B(n_1523),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1559),
.Y(n_1604)
);

INVxp33_ASAP7_75t_L g1605 ( 
.A(n_1549),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1545),
.B(n_1522),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1549),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1549),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1545),
.B(n_1531),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1549),
.B(n_1533),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1562),
.B(n_1532),
.C(n_1505),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1545),
.B(n_1543),
.Y(n_1612)
);

NOR3xp33_ASAP7_75t_SL g1613 ( 
.A(n_1548),
.B(n_1539),
.C(n_1536),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1549),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1548),
.B(n_1496),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1557),
.B(n_1533),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1573),
.B(n_1522),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1573),
.B(n_1518),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1619)
);

NAND4xp75_ASAP7_75t_L g1620 ( 
.A(n_1613),
.B(n_1516),
.C(n_1562),
.D(n_1563),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1583),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1593),
.B(n_1557),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1588),
.B(n_1573),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1586),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1581),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1588),
.B(n_1573),
.Y(n_1626)
);

INVxp33_ASAP7_75t_L g1627 ( 
.A(n_1591),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1580),
.B(n_1562),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1586),
.B(n_1568),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1590),
.B(n_1563),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1579),
.B(n_1563),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1578),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1593),
.B(n_1557),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1594),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1611),
.B(n_1565),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1583),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1598),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1601),
.B(n_1568),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1598),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1599),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1585),
.B(n_1553),
.C(n_1474),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1599),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1600),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1600),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_L g1645 ( 
.A(n_1595),
.B(n_1553),
.C(n_1474),
.Y(n_1645)
);

NAND4xp25_ASAP7_75t_L g1646 ( 
.A(n_1577),
.B(n_1553),
.C(n_1557),
.D(n_1540),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1589),
.B(n_1565),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1584),
.B(n_1557),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1601),
.B(n_1556),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1584),
.B(n_1550),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1602),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1592),
.B(n_1550),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1592),
.B(n_1550),
.Y(n_1653)
);

AOI211xp5_ASAP7_75t_SL g1654 ( 
.A1(n_1582),
.A2(n_1553),
.B(n_1540),
.C(n_1546),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1612),
.B(n_1565),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1622),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1620),
.A2(n_1516),
.B1(n_1478),
.B2(n_1488),
.Y(n_1657)
);

AOI222xp33_ASAP7_75t_L g1658 ( 
.A1(n_1635),
.A2(n_1516),
.B1(n_1554),
.B2(n_1615),
.C1(n_1603),
.C2(n_1574),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1631),
.A2(n_1578),
.B(n_1609),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1625),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1624),
.B(n_1634),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1621),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1632),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1621),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1639),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1624),
.B(n_1612),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1639),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1627),
.A2(n_1488),
.B1(n_1587),
.B2(n_1597),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1628),
.A2(n_1602),
.B1(n_1604),
.B2(n_1554),
.C(n_1596),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1649),
.B(n_1629),
.Y(n_1670)
);

NAND4xp75_ASAP7_75t_L g1671 ( 
.A(n_1623),
.B(n_1607),
.C(n_1610),
.D(n_1616),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1622),
.B(n_1619),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1620),
.B(n_1606),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1626),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1646),
.B(n_1608),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1650),
.B(n_1652),
.Y(n_1676)
);

NAND4xp25_ASAP7_75t_L g1677 ( 
.A(n_1654),
.B(n_1614),
.C(n_1610),
.D(n_1616),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1649),
.B(n_1606),
.Y(n_1678)
);

NAND2x1_ASAP7_75t_L g1679 ( 
.A(n_1633),
.B(n_1607),
.Y(n_1679)
);

OAI322xp33_ASAP7_75t_L g1680 ( 
.A1(n_1630),
.A2(n_1604),
.A3(n_1617),
.B1(n_1618),
.B2(n_1587),
.C1(n_1597),
.C2(n_1556),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1640),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1633),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1678),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1660),
.B(n_1605),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1658),
.B(n_1663),
.C(n_1669),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1672),
.B(n_1650),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1662),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1664),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1665),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1667),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1670),
.B(n_1648),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1673),
.A2(n_1645),
.B1(n_1641),
.B2(n_1655),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1674),
.B(n_1652),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1659),
.B(n_1653),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1682),
.B(n_1653),
.Y(n_1695)
);

OAI322xp33_ASAP7_75t_L g1696 ( 
.A1(n_1659),
.A2(n_1638),
.A3(n_1629),
.B1(n_1651),
.B2(n_1640),
.C1(n_1642),
.C2(n_1643),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1681),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1661),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1657),
.A2(n_1638),
.B1(n_1647),
.B2(n_1651),
.C(n_1642),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1671),
.A2(n_1540),
.B1(n_1546),
.B2(n_1619),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1685),
.A2(n_1663),
.B(n_1675),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_L g1702 ( 
.A(n_1684),
.B(n_1669),
.C(n_1677),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1683),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1695),
.Y(n_1704)
);

A2O1A1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1694),
.A2(n_1668),
.B(n_1666),
.C(n_1679),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1687),
.Y(n_1706)
);

BUFx2_ASAP7_75t_L g1707 ( 
.A(n_1686),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1698),
.B(n_1676),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1688),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1698),
.A2(n_1684),
.B1(n_1692),
.B2(n_1699),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1707),
.B(n_1691),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1710),
.A2(n_1693),
.B1(n_1668),
.B2(n_1682),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_L g1713 ( 
.A(n_1701),
.B(n_1690),
.C(n_1689),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1703),
.Y(n_1714)
);

NOR3xp33_ASAP7_75t_SL g1715 ( 
.A(n_1701),
.B(n_1702),
.C(n_1705),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1704),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_SL g1717 ( 
.A(n_1708),
.B(n_1696),
.Y(n_1717)
);

AND2x4_ASAP7_75t_SL g1718 ( 
.A(n_1706),
.B(n_1656),
.Y(n_1718)
);

O2A1O1Ixp5_ASAP7_75t_SL g1719 ( 
.A1(n_1709),
.A2(n_1697),
.B(n_1643),
.C(n_1700),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1711),
.B(n_1636),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1715),
.A2(n_1644),
.B1(n_1637),
.B2(n_1546),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1717),
.B(n_1680),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1718),
.B(n_1716),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1713),
.Y(n_1724)
);

NAND4xp25_ASAP7_75t_L g1725 ( 
.A(n_1722),
.B(n_1712),
.C(n_1714),
.D(n_1719),
.Y(n_1725)
);

NAND4xp25_ASAP7_75t_L g1726 ( 
.A(n_1723),
.B(n_1540),
.C(n_1448),
.D(n_1537),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1724),
.A2(n_1524),
.B1(n_1574),
.B2(n_1567),
.C(n_1564),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1720),
.Y(n_1728)
);

AOI321xp33_ASAP7_75t_L g1729 ( 
.A1(n_1721),
.A2(n_1491),
.A3(n_1466),
.B1(n_1456),
.B2(n_1552),
.C(n_1561),
.Y(n_1729)
);

AOI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1722),
.A2(n_1524),
.B1(n_1574),
.B2(n_1567),
.C(n_1564),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1728),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1725),
.B(n_1576),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1729),
.B(n_1571),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1727),
.B(n_1559),
.Y(n_1734)
);

NOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1726),
.B(n_1559),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1731),
.B(n_1730),
.C(n_1488),
.Y(n_1736)
);

NOR4xp75_ASAP7_75t_L g1737 ( 
.A(n_1734),
.B(n_1571),
.C(n_1558),
.D(n_1560),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1733),
.B(n_1571),
.Y(n_1738)
);

OAI211xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1736),
.A2(n_1732),
.B(n_1735),
.C(n_1576),
.Y(n_1739)
);

NAND4xp75_ASAP7_75t_L g1740 ( 
.A(n_1739),
.B(n_1738),
.C(n_1737),
.D(n_1551),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1740),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1740),
.Y(n_1742)
);

OA22x2_ASAP7_75t_L g1743 ( 
.A1(n_1742),
.A2(n_1569),
.B1(n_1566),
.B2(n_1576),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1741),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1743),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1744),
.A2(n_1551),
.B(n_1561),
.Y(n_1746)
);

OAI21xp33_ASAP7_75t_L g1747 ( 
.A1(n_1745),
.A2(n_1746),
.B(n_1569),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1747),
.A2(n_1551),
.B1(n_1564),
.B2(n_1567),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1574),
.B1(n_1541),
.B2(n_1567),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1749),
.A2(n_1569),
.B1(n_1566),
.B2(n_1541),
.C(n_1564),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1491),
.B(n_1566),
.C(n_1552),
.Y(n_1751)
);


endmodule