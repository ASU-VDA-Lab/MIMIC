module fake_aes_1844_n_42 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_9), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
INVx1_ASAP7_75t_SL g14 ( .A(n_5), .Y(n_14) );
NOR2xp33_ASAP7_75t_R g15 ( .A(n_5), .B(n_2), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_3), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_8), .Y(n_17) );
OR2x2_ASAP7_75t_L g18 ( .A(n_11), .B(n_0), .Y(n_18) );
AOI21x1_ASAP7_75t_L g19 ( .A1(n_11), .A2(n_10), .B(n_3), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_16), .B(n_1), .C(n_4), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_13), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_13), .Y(n_22) );
BUFx12f_ASAP7_75t_L g23 ( .A(n_18), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_22), .B(n_17), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_21), .B(n_12), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_22), .B1(n_21), .B2(n_18), .Y(n_27) );
OAI31xp33_ASAP7_75t_SL g28 ( .A1(n_25), .A2(n_14), .A3(n_20), .B(n_15), .Y(n_28) );
AOI21x1_ASAP7_75t_L g29 ( .A1(n_24), .A2(n_19), .B(n_21), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_23), .Y(n_30) );
AO21x1_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_19), .B(n_26), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
NOR2xp67_ASAP7_75t_SL g33 ( .A(n_30), .B(n_23), .Y(n_33) );
AOI21xp33_ASAP7_75t_SL g34 ( .A1(n_32), .A2(n_28), .B(n_4), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_33), .B(n_26), .Y(n_35) );
OAI211xp5_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_15), .B(n_20), .C(n_14), .Y(n_36) );
AOI22xp33_ASAP7_75t_SL g37 ( .A1(n_36), .A2(n_24), .B1(n_6), .B2(n_7), .Y(n_37) );
NOR3xp33_ASAP7_75t_SL g38 ( .A(n_35), .B(n_1), .C(n_6), .Y(n_38) );
A2O1A1Ixp33_ASAP7_75t_L g39 ( .A1(n_34), .A2(n_31), .B(n_8), .C(n_7), .Y(n_39) );
CKINVDCx20_ASAP7_75t_R g40 ( .A(n_38), .Y(n_40) );
CKINVDCx20_ASAP7_75t_R g41 ( .A(n_37), .Y(n_41) );
AOI22xp33_ASAP7_75t_SL g42 ( .A1(n_41), .A2(n_29), .B1(n_39), .B2(n_40), .Y(n_42) );
endmodule