module fake_jpeg_13802_n_417 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_417);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_417;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_39),
.B(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_16),
.B(n_15),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_48),
.Y(n_107)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_27),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_66),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_67),
.Y(n_112)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_38),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_70),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_74),
.Y(n_80)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_27),
.Y(n_101)
);

INVx2_ASAP7_75t_R g73 ( 
.A(n_31),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_33),
.CON(n_96),
.SN(n_96)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_18),
.B(n_15),
.Y(n_74)
);

NAND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_53),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_77),
.B(n_41),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_14),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_108),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_90),
.A2(n_102),
.B1(n_106),
.B2(n_41),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_45),
.A2(n_60),
.B1(n_63),
.B2(n_57),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_93),
.A2(n_116),
.B1(n_59),
.B2(n_51),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_101),
.B(n_111),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_48),
.A2(n_26),
.B1(n_36),
.B2(n_35),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_72),
.A2(n_26),
.B1(n_36),
.B2(n_35),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_104),
.A2(n_114),
.B1(n_19),
.B2(n_20),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_26),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_73),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_53),
.A2(n_25),
.B1(n_36),
.B2(n_34),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_73),
.B(n_14),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_14),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_47),
.A2(n_25),
.B1(n_34),
.B2(n_33),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_33),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_119),
.B(n_139),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_120),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_77),
.A2(n_40),
.B1(n_56),
.B2(n_61),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_129),
.B1(n_149),
.B2(n_155),
.Y(n_159)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_54),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_127),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_125),
.B(n_140),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_64),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_77),
.A2(n_25),
.B1(n_20),
.B2(n_34),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_67),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_134),
.C(n_111),
.Y(n_172)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_133),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_68),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_53),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_77),
.A2(n_42),
.B1(n_46),
.B2(n_62),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_147),
.B1(n_150),
.B2(n_157),
.Y(n_168)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_148),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_92),
.B(n_19),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_20),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_153),
.B(n_154),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_44),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_84),
.A2(n_58),
.B1(n_41),
.B2(n_23),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_158),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_114),
.A2(n_55),
.B1(n_52),
.B2(n_49),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_78),
.B1(n_104),
.B2(n_115),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_161),
.A2(n_138),
.B1(n_123),
.B2(n_118),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_175),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_96),
.B(n_113),
.C(n_111),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_139),
.B(n_79),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_78),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_135),
.C(n_141),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_111),
.B1(n_115),
.B2(n_109),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_185),
.B1(n_107),
.B2(n_84),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_122),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_181),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_119),
.A2(n_87),
.B1(n_95),
.B2(n_109),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_107),
.Y(n_211)
);

AO22x1_ASAP7_75t_SL g181 ( 
.A1(n_130),
.A2(n_103),
.B1(n_100),
.B2(n_50),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_87),
.B1(n_79),
.B2(n_95),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_113),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_23),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_79),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_196),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_198),
.B(n_208),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_192),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_205),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_125),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_201),
.B(n_206),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_152),
.B(n_144),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_203),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_231),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_191),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_117),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_209),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_210),
.B(n_228),
.Y(n_252)
);

A2O1A1O1Ixp25_ASAP7_75t_L g259 ( 
.A1(n_212),
.A2(n_181),
.B(n_197),
.C(n_194),
.D(n_193),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_168),
.A2(n_145),
.B1(n_137),
.B2(n_128),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_168),
.A2(n_120),
.B1(n_156),
.B2(n_142),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_126),
.B1(n_136),
.B2(n_99),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_215),
.A2(n_176),
.B1(n_188),
.B2(n_184),
.Y(n_268)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

CKINVDCx11_ASAP7_75t_R g217 ( 
.A(n_190),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_226),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_219),
.C(n_221),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_143),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_220),
.A2(n_178),
.B1(n_194),
.B2(n_193),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_146),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_179),
.A2(n_99),
.B1(n_89),
.B2(n_38),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_222),
.A2(n_223),
.B1(n_187),
.B2(n_176),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_171),
.A2(n_89),
.B1(n_38),
.B2(n_32),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_172),
.A2(n_32),
.B(n_24),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_187),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_32),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_230),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_162),
.B(n_44),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_162),
.B(n_24),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_24),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_163),
.B(n_23),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_233),
.Y(n_254)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_169),
.Y(n_234)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_163),
.B(n_1),
.C(n_2),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_181),
.C(n_178),
.Y(n_265)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_165),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_253),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_229),
.A2(n_159),
.B1(n_196),
.B2(n_161),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_250),
.A2(n_268),
.B1(n_227),
.B2(n_177),
.Y(n_293)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_251),
.Y(n_279)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_199),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_256),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_201),
.B(n_195),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_218),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_225),
.B(n_224),
.Y(n_290)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_199),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_266),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_206),
.B(n_195),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_264),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_221),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_205),
.B(n_184),
.Y(n_266)
);

OAI32xp33_ASAP7_75t_L g267 ( 
.A1(n_202),
.A2(n_229),
.A3(n_233),
.B1(n_230),
.B2(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_231),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_202),
.A2(n_183),
.B1(n_182),
.B2(n_169),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_207),
.B1(n_211),
.B2(n_222),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_274),
.B(n_284),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_266),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_286),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_245),
.A2(n_203),
.B1(n_204),
.B2(n_225),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_276),
.A2(n_293),
.B1(n_301),
.B2(n_242),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_228),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_212),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_281),
.A2(n_288),
.B(n_297),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_285),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_237),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_219),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_294),
.C(n_258),
.Y(n_303)
);

OA21x2_ASAP7_75t_L g288 ( 
.A1(n_239),
.A2(n_211),
.B(n_213),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_289),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_290),
.B(n_295),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_231),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_241),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_255),
.Y(n_308)
);

A2O1A1O1Ixp25_ASAP7_75t_L g297 ( 
.A1(n_242),
.A2(n_235),
.B(n_217),
.C(n_209),
.D(n_223),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_244),
.A2(n_209),
.B(n_177),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_252),
.B(n_227),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_299),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_239),
.A2(n_235),
.B1(n_183),
.B2(n_182),
.Y(n_300)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_300),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_257),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_302),
.A2(n_309),
.B1(n_321),
.B2(n_289),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_311),
.C(n_312),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_246),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_310),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_319),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_288),
.A2(n_262),
.B1(n_257),
.B2(n_260),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_246),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_265),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_274),
.B(n_254),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_291),
.B1(n_278),
.B2(n_283),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_254),
.C(n_269),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_317),
.C(n_324),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_267),
.C(n_248),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_292),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_271),
.B1(n_261),
.B2(n_251),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_272),
.Y(n_323)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_323),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_240),
.C(n_270),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_325),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_280),
.B(n_296),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_340),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_329),
.A2(n_336),
.B1(n_337),
.B2(n_339),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_283),
.Y(n_330)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_330),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_321),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_333),
.B(n_345),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_322),
.A2(n_304),
.B1(n_291),
.B2(n_280),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_304),
.A2(n_278),
.B1(n_277),
.B2(n_290),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_318),
.Y(n_338)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_338),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_317),
.A2(n_277),
.B1(n_282),
.B2(n_271),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_341),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_273),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_344),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_299),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_307),
.A2(n_299),
.B1(n_297),
.B2(n_301),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_302),
.A2(n_298),
.B1(n_240),
.B2(n_247),
.Y(n_346)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_315),
.A2(n_247),
.B(n_270),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_347),
.B(n_307),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_324),
.A2(n_253),
.B1(n_3),
.B2(n_4),
.Y(n_348)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_348),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_328),
.B(n_313),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_354),
.Y(n_366)
);

NOR3xp33_ASAP7_75t_SL g353 ( 
.A(n_330),
.B(n_306),
.C(n_311),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_353),
.A2(n_335),
.B1(n_6),
.B2(n_7),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_312),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_310),
.C(n_313),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_355),
.B(n_356),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_343),
.B(n_316),
.C(n_320),
.Y(n_356)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_360),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_2),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_362),
.C(n_348),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_4),
.C(n_5),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_369),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_356),
.A2(n_339),
.B(n_331),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_5),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_332),
.C(n_347),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_362),
.A2(n_337),
.B(n_349),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_370),
.A2(n_6),
.B(n_8),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_359),
.A2(n_340),
.B1(n_346),
.B2(n_332),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_372),
.B(n_6),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_336),
.C(n_327),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_374),
.Y(n_385)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_357),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_363),
.A2(n_329),
.B1(n_345),
.B2(n_334),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_375),
.B(n_379),
.Y(n_390)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_351),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_361),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_378),
.A2(n_365),
.B1(n_353),
.B2(n_7),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_5),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_376),
.A2(n_364),
.B(n_355),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_382),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_354),
.C(n_352),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_383),
.B(n_386),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_384),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_5),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_388),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_6),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_367),
.C(n_366),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_8),
.Y(n_400)
);

OAI21xp33_ASAP7_75t_L g392 ( 
.A1(n_385),
.A2(n_372),
.B(n_375),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_391),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_396),
.B(n_9),
.Y(n_406)
);

NOR2x1_ASAP7_75t_SL g397 ( 
.A(n_383),
.B(n_366),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_397),
.A2(n_380),
.B(n_386),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_388),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_399),
.B(n_400),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_401),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_403),
.B(n_406),
.C(n_398),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_390),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_404),
.A2(n_405),
.B(n_407),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_9),
.C(n_11),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_395),
.B(n_9),
.C(n_12),
.Y(n_407)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_410),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_400),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_411),
.B(n_409),
.C(n_408),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_412),
.A2(n_392),
.B1(n_402),
.B2(n_12),
.Y(n_414)
);

AO21x1_ASAP7_75t_L g415 ( 
.A1(n_414),
.A2(n_413),
.B(n_13),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_415),
.B(n_13),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_13),
.Y(n_417)
);


endmodule