module fake_aes_5048_n_15 (n_1, n_2, n_4, n_3, n_5, n_0, n_15);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_9;
wire n_14;
wire n_10;
wire n_7;
wire n_8;
INVx2_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
NAND2xp5_ASAP7_75t_SL g7 ( .A(n_0), .B(n_2), .Y(n_7) );
OR2x6_ASAP7_75t_L g8 ( .A(n_5), .B(n_1), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_0), .B(n_3), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
INVxp67_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
NOR4xp25_ASAP7_75t_L g14 ( .A(n_13), .B(n_7), .C(n_11), .D(n_8), .Y(n_14) );
INVx2_ASAP7_75t_SL g15 ( .A(n_14), .Y(n_15) );
endmodule