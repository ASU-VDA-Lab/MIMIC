module real_jpeg_25395_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_176;
wire n_166;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_1),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_2),
.B(n_70),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_2),
.A2(n_35),
.B(n_54),
.C(n_150),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_2),
.B(n_39),
.C(n_92),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_2),
.A2(n_30),
.B1(n_51),
.B2(n_52),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_2),
.A2(n_82),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_2),
.B(n_63),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_4),
.A2(n_51),
.B1(n_52),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_4),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_88),
.Y(n_126)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_6),
.A2(n_27),
.B1(n_35),
.B2(n_59),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_59),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_59),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_45),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_9),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_27),
.B1(n_35),
.B2(n_62),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_10),
.A2(n_62),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_62),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_62),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_11),
.A2(n_32),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_11),
.A2(n_27),
.B1(n_35),
.B2(n_67),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_67),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_67),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_15),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_36)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_15),
.Y(n_129)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_15),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_15),
.A2(n_37),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_15),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_111),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_78),
.B1(n_79),
.B2(n_110),
.Y(n_20)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_21),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_48),
.CI(n_64),
.CON(n_21),
.SN(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_23),
.A2(n_24),
.B1(n_36),
.B2(n_118),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_33),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_25),
.A2(n_26),
.B1(n_74),
.B2(n_75),
.Y(n_77)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_34),
.C(n_35),
.Y(n_33)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_27),
.A2(n_35),
.B1(n_54),
.B2(n_55),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_29),
.A2(n_30),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_30),
.A2(n_51),
.B(n_55),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_30),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_30),
.B(n_95),
.Y(n_192)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_36),
.Y(n_118)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_37),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_38),
.A2(n_39),
.B1(n_92),
.B2(n_94),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_38),
.B(n_183),
.Y(n_182)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_42),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_81)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_42),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_44),
.A2(n_82),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_57),
.B(n_60),
.Y(n_48)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_49),
.A2(n_60),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_50),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_52),
.B1(n_92),
.B2(n_94),
.Y(n_91)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_52),
.B(n_171),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_58),
.A2(n_63),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_104),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B(n_71),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_106),
.B(n_109),
.Y(n_105)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_97),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_82),
.A2(n_179),
.B(n_187),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_95),
.B2(n_96),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_95),
.B(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_89),
.A2(n_143),
.B(n_145),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_89),
.A2(n_145),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_90),
.A2(n_144),
.B1(n_146),
.B2(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

BUFx24_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_95),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_95),
.A2(n_100),
.B(n_160),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.C(n_105),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_101),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_119),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_112),
.A2(n_113),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_125),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_212),
.B(n_218),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_164),
.B(n_211),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_156),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_135),
.B(n_156),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_140),
.B2(n_155),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_136),
.B(n_142),
.C(n_147),
.Y(n_217)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_147),
.B2(n_148),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_149),
.B(n_151),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_153),
.A2(n_177),
.B(n_189),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.C(n_161),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_158),
.A2(n_161),
.B1(n_162),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_205),
.B(n_210),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_195),
.B(n_204),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_180),
.B(n_194),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_175),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_190),
.B(n_193),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_192),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_203),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_202),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_209)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_209),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_217),
.Y(n_218)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);


endmodule