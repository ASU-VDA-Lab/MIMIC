module fake_jpeg_24366_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_2),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_2),
.B(n_1),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_15),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_11),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_20),
.B(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_5),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_11),
.A2(n_6),
.B1(n_12),
.B2(n_7),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_23),
.B(n_17),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_11),
.B1(n_7),
.B2(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_14),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_31),
.B1(n_26),
.B2(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_15),
.Y(n_30)
);

AOI21x1_ASAP7_75t_SL g31 ( 
.A1(n_21),
.A2(n_20),
.B(n_14),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_18),
.B(n_24),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_14),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_10),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_38),
.C(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_10),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_33),
.B(n_9),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.C(n_27),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_8),
.B(n_19),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.C(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_45),
.B(n_19),
.Y(n_46)
);


endmodule