module real_jpeg_11226_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_1),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_2),
.A2(n_32),
.B(n_39),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_2),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_2),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_22),
.Y(n_21)
);

A2O1A1O1Ixp25_ASAP7_75t_L g57 ( 
.A1(n_8),
.A2(n_21),
.B(n_22),
.C(n_58),
.D(n_60),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_8),
.B(n_75),
.Y(n_74)
);

A2O1A1O1Ixp25_ASAP7_75t_L g92 ( 
.A1(n_8),
.A2(n_30),
.B(n_49),
.C(n_85),
.D(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_8),
.B(n_59),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_8),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g126 ( 
.A1(n_8),
.A2(n_40),
.B(n_108),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_43),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_9),
.A2(n_26),
.B1(n_30),
.B2(n_43),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_10),
.A2(n_26),
.B1(n_30),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_55),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_11),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_12),
.A2(n_26),
.B1(n_30),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_12),
.A2(n_22),
.B1(n_23),
.B2(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_47),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_88),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_87),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_63),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_17),
.B(n_63),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_44),
.C(n_57),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_18),
.A2(n_19),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_31),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_24),
.B1(n_27),
.B2(n_30),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_29),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_23),
.A2(n_28),
.B(n_29),
.C(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_26),
.A2(n_50),
.B(n_52),
.C(n_53),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_50),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_33),
.A2(n_40),
.B1(n_41),
.B2(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_35),
.B1(n_50),
.B2(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_34),
.B(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_34),
.B(n_128),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_35),
.A2(n_52),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_39),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_42),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_40),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_40),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_41),
.A2(n_114),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_41),
.B(n_122),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_44),
.A2(n_45),
.B1(n_57),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_54),
.B2(n_56),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_46),
.A2(n_56),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_48),
.A2(n_54),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_49),
.B(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_53),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_56),
.B(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_57),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_67),
.B(n_68),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_81),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_70),
.B2(n_80),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_71),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_74),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_132),
.B(n_138),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_110),
.B(n_131),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_98),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_98),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_92),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_93),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_106),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_103),
.C(n_106),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_119),
.B(n_130),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_117),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_125),
.B(n_129),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_133),
.B(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);


endmodule