module fake_jpeg_15905_n_212 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_212);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_49),
.B(n_56),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_27),
.B1(n_24),
.B2(n_23),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_51),
.B1(n_67),
.B2(n_73),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_27),
.B1(n_24),
.B2(n_33),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_26),
.B1(n_20),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_48),
.B1(n_42),
.B2(n_32),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_1),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_54),
.A2(n_57),
.B1(n_63),
.B2(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_34),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_28),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_62),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_1),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_22),
.B1(n_29),
.B2(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_74),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_21),
.B1(n_32),
.B2(n_17),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_86),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_63),
.B1(n_64),
.B2(n_61),
.Y(n_107)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_17),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_80),
.B(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_35),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_48),
.C(n_39),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_94),
.B1(n_103),
.B2(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_31),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_11),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_88),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_9),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_39),
.C(n_35),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_57),
.A2(n_32),
.B1(n_2),
.B2(n_3),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_101),
.B1(n_79),
.B2(n_66),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_74),
.Y(n_126)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_42),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_71),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_74),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_58),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_63),
.B(n_70),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_105),
.A2(n_108),
.B(n_114),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_111),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_113),
.B1(n_94),
.B2(n_102),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_53),
.B(n_59),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_64),
.B1(n_61),
.B2(n_53),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_53),
.B(n_6),
.Y(n_114)
);

BUFx24_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_77),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_74),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_78),
.B(n_12),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_78),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_134),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_132),
.B1(n_117),
.B2(n_122),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_76),
.B1(n_93),
.B2(n_101),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_135),
.B1(n_144),
.B2(n_107),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_75),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_105),
.A2(n_97),
.B1(n_84),
.B2(n_96),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_114),
.A2(n_72),
.B1(n_100),
.B2(n_88),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_106),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_123),
.B(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_143),
.B(n_125),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_152),
.Y(n_175)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_158),
.B1(n_132),
.B2(n_128),
.C(n_115),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_112),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_153),
.B(n_159),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_110),
.C(n_116),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_163),
.C(n_135),
.Y(n_167)
);

XOR2x2_ASAP7_75t_SL g168 ( 
.A(n_157),
.B(n_146),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_111),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_161),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_117),
.B1(n_122),
.B2(n_92),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_115),
.C(n_9),
.Y(n_163)
);

AO221x1_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_148),
.B1(n_137),
.B2(n_147),
.C(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_171),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_SL g179 ( 
.A(n_168),
.B(n_172),
.C(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_146),
.C(n_140),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_128),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_156),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_132),
.A3(n_130),
.B1(n_133),
.B2(n_139),
.C1(n_127),
.C2(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_5),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_177),
.A2(n_176),
.B1(n_171),
.B2(n_173),
.Y(n_183)
);

OA21x2_ASAP7_75t_SL g190 ( 
.A1(n_179),
.A2(n_180),
.B(n_182),
.Y(n_190)
);

AO22x2_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_161),
.B1(n_150),
.B2(n_164),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_180),
.A2(n_182),
.B1(n_169),
.B2(n_6),
.Y(n_194)
);

AOI22x1_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_154),
.B1(n_164),
.B2(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_163),
.C(n_115),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_185),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_174),
.B(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_190),
.A2(n_180),
.B1(n_179),
.B2(n_185),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_173),
.B(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_195),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_5),
.Y(n_201)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_199),
.C(n_191),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_181),
.C(n_184),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_201),
.B(n_194),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_193),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_203),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_204),
.A2(n_196),
.B(n_200),
.C(n_199),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_188),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_205),
.A2(n_8),
.B(n_14),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_207),
.A2(n_208),
.B(n_15),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_210),
.C(n_7),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_SL g210 ( 
.A(n_206),
.B(n_14),
.C(n_7),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_7),
.Y(n_212)
);


endmodule