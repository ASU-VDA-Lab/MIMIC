module fake_jpeg_20674_n_162 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_162);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_0),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_28),
.Y(n_58)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_45),
.B(n_58),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_27),
.B1(n_25),
.B2(n_21),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_56),
.B1(n_62),
.B2(n_27),
.Y(n_67)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_57),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_61),
.B(n_20),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_26),
.B1(n_23),
.B2(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_70),
.Y(n_95)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_16),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_5),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_72),
.B(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_17),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_25),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_74),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_80),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_42),
.B1(n_21),
.B2(n_22),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_79),
.B1(n_59),
.B2(n_57),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_22),
.B1(n_39),
.B2(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_20),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_39),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_84),
.B(n_53),
.Y(n_91)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_20),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_2),
.C(n_3),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_88),
.C(n_54),
.Y(n_93)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_87),
.A2(n_59),
.B1(n_61),
.B2(n_43),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_2),
.C(n_3),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_103),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_43),
.C(n_48),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_88),
.C(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_63),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_47),
.B1(n_8),
.B2(n_11),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_86),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_47),
.B1(n_11),
.B2(n_12),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_108),
.B1(n_98),
.B2(n_94),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_69),
.A2(n_7),
.B1(n_12),
.B2(n_14),
.Y(n_108)
);

NOR4xp25_ASAP7_75t_SL g109 ( 
.A(n_74),
.B(n_7),
.C(n_79),
.D(n_82),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_98),
.B(n_81),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_112),
.B(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_107),
.B(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_113),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_82),
.B(n_75),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_70),
.C(n_75),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_105),
.B1(n_92),
.B2(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_77),
.Y(n_121)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_93),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_118),
.B(n_120),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_91),
.B(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

OAI321xp33_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_119),
.A3(n_117),
.B1(n_109),
.B2(n_114),
.C(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_138),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_115),
.B1(n_122),
.B2(n_90),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_87),
.B1(n_96),
.B2(n_83),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_140),
.A2(n_100),
.B(n_96),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_77),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_142),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_97),
.C(n_100),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_132),
.C(n_134),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_143),
.A2(n_134),
.B1(n_132),
.B2(n_128),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_147),
.C(n_143),
.Y(n_153)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_125),
.B(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_146),
.B(n_142),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_138),
.B(n_141),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_144),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_151),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_153),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_155),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

NAND2x1_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_145),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_96),
.A3(n_149),
.B1(n_150),
.B2(n_155),
.C1(n_157),
.C2(n_156),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_159),
.B(n_158),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_161),
.Y(n_162)
);


endmodule