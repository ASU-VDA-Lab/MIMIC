module fake_netlist_1_3138_n_727 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_727);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_727;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_311;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_386;
wire n_432;
wire n_659;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_580;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_565;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_573;
wire n_673;
wire n_669;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_409;
wire n_315;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_615;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_535;
wire n_530;
wire n_358;
wire n_267;
wire n_456;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_602;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_538;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_695;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_709;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g240 ( .A(n_120), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_163), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_226), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_217), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_47), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_56), .Y(n_245) );
BUFx10_ASAP7_75t_L g246 ( .A(n_80), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_206), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_223), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_10), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_156), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_98), .Y(n_251) );
INVxp67_ASAP7_75t_L g252 ( .A(n_2), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_131), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_201), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_85), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_110), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_216), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_205), .Y(n_258) );
INVxp67_ASAP7_75t_L g259 ( .A(n_0), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_185), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_86), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_237), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_49), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_29), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_60), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_220), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_160), .B(n_155), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_8), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_25), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_171), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_41), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_200), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_97), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_221), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_104), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_197), .Y(n_276) );
CKINVDCx16_ASAP7_75t_R g277 ( .A(n_10), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_51), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_3), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_184), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_5), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_37), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_67), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_126), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_194), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_88), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_239), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_207), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_84), .B(n_121), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_174), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_218), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_202), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_1), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_118), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_142), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_212), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_152), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_159), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_219), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_11), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_170), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_213), .Y(n_302) );
CKINVDCx14_ASAP7_75t_R g303 ( .A(n_35), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_108), .Y(n_304) );
CKINVDCx11_ASAP7_75t_R g305 ( .A(n_78), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_25), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_95), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_129), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_134), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_224), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_111), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_54), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_187), .Y(n_313) );
CKINVDCx14_ASAP7_75t_R g314 ( .A(n_232), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_69), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_193), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_234), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_113), .Y(n_318) );
CKINVDCx16_ASAP7_75t_R g319 ( .A(n_208), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_132), .Y(n_320) );
NOR2xp67_ASAP7_75t_L g321 ( .A(n_145), .B(n_122), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_119), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_71), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_96), .Y(n_324) );
CKINVDCx16_ASAP7_75t_R g325 ( .A(n_76), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_178), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_1), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_222), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_137), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_94), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_157), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_161), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_9), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_141), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_229), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_87), .Y(n_336) );
INVxp33_ASAP7_75t_L g337 ( .A(n_189), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_91), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_17), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_183), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_167), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_101), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_106), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_68), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_148), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_19), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_20), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_265), .Y(n_348) );
OA21x2_ASAP7_75t_L g349 ( .A1(n_241), .A2(n_27), .B(n_26), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_240), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_243), .Y(n_351) );
INVx4_ASAP7_75t_L g352 ( .A(n_283), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_265), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_247), .A2(n_30), .B(n_28), .Y(n_354) );
NAND2xp33_ASAP7_75t_L g355 ( .A(n_244), .B(n_31), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_333), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_264), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_334), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_277), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_249), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_240), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_252), .Y(n_362) );
OA21x2_ASAP7_75t_L g363 ( .A1(n_242), .A2(n_33), .B(n_32), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_278), .A2(n_36), .B(n_34), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_268), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_252), .A2(n_3), .B1(n_0), .B2(n_2), .Y(n_366) );
BUFx8_ASAP7_75t_SL g367 ( .A(n_346), .Y(n_367) );
NOR2x1_ASAP7_75t_L g368 ( .A(n_269), .B(n_38), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_356), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_351), .Y(n_370) );
INVx2_ASAP7_75t_SL g371 ( .A(n_352), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_350), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_352), .B(n_337), .Y(n_373) );
CKINVDCx16_ASAP7_75t_R g374 ( .A(n_359), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_362), .B(n_259), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_365), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_348), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_354), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_359), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_364), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_353), .B(n_285), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_350), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_357), .B(n_331), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_360), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_370), .Y(n_385) );
NOR3xp33_ASAP7_75t_L g386 ( .A(n_374), .B(n_366), .C(n_325), .Y(n_386) );
INVx5_ASAP7_75t_L g387 ( .A(n_376), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_373), .B(n_358), .Y(n_388) );
O2A1O1Ixp5_ASAP7_75t_L g389 ( .A1(n_378), .A2(n_251), .B(n_254), .C(n_253), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_377), .B(n_355), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_373), .B(n_319), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_384), .A2(n_355), .B1(n_281), .B2(n_306), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_375), .B(n_259), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_371), .B(n_279), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_381), .B(n_368), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_369), .Y(n_396) );
BUFx6f_ASAP7_75t_SL g397 ( .A(n_379), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_383), .B(n_303), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_383), .A2(n_327), .B1(n_339), .B2(n_300), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_379), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_380), .Y(n_401) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_382), .A2(n_280), .B(n_256), .C(n_257), .Y(n_402) );
INVx8_ASAP7_75t_L g403 ( .A(n_372), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_372), .A2(n_314), .B1(n_305), .B2(n_255), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_401), .A2(n_363), .B(n_349), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_390), .A2(n_363), .B(n_349), .Y(n_406) );
O2A1O1Ixp5_ASAP7_75t_L g407 ( .A1(n_389), .A2(n_343), .B(n_345), .C(n_267), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_390), .A2(n_363), .B(n_349), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_388), .B(n_367), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_397), .A2(n_263), .B1(n_273), .B2(n_271), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_393), .B(n_293), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_392), .A2(n_294), .B1(n_304), .B2(n_280), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_398), .B(n_347), .Y(n_413) );
NOR2xp67_ASAP7_75t_L g414 ( .A(n_400), .B(n_4), .Y(n_414) );
O2A1O1Ixp33_ASAP7_75t_L g415 ( .A1(n_386), .A2(n_258), .B(n_270), .C(n_262), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_395), .A2(n_274), .B(n_272), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_395), .A2(n_276), .B(n_275), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_391), .B(n_367), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_387), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_385), .Y(n_420) );
O2A1O1Ixp33_ASAP7_75t_L g421 ( .A1(n_396), .A2(n_288), .B(n_290), .C(n_284), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_387), .B(n_248), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_394), .B(n_250), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_387), .Y(n_424) );
INVx5_ASAP7_75t_L g425 ( .A(n_387), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_397), .B(n_246), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_420), .Y(n_427) );
AO32x2_ASAP7_75t_L g428 ( .A1(n_412), .A2(n_399), .A3(n_402), .B1(n_404), .B2(n_350), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_406), .A2(n_403), .B(n_289), .Y(n_429) );
AOI21x1_ASAP7_75t_L g430 ( .A1(n_405), .A2(n_321), .B(n_301), .Y(n_430) );
INVx5_ASAP7_75t_L g431 ( .A(n_419), .Y(n_431) );
OR2x6_ASAP7_75t_L g432 ( .A(n_415), .B(n_403), .Y(n_432) );
AO32x2_ASAP7_75t_L g433 ( .A1(n_421), .A2(n_361), .A3(n_350), .B1(n_246), .B2(n_7), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_416), .A2(n_302), .B(n_310), .C(n_291), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_414), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_409), .A2(n_317), .B1(n_322), .B2(n_313), .C(n_312), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_411), .B(n_403), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_413), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_419), .Y(n_439) );
OR2x6_ASAP7_75t_L g440 ( .A(n_418), .B(n_324), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_408), .A2(n_328), .B(n_326), .Y(n_441) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_407), .A2(n_335), .B(n_330), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_417), .B(n_340), .Y(n_443) );
NOR3xp33_ASAP7_75t_L g444 ( .A(n_410), .B(n_344), .C(n_260), .Y(n_444) );
AO31x2_ASAP7_75t_L g445 ( .A1(n_424), .A2(n_361), .A3(n_298), .B(n_245), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_425), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_423), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_422), .A2(n_266), .B(n_261), .Y(n_448) );
OAI21x1_ASAP7_75t_L g449 ( .A1(n_425), .A2(n_298), .B(n_245), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_426), .Y(n_450) );
AO31x2_ASAP7_75t_L g451 ( .A1(n_425), .A2(n_361), .A3(n_298), .B(n_342), .Y(n_451) );
OAI21x1_ASAP7_75t_L g452 ( .A1(n_405), .A2(n_40), .B(n_39), .Y(n_452) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_430), .A2(n_361), .B(n_307), .Y(n_453) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_429), .A2(n_286), .B(n_282), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_427), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_441), .A2(n_292), .B(n_287), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_431), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_447), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_444), .B(n_6), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_431), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_436), .B(n_7), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_440), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_446), .B(n_437), .Y(n_463) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_452), .A2(n_296), .B(n_295), .Y(n_464) );
INVxp67_ASAP7_75t_L g465 ( .A(n_440), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_442), .A2(n_299), .B(n_297), .Y(n_466) );
AO31x2_ASAP7_75t_L g467 ( .A1(n_434), .A2(n_443), .A3(n_435), .B(n_439), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_432), .Y(n_468) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_449), .A2(n_309), .B(n_308), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_432), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_433), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_450), .Y(n_472) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_445), .A2(n_315), .B(n_311), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_445), .Y(n_474) );
OAI21x1_ASAP7_75t_L g475 ( .A1(n_448), .A2(n_43), .B(n_42), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_428), .Y(n_476) );
OAI21x1_ASAP7_75t_L g477 ( .A1(n_451), .A2(n_45), .B(n_44), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_428), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_431), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_438), .B(n_12), .Y(n_480) );
OAI21x1_ASAP7_75t_L g481 ( .A1(n_452), .A2(n_48), .B(n_46), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_438), .A2(n_318), .B1(n_320), .B2(n_316), .Y(n_482) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_430), .A2(n_329), .B(n_323), .Y(n_483) );
OAI21x1_ASAP7_75t_SL g484 ( .A1(n_439), .A2(n_13), .B(n_14), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_440), .B(n_332), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_429), .A2(n_338), .B(n_336), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_429), .A2(n_341), .B(n_52), .Y(n_487) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_430), .A2(n_53), .B(n_50), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_455), .Y(n_489) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_474), .A2(n_15), .B(n_16), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g491 ( .A1(n_461), .A2(n_15), .B1(n_16), .B2(n_17), .C(n_18), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_460), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_471), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_480), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_465), .B(n_472), .Y(n_495) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_474), .A2(n_21), .B(n_22), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_462), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_459), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_471), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_463), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_487), .A2(n_23), .B(n_24), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_479), .B(n_24), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_463), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_457), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_467), .B(n_55), .Y(n_505) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_453), .A2(n_57), .B(n_58), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_467), .B(n_59), .Y(n_507) );
INVxp67_ASAP7_75t_SL g508 ( .A(n_478), .Y(n_508) );
OR2x6_ASAP7_75t_L g509 ( .A(n_468), .B(n_61), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_470), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_485), .B(n_238), .Y(n_511) );
INVx3_ASAP7_75t_L g512 ( .A(n_467), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_484), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_482), .B(n_62), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_475), .B(n_63), .Y(n_515) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_476), .A2(n_64), .B(n_65), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_481), .B(n_66), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_483), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_469), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_473), .Y(n_520) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_477), .A2(n_70), .B(n_72), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_473), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_454), .B(n_73), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_469), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_464), .Y(n_525) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_486), .A2(n_74), .B(n_75), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_466), .B(n_77), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_464), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_488), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_456), .B(n_79), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_488), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_471), .A2(n_81), .B(n_82), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_458), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_458), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_474), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_455), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_458), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_458), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_465), .B(n_83), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_455), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_455), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_493), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_498), .B(n_89), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_499), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_509), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_533), .B(n_90), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_535), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_492), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_534), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_537), .B(n_538), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_536), .B(n_236), .Y(n_551) );
NOR2x1_ASAP7_75t_L g552 ( .A(n_509), .B(n_92), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_540), .B(n_93), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_541), .B(n_235), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_489), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_495), .B(n_233), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_502), .B(n_99), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_504), .B(n_500), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_509), .B(n_100), .Y(n_559) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_490), .B(n_102), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_510), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_503), .Y(n_562) );
INVx4_ASAP7_75t_L g563 ( .A(n_517), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_490), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_494), .B(n_231), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_529), .A2(n_103), .B(n_105), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_496), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_539), .B(n_107), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_511), .B(n_109), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_491), .B(n_112), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_514), .B(n_114), .Y(n_572) );
INVx2_ASAP7_75t_SL g573 ( .A(n_497), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_491), .B(n_115), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_513), .B(n_116), .Y(n_575) );
BUFx2_ASAP7_75t_L g576 ( .A(n_523), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_501), .B(n_117), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_501), .B(n_123), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_530), .B(n_230), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_518), .B(n_124), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_527), .B(n_125), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_508), .B(n_127), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_528), .Y(n_583) );
AND2x4_ASAP7_75t_L g584 ( .A(n_525), .B(n_128), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_525), .B(n_228), .Y(n_585) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_515), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_512), .B(n_130), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_512), .B(n_227), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_532), .B(n_133), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_519), .B(n_135), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_524), .Y(n_591) );
NOR2x1p5_ASAP7_75t_L g592 ( .A(n_505), .B(n_136), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_507), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_520), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_520), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_522), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_526), .B(n_138), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_526), .B(n_139), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_516), .Y(n_599) );
BUFx2_ASAP7_75t_L g600 ( .A(n_521), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_506), .B(n_225), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_531), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_549), .B(n_529), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_558), .B(n_506), .Y(n_604) );
INVx3_ASAP7_75t_L g605 ( .A(n_563), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_542), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_548), .B(n_516), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_563), .B(n_140), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_555), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_561), .B(n_143), .Y(n_610) );
BUFx2_ASAP7_75t_SL g611 ( .A(n_573), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_550), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_552), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_545), .B(n_144), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_547), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_562), .B(n_146), .Y(n_616) );
NAND2x1_ASAP7_75t_L g617 ( .A(n_545), .B(n_147), .Y(n_617) );
NAND2x1_ASAP7_75t_L g618 ( .A(n_564), .B(n_149), .Y(n_618) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_586), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_559), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_576), .B(n_150), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_556), .B(n_151), .Y(n_622) );
INVx4_ASAP7_75t_L g623 ( .A(n_559), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_542), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_544), .Y(n_625) );
NAND2x1_ASAP7_75t_SL g626 ( .A(n_575), .B(n_577), .Y(n_626) );
AND2x4_ASAP7_75t_L g627 ( .A(n_586), .B(n_153), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_583), .B(n_154), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_543), .B(n_158), .Y(n_629) );
BUFx2_ASAP7_75t_L g630 ( .A(n_586), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_557), .B(n_162), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_594), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_582), .Y(n_633) );
INVx2_ASAP7_75t_SL g634 ( .A(n_551), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_565), .B(n_164), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_595), .B(n_165), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_575), .Y(n_637) );
AND2x4_ASAP7_75t_L g638 ( .A(n_595), .B(n_166), .Y(n_638) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_590), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_596), .Y(n_640) );
BUFx2_ASAP7_75t_L g641 ( .A(n_590), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_591), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_570), .B(n_168), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_602), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_602), .B(n_169), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_568), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_584), .Y(n_647) );
INVx4_ASAP7_75t_L g648 ( .A(n_572), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_566), .B(n_172), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_620), .Y(n_650) );
INVx2_ASAP7_75t_SL g651 ( .A(n_605), .Y(n_651) );
NAND2x1p5_ASAP7_75t_L g652 ( .A(n_623), .B(n_569), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_644), .Y(n_653) );
BUFx2_ASAP7_75t_L g654 ( .A(n_623), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_615), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_612), .B(n_593), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_609), .B(n_593), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_632), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_605), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_640), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_606), .B(n_560), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_641), .A2(n_592), .B1(n_580), .B2(n_578), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_606), .Y(n_663) );
NAND2x1_ASAP7_75t_SL g664 ( .A(n_648), .B(n_584), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_604), .B(n_600), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_624), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_633), .B(n_639), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_603), .B(n_553), .Y(n_668) );
NAND4xp25_ASAP7_75t_SL g669 ( .A(n_611), .B(n_574), .C(n_571), .D(n_581), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_648), .B(n_579), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_637), .B(n_587), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_642), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_630), .B(n_588), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_625), .B(n_585), .Y(n_674) );
NOR2xp67_ASAP7_75t_L g675 ( .A(n_613), .B(n_599), .Y(n_675) );
NOR2xp67_ASAP7_75t_L g676 ( .A(n_647), .B(n_597), .Y(n_676) );
INVxp67_ASAP7_75t_SL g677 ( .A(n_653), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_669), .A2(n_634), .B1(n_647), .B2(n_621), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_655), .Y(n_679) );
INVx2_ASAP7_75t_SL g680 ( .A(n_654), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_672), .B(n_646), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_667), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_658), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_650), .B(n_607), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_659), .B(n_608), .Y(n_685) );
AND3x2_ASAP7_75t_L g686 ( .A(n_670), .B(n_608), .C(n_614), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_660), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_663), .Y(n_688) );
INVx2_ASAP7_75t_SL g689 ( .A(n_651), .Y(n_689) );
INVx1_ASAP7_75t_SL g690 ( .A(n_659), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_666), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_656), .B(n_635), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_657), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_678), .A2(n_662), .B1(n_676), .B2(n_671), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_680), .A2(n_664), .B(n_626), .C(n_676), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_689), .A2(n_692), .B1(n_677), .B2(n_662), .C(n_652), .Y(n_696) );
A2O1A1Ixp33_ASAP7_75t_L g697 ( .A1(n_682), .A2(n_622), .B(n_617), .C(n_675), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_693), .B(n_665), .Y(n_698) );
AOI21xp33_ASAP7_75t_SL g699 ( .A1(n_685), .A2(n_614), .B(n_628), .Y(n_699) );
AOI21xp33_ASAP7_75t_SL g700 ( .A1(n_686), .A2(n_636), .B(n_643), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_690), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g702 ( .A1(n_692), .A2(n_675), .B1(n_668), .B2(n_618), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_684), .A2(n_673), .B1(n_674), .B2(n_661), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_695), .A2(n_681), .B(n_679), .Y(n_704) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_694), .A2(n_683), .B(n_681), .Y(n_705) );
AOI31xp33_ASAP7_75t_L g706 ( .A1(n_700), .A2(n_631), .A3(n_610), .B(n_649), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_694), .A2(n_697), .B1(n_703), .B2(n_699), .Y(n_707) );
OAI22xp5_ASAP7_75t_SL g708 ( .A1(n_701), .A2(n_645), .B1(n_638), .B2(n_627), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_702), .A2(n_691), .B1(n_688), .B2(n_687), .Y(n_709) );
OAI322xp33_ASAP7_75t_L g710 ( .A1(n_698), .A2(n_546), .A3(n_616), .B1(n_629), .B2(n_589), .C1(n_601), .C2(n_554), .Y(n_710) );
NAND3xp33_ASAP7_75t_SL g711 ( .A(n_700), .B(n_567), .C(n_598), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_696), .A2(n_619), .B1(n_175), .B2(n_176), .Y(n_712) );
AOI211xp5_ASAP7_75t_L g713 ( .A1(n_700), .A2(n_173), .B(n_177), .C(n_179), .Y(n_713) );
AOI211xp5_ASAP7_75t_L g714 ( .A1(n_700), .A2(n_180), .B(n_181), .C(n_182), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_711), .B(n_707), .C(n_712), .Y(n_715) );
NAND3xp33_ASAP7_75t_L g716 ( .A(n_705), .B(n_709), .C(n_714), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_706), .A2(n_704), .B(n_708), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g718 ( .A(n_715), .B(n_713), .C(n_710), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_716), .A2(n_186), .B1(n_188), .B2(n_190), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g720 ( .A(n_718), .B(n_717), .C(n_191), .D(n_192), .Y(n_720) );
OAI21x1_ASAP7_75t_SL g721 ( .A1(n_720), .A2(n_719), .B(n_196), .Y(n_721) );
AOI21x1_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_195), .B(n_198), .Y(n_722) );
AND2x4_ASAP7_75t_L g723 ( .A(n_722), .B(n_199), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_723), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_724), .A2(n_203), .B(n_204), .Y(n_725) );
OA21x2_ASAP7_75t_L g726 ( .A1(n_725), .A2(n_209), .B(n_210), .Y(n_726) );
AOI22xp5_ASAP7_75t_SL g727 ( .A1(n_726), .A2(n_211), .B1(n_214), .B2(n_215), .Y(n_727) );
endmodule