module fake_jpeg_29120_n_88 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_88);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_88;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx3_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_21),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_17),
.Y(n_28)
);

CKINVDCx9p33_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_23),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_15),
.B1(n_21),
.B2(n_11),
.Y(n_37)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_12),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_18),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_38),
.B1(n_20),
.B2(n_18),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_20),
.B1(n_21),
.B2(n_19),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_42),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_26),
.B1(n_22),
.B2(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_22),
.B1(n_11),
.B2(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_12),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_14),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_45),
.C(n_47),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_52),
.C(n_38),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_37),
.C(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_54),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_22),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_46),
.B(n_39),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_46),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_38),
.B1(n_36),
.B2(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_59),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_16),
.C(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_63),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_36),
.B1(n_9),
.B2(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_33),
.B1(n_18),
.B2(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_19),
.B1(n_29),
.B2(n_27),
.Y(n_63)
);

NOR4xp25_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_46),
.C(n_2),
.D(n_3),
.Y(n_66)
);

OA21x2_ASAP7_75t_SL g71 ( 
.A1(n_66),
.A2(n_0),
.B(n_2),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_9),
.B1(n_13),
.B2(n_19),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_63),
.C(n_62),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_72),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_R g72 ( 
.A1(n_68),
.A2(n_56),
.B(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_74),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_68),
.C(n_65),
.Y(n_77)
);

AOI321xp33_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_9),
.A3(n_13),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_79),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_29),
.C(n_27),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_73),
.B(n_67),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_82),
.C(n_19),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_78),
.A3(n_29),
.B1(n_27),
.B2(n_31),
.C1(n_0),
.C2(n_7),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_4),
.B(n_6),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_4),
.C(n_6),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_86),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_4),
.Y(n_88)
);


endmodule