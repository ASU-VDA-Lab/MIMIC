module fake_jpeg_4656_n_232 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_232);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_14),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_16),
.B1(n_15),
.B2(n_26),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_42),
.B1(n_51),
.B2(n_15),
.Y(n_56)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_15),
.B1(n_26),
.B2(n_16),
.Y(n_42)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_26),
.B1(n_16),
.B2(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_53),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_16),
.B1(n_15),
.B2(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_30),
.Y(n_84)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_64),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_20),
.B1(n_37),
.B2(n_22),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_63),
.B1(n_70),
.B2(n_72),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_20),
.B1(n_37),
.B2(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_33),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_20),
.B1(n_22),
.B2(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_36),
.B1(n_33),
.B2(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_40),
.B(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_40),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_43),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_54),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_44),
.B1(n_39),
.B2(n_19),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_38),
.B1(n_51),
.B2(n_44),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_30),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_95),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_19),
.B1(n_27),
.B2(n_21),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_27),
.B1(n_21),
.B2(n_17),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_39),
.B1(n_30),
.B2(n_23),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_71),
.B1(n_68),
.B2(n_66),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_18),
.B1(n_23),
.B2(n_30),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_96),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_43),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_43),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_1),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_100),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_64),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_23),
.B(n_18),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_111),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_63),
.B(n_55),
.C(n_43),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_118),
.B1(n_93),
.B2(n_75),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_43),
.B1(n_66),
.B2(n_59),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_115),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_74),
.C(n_9),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_74),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_59),
.B1(n_14),
.B2(n_8),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_93),
.B(n_75),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_85),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_129),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_96),
.B1(n_88),
.B2(n_84),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_122),
.A2(n_116),
.B1(n_86),
.B2(n_14),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_107),
.B1(n_80),
.B2(n_84),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_136),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_85),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_141),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_110),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_107),
.B1(n_98),
.B2(n_112),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_153),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_104),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_147),
.C(n_148),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_101),
.C(n_109),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_117),
.C(n_105),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_150),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_106),
.B(n_91),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_91),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_137),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_129),
.B1(n_160),
.B2(n_161),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_136),
.B(n_48),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_159),
.B(n_134),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_48),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_120),
.C(n_122),
.Y(n_173)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_156),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_128),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_173),
.A2(n_153),
.B(n_152),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_123),
.C(n_121),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_175),
.C(n_152),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_123),
.C(n_127),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_130),
.B1(n_134),
.B2(n_131),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_142),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_174),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_182),
.B(n_190),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_184),
.C(n_188),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_169),
.B1(n_164),
.B2(n_167),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_150),
.C(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_166),
.B(n_145),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_165),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_192),
.C(n_199),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_175),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_200),
.B(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_181),
.B(n_144),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_179),
.B(n_186),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_163),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_180),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_208),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_206),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_185),
.B(n_178),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_209),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_182),
.C(n_177),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_164),
.B(n_130),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_151),
.B(n_158),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_210),
.B(n_201),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_7),
.A3(n_12),
.B1(n_11),
.B2(n_6),
.C1(n_45),
.C2(n_14),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_203),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_151),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_191),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_214),
.B(n_2),
.Y(n_222)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_193),
.C(n_10),
.Y(n_215)
);

AOI21x1_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_10),
.B(n_12),
.Y(n_218)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_220),
.B(n_221),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_7),
.C(n_3),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_216),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_215),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_222),
.B(n_217),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_224),
.A2(n_45),
.B(n_3),
.Y(n_228)
);

AOI21x1_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_228),
.B(n_226),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_229),
.A2(n_225),
.B(n_3),
.Y(n_230)
);

AOI321xp33_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_218),
.C(n_227),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_2),
.Y(n_232)
);


endmodule