module fake_jpeg_28254_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_25),
.Y(n_30)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_0),
.C(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_20),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_20),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_42),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_52),
.B(n_13),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

FAx1_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_28),
.CI(n_26),
.CON(n_42),
.SN(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_48),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_17),
.B1(n_19),
.B2(n_13),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_25),
.B(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_42),
.B1(n_50),
.B2(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_65),
.B(n_63),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_61),
.C(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_42),
.B1(n_24),
.B2(n_26),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_24),
.B1(n_25),
.B2(n_48),
.Y(n_74)
);

A2O1A1O1Ixp25_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_46),
.B(n_64),
.C(n_16),
.D(n_14),
.Y(n_77)
);

A2O1A1O1Ixp25_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_82),
.B(n_12),
.C(n_22),
.D(n_11),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_75),
.B1(n_58),
.B2(n_60),
.Y(n_87)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_14),
.B(n_12),
.C(n_22),
.D(n_10),
.Y(n_82)
);

XNOR2x1_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_11),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_56),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_69),
.B(n_74),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_88),
.C(n_89),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_79),
.Y(n_89)
);

INVxp67_ASAP7_75t_SL g92 ( 
.A(n_88),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_96),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_78),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_97),
.C(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_90),
.B(n_58),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_4),
.B(n_6),
.C(n_9),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_98),
.B(n_10),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_102),
.Y(n_104)
);


endmodule