module fake_netlist_5_2522_n_358 (n_91, n_82, n_10, n_24, n_86, n_83, n_61, n_90, n_75, n_101, n_65, n_78, n_74, n_57, n_96, n_37, n_108, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_42, n_22, n_1, n_45, n_46, n_21, n_94, n_38, n_105, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_85, n_95, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_28, n_89, n_70, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_358);

input n_91;
input n_82;
input n_10;
input n_24;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_57;
input n_96;
input n_37;
input n_108;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_42;
input n_22;
input n_1;
input n_45;
input n_46;
input n_21;
input n_94;
input n_38;
input n_105;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_85;
input n_95;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_28;
input n_89;
input n_70;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;

output n_358;

wire n_137;
wire n_294;
wire n_318;
wire n_194;
wire n_316;
wire n_248;
wire n_124;
wire n_136;
wire n_146;
wire n_315;
wire n_268;
wire n_127;
wire n_235;
wire n_226;
wire n_353;
wire n_351;
wire n_111;
wire n_155;
wire n_116;
wire n_284;
wire n_245;
wire n_139;
wire n_280;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_244;
wire n_173;
wire n_198;
wire n_247;
wire n_314;
wire n_321;
wire n_292;
wire n_212;
wire n_119;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_147;
wire n_307;
wire n_150;
wire n_209;
wire n_259;
wire n_301;
wire n_186;
wire n_134;
wire n_191;
wire n_171;
wire n_153;
wire n_341;
wire n_204;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_122;
wire n_282;
wire n_331;
wire n_325;
wire n_132;
wire n_281;
wire n_240;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_123;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_267;
wire n_297;
wire n_156;
wire n_225;
wire n_219;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_211;
wire n_218;
wire n_181;
wire n_290;
wire n_221;
wire n_178;
wire n_287;
wire n_344;
wire n_141;
wire n_355;
wire n_336;
wire n_145;
wire n_337;
wire n_313;
wire n_216;
wire n_168;
wire n_164;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_144;
wire n_114;
wire n_165;
wire n_213;
wire n_129;
wire n_342;
wire n_197;
wire n_236;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_277;
wire n_338;
wire n_149;
wire n_333;
wire n_309;
wire n_130;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_112;
wire n_239;
wire n_310;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_118;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_312;
wire n_345;
wire n_210;
wire n_176;
wire n_182;
wire n_143;
wire n_354;
wire n_237;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_229;
wire n_177;
wire n_117;
wire n_326;
wire n_233;
wire n_205;
wire n_113;
wire n_246;
wire n_179;
wire n_125;
wire n_269;
wire n_128;
wire n_285;
wire n_120;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_154;
wire n_148;
wire n_300;
wire n_159;
wire n_334;
wire n_175;
wire n_262;
wire n_238;
wire n_319;
wire n_121;
wire n_242;
wire n_200;
wire n_162;
wire n_222;
wire n_115;
wire n_324;
wire n_199;
wire n_187;
wire n_348;
wire n_166;
wire n_256;
wire n_305;
wire n_278;
wire n_110;

INVxp33_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_38),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_78),
.Y(n_112)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_19),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_5),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_16),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_47),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_17),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_43),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_65),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_14),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_27),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_21),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_25),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_53),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_92),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_4),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_48),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_32),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_35),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_18),
.Y(n_145)
);

INVx4_ASAP7_75t_R g146 ( 
.A(n_87),
.Y(n_146)
);

NOR2xp67_ASAP7_75t_L g147 ( 
.A(n_29),
.B(n_55),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_85),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_46),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_45),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_15),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_36),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_82),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_42),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_61),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_10),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_2),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_111),
.B(n_0),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_51),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_115),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_52),
.B(n_106),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_109),
.B(n_0),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

AND2x4_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_1),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

CKINVDCx6p67_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_2),
.Y(n_174)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g178 ( 
.A(n_110),
.B(n_54),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_109),
.B(n_3),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_179),
.B1(n_163),
.B2(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_112),
.Y(n_182)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_112),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_113),
.Y(n_185)
);

AND2x4_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_113),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_178),
.B(n_151),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_178),
.B(n_151),
.Y(n_191)
);

NAND2xp33_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_133),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_131),
.B1(n_133),
.B2(n_120),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_173),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_119),
.Y(n_201)
);

AO21x2_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_147),
.B(n_131),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

OR2x6_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_121),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_122),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_203),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_116),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_197),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_123),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_128),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_125),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_134),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_139),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_181),
.B(n_161),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_133),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_142),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_148),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_SL g231 ( 
.A(n_196),
.B(n_159),
.C(n_158),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_204),
.B(n_126),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_187),
.A2(n_145),
.B(n_129),
.Y(n_233)
);

OR2x6_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_127),
.Y(n_234)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_149),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_196),
.B(n_156),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_157),
.B(n_155),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

NAND2x1p5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_198),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_202),
.Y(n_245)
);

O2A1O1Ixp5_ASAP7_75t_SL g246 ( 
.A1(n_225),
.A2(n_143),
.B(n_154),
.C(n_153),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_138),
.B1(n_135),
.B2(n_152),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

OAI221xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_150),
.B1(n_136),
.B2(n_137),
.C(n_132),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_221),
.A2(n_146),
.B1(n_183),
.B2(n_202),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_183),
.B(n_133),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_216),
.A2(n_183),
.B1(n_133),
.B2(n_56),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_211),
.A2(n_230),
.B1(n_222),
.B2(n_218),
.Y(n_255)
);

O2A1O1Ixp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_50),
.B(n_103),
.C(n_101),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_212),
.B(n_4),
.Y(n_257)
);

OR2x6_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_6),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_6),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_226),
.A2(n_218),
.B(n_214),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_57),
.B(n_100),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_215),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_7),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

O2A1O1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

AO31x2_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_239),
.A3(n_229),
.B(n_227),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_212),
.Y(n_271)
);

O2A1O1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_232),
.B(n_219),
.C(n_212),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_243),
.A2(n_266),
.B(n_242),
.Y(n_273)
);

AO32x2_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_8),
.A3(n_215),
.B1(n_219),
.B2(n_12),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_235),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

AOI221x1_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_11),
.B1(n_20),
.B2(n_22),
.C(n_23),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_247),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_280)
);

O2A1O1Ixp33_ASAP7_75t_SL g281 ( 
.A1(n_257),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_263),
.A2(n_37),
.B(n_39),
.Y(n_283)
);

AO31x2_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_40),
.A3(n_41),
.B(n_44),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_59),
.B(n_69),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_265),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_258),
.B1(n_262),
.B2(n_241),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_248),
.B1(n_258),
.B2(n_261),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_256),
.B(n_248),
.C(n_246),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_70),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_277),
.B(n_269),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_269),
.B1(n_278),
.B2(n_280),
.Y(n_295)
);

OAI221xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.C(n_76),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_283),
.Y(n_297)
);

OA21x2_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_77),
.B(n_79),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_270),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_270),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_297),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_270),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

OR2x6_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_285),
.Y(n_306)
);

AND2x4_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_284),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_284),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_284),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_274),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_274),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_300),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_309),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_307),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_307),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_313),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_307),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

OAI211xp5_ASAP7_75t_SL g328 ( 
.A1(n_319),
.A2(n_287),
.B(n_296),
.C(n_294),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_298),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_318),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_315),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_315),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_315),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_326),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_330),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_315),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_324),
.Y(n_338)
);

OAI322xp33_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_331),
.A3(n_320),
.B1(n_327),
.B2(n_321),
.C1(n_323),
.C2(n_325),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_329),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_338),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_340),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_334),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_341),
.B(n_336),
.Y(n_344)
);

AOI221xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_339),
.B1(n_342),
.B2(n_328),
.C(n_333),
.Y(n_345)
);

OAI321xp33_ASAP7_75t_L g346 ( 
.A1(n_343),
.A2(n_328),
.A3(n_337),
.B1(n_306),
.B2(n_295),
.C(n_290),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_345),
.B(n_321),
.Y(n_347)
);

NAND4xp25_ASAP7_75t_L g348 ( 
.A(n_346),
.B(n_80),
.C(n_83),
.D(n_84),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_89),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_349),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_350),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_347),
.B1(n_306),
.B2(n_298),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_352),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_352),
.B(n_90),
.Y(n_354)
);

NAND3xp33_ASAP7_75t_L g355 ( 
.A(n_353),
.B(n_298),
.C(n_93),
.Y(n_355)
);

OAI21x1_ASAP7_75t_L g356 ( 
.A1(n_354),
.A2(n_91),
.B(n_94),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_356),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_355),
.B(n_107),
.Y(n_358)
);


endmodule