module fake_aes_7665_n_141 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_141);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_141;
wire n_117;
wire n_44;
wire n_133;
wire n_81;
wire n_69;
wire n_22;
wire n_57;
wire n_88;
wire n_52;
wire n_26;
wire n_50;
wire n_33;
wire n_102;
wire n_73;
wire n_49;
wire n_119;
wire n_115;
wire n_97;
wire n_80;
wire n_107;
wire n_60;
wire n_114;
wire n_121;
wire n_41;
wire n_35;
wire n_94;
wire n_65;
wire n_125;
wire n_130;
wire n_103;
wire n_19;
wire n_87;
wire n_137;
wire n_104;
wire n_98;
wire n_74;
wire n_29;
wire n_45;
wire n_85;
wire n_101;
wire n_62;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_23;
wire n_91;
wire n_108;
wire n_116;
wire n_139;
wire n_16;
wire n_113;
wire n_95;
wire n_124;
wire n_128;
wire n_129;
wire n_120;
wire n_70;
wire n_17;
wire n_63;
wire n_71;
wire n_90;
wire n_56;
wire n_135;
wire n_42;
wire n_24;
wire n_78;
wire n_127;
wire n_40;
wire n_111;
wire n_79;
wire n_38;
wire n_64;
wire n_46;
wire n_31;
wire n_58;
wire n_122;
wire n_138;
wire n_126;
wire n_118;
wire n_32;
wire n_84;
wire n_131;
wire n_112;
wire n_55;
wire n_86;
wire n_75;
wire n_105;
wire n_72;
wire n_136;
wire n_43;
wire n_76;
wire n_89;
wire n_68;
wire n_27;
wire n_53;
wire n_67;
wire n_77;
wire n_20;
wire n_54;
wire n_123;
wire n_83;
wire n_28;
wire n_48;
wire n_100;
wire n_92;
wire n_25;
wire n_30;
wire n_59;
wire n_18;
wire n_110;
wire n_66;
wire n_134;
wire n_82;
wire n_106;
wire n_61;
wire n_21;
wire n_99;
wire n_109;
wire n_93;
wire n_132;
wire n_51;
wire n_140;
wire n_96;
wire n_39;
INVx2_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
INVx2_ASAP7_75t_SL g18 ( .A(n_2), .Y(n_18) );
BUFx3_ASAP7_75t_L g19 ( .A(n_5), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_9), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_10), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_8), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_15), .Y(n_23) );
BUFx2_ASAP7_75t_L g24 ( .A(n_11), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_2), .Y(n_25) );
BUFx2_ASAP7_75t_L g26 ( .A(n_4), .Y(n_26) );
BUFx5_ASAP7_75t_L g27 ( .A(n_14), .Y(n_27) );
BUFx6f_ASAP7_75t_L g28 ( .A(n_19), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_17), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_26), .B(n_24), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_27), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_27), .Y(n_32) );
INVx2_ASAP7_75t_L g33 ( .A(n_27), .Y(n_33) );
INVx2_ASAP7_75t_L g34 ( .A(n_27), .Y(n_34) );
INVx3_ASAP7_75t_L g35 ( .A(n_20), .Y(n_35) );
AND2x4_ASAP7_75t_L g36 ( .A(n_25), .B(n_0), .Y(n_36) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_18), .B(n_0), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_18), .B(n_1), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_31), .Y(n_39) );
AO22x2_ASAP7_75t_L g40 ( .A1(n_30), .A2(n_21), .B1(n_22), .B2(n_20), .Y(n_40) );
BUFx10_ASAP7_75t_L g41 ( .A(n_36), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_31), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_32), .Y(n_43) );
OA21x2_ASAP7_75t_L g44 ( .A1(n_29), .A2(n_22), .B(n_21), .Y(n_44) );
NAND2xp5_ASAP7_75t_L g45 ( .A(n_29), .B(n_16), .Y(n_45) );
AND2x4_ASAP7_75t_L g46 ( .A(n_36), .B(n_35), .Y(n_46) );
INVx2_ASAP7_75t_L g47 ( .A(n_32), .Y(n_47) );
INVx1_ASAP7_75t_L g48 ( .A(n_33), .Y(n_48) );
NAND2x1p5_ASAP7_75t_L g49 ( .A(n_36), .B(n_23), .Y(n_49) );
INVx2_ASAP7_75t_SL g50 ( .A(n_41), .Y(n_50) );
BUFx6f_ASAP7_75t_L g51 ( .A(n_41), .Y(n_51) );
BUFx4_ASAP7_75t_SL g52 ( .A(n_40), .Y(n_52) );
BUFx6f_ASAP7_75t_L g53 ( .A(n_41), .Y(n_53) );
INVx2_ASAP7_75t_L g54 ( .A(n_47), .Y(n_54) );
INVx8_ASAP7_75t_L g55 ( .A(n_46), .Y(n_55) );
NAND3xp33_ASAP7_75t_L g56 ( .A(n_44), .B(n_38), .C(n_37), .Y(n_56) );
NOR2xp67_ASAP7_75t_L g57 ( .A(n_45), .B(n_35), .Y(n_57) );
OAI21x1_ASAP7_75t_L g58 ( .A1(n_49), .A2(n_35), .B(n_34), .Y(n_58) );
INVx3_ASAP7_75t_L g59 ( .A(n_49), .Y(n_59) );
NAND3xp33_ASAP7_75t_L g60 ( .A(n_44), .B(n_35), .C(n_34), .Y(n_60) );
INVx1_ASAP7_75t_L g61 ( .A(n_44), .Y(n_61) );
INVx2_ASAP7_75t_L g62 ( .A(n_39), .Y(n_62) );
HB1xp67_ASAP7_75t_L g63 ( .A(n_52), .Y(n_63) );
BUFx6f_ASAP7_75t_L g64 ( .A(n_51), .Y(n_64) );
INVx2_ASAP7_75t_L g65 ( .A(n_62), .Y(n_65) );
AOI21xp5_ASAP7_75t_L g66 ( .A1(n_50), .A2(n_48), .B(n_42), .Y(n_66) );
INVx2_ASAP7_75t_L g67 ( .A(n_62), .Y(n_67) );
INVx2_ASAP7_75t_L g68 ( .A(n_62), .Y(n_68) );
NAND2xp5_ASAP7_75t_SL g69 ( .A(n_53), .B(n_43), .Y(n_69) );
BUFx6f_ASAP7_75t_L g70 ( .A(n_59), .Y(n_70) );
INVx5_ASAP7_75t_L g71 ( .A(n_55), .Y(n_71) );
INVx5_ASAP7_75t_L g72 ( .A(n_55), .Y(n_72) );
INVx4_ASAP7_75t_L g73 ( .A(n_55), .Y(n_73) );
AOI21xp5_ASAP7_75t_L g74 ( .A1(n_54), .A2(n_56), .B(n_61), .Y(n_74) );
INVx2_ASAP7_75t_L g75 ( .A(n_65), .Y(n_75) );
OR2x6_ASAP7_75t_L g76 ( .A(n_63), .B(n_58), .Y(n_76) );
OAI21xp5_ASAP7_75t_L g77 ( .A1(n_74), .A2(n_60), .B(n_57), .Y(n_77) );
BUFx6f_ASAP7_75t_L g78 ( .A(n_64), .Y(n_78) );
INVx3_ASAP7_75t_L g79 ( .A(n_71), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_65), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_67), .Y(n_81) );
BUFx4f_ASAP7_75t_SL g82 ( .A(n_73), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_72), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_68), .Y(n_84) );
OR2x6_ASAP7_75t_L g85 ( .A(n_70), .B(n_28), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_78), .Y(n_86) );
AO21x2_ASAP7_75t_L g87 ( .A1(n_77), .A2(n_69), .B(n_66), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_83), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_75), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_80), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_81), .Y(n_91) );
OR2x6_ASAP7_75t_L g92 ( .A(n_76), .B(n_3), .Y(n_92) );
INVx4_ASAP7_75t_L g93 ( .A(n_82), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_84), .Y(n_94) );
INVx3_ASAP7_75t_SL g95 ( .A(n_79), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_89), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_90), .Y(n_97) );
BUFx3_ASAP7_75t_L g98 ( .A(n_93), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_91), .Y(n_99) );
NAND2xp33_ASAP7_75t_R g100 ( .A(n_92), .B(n_85), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_94), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_86), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_86), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_86), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_88), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_86), .Y(n_106) );
INVx2_ASAP7_75t_SL g107 ( .A(n_95), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_100), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_96), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_97), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_99), .Y(n_111) );
AND2x4_ASAP7_75t_L g112 ( .A(n_102), .B(n_87), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_101), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_98), .Y(n_114) );
OR2x2_ASAP7_75t_L g115 ( .A(n_105), .B(n_12), .Y(n_115) );
AND2x4_ASAP7_75t_SL g116 ( .A(n_107), .B(n_13), .Y(n_116) );
AND2x2_ASAP7_75t_L g117 ( .A(n_103), .B(n_104), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_103), .B(n_104), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_106), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_108), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_109), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_112), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_117), .B(n_118), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_110), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_114), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_116), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_110), .B(n_113), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_111), .Y(n_128) );
NOR2xp67_ASAP7_75t_SL g129 ( .A(n_126), .B(n_115), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_125), .B(n_119), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_123), .Y(n_131) );
NAND2x1p5_ASAP7_75t_L g132 ( .A(n_129), .B(n_120), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_131), .B(n_122), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_132), .B(n_130), .Y(n_134) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_134), .B(n_133), .Y(n_135) );
INVx1_ASAP7_75t_SL g136 ( .A(n_135), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_136), .Y(n_137) );
BUFx2_ASAP7_75t_L g138 ( .A(n_137), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_138), .Y(n_139) );
INVx1_ASAP7_75t_SL g140 ( .A(n_139), .Y(n_140) );
AOI221xp5_ASAP7_75t_L g141 ( .A1(n_140), .A2(n_128), .B1(n_127), .B2(n_124), .C(n_121), .Y(n_141) );
endmodule