module fake_jpeg_1861_n_408 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_408);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_408;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_11),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_54),
.B(n_56),
.Y(n_136)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_55),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_10),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_57),
.B(n_59),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_20),
.B(n_10),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_62),
.B(n_69),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_23),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g130 ( 
.A(n_63),
.Y(n_130)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_66),
.Y(n_149)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_24),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_72),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_73),
.B(n_74),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_12),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_29),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_79),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_82),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_25),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_96),
.Y(n_143)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_86),
.Y(n_181)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_40),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_92),
.Y(n_142)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_20),
.B(n_12),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_33),
.Y(n_97)
);

BUFx16f_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_22),
.B(n_7),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_105),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_22),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_106),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_103),
.B(n_111),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_104),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_25),
.B(n_7),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_47),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_47),
.B(n_13),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_109),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_13),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_34),
.B1(n_44),
.B2(n_42),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_113),
.A2(n_122),
.B1(n_155),
.B2(n_161),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_114),
.B(n_115),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_52),
.B1(n_53),
.B2(n_34),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_116),
.A2(n_126),
.B1(n_129),
.B2(n_161),
.Y(n_201)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_60),
.A2(n_53),
.B1(n_41),
.B2(n_42),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_76),
.B1(n_80),
.B2(n_82),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_91),
.A2(n_28),
.B1(n_38),
.B2(n_36),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_127),
.A2(n_159),
.B1(n_155),
.B2(n_122),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_44),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_128),
.B(n_160),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_86),
.A2(n_41),
.B1(n_50),
.B2(n_28),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_141),
.B(n_152),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_79),
.B(n_50),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_89),
.A2(n_19),
.B1(n_38),
.B2(n_36),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_68),
.A2(n_26),
.B1(n_19),
.B2(n_49),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_26),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_63),
.A2(n_32),
.B1(n_4),
.B2(n_5),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_66),
.B(n_13),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_169),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_77),
.B(n_14),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_78),
.A2(n_32),
.B1(n_16),
.B2(n_5),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_170),
.A2(n_151),
.B1(n_163),
.B2(n_176),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_67),
.B(n_16),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_175),
.B(n_112),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_75),
.B(n_3),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_177),
.B(n_180),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_103),
.B(n_3),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_90),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_183),
.B(n_190),
.Y(n_252)
);

OR2x4_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_65),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_184),
.Y(n_258)
);

OR2x2_ASAP7_75t_SL g185 ( 
.A(n_137),
.B(n_71),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g279 ( 
.A(n_185),
.B(n_219),
.Y(n_279)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_186),
.Y(n_265)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_188),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_127),
.A2(n_95),
.B1(n_64),
.B2(n_61),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_3),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_191),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_70),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_193),
.B(n_199),
.Y(n_255)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_142),
.Y(n_195)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_196),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_135),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_202),
.Y(n_251)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_136),
.B(n_71),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_200),
.Y(n_282)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_206),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_177),
.A2(n_4),
.B(n_5),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_204),
.B(n_226),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_171),
.A2(n_4),
.B1(n_149),
.B2(n_179),
.Y(n_205)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_159),
.A2(n_4),
.B1(n_173),
.B2(n_178),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_207),
.A2(n_167),
.B1(n_158),
.B2(n_118),
.Y(n_244)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_210),
.B(n_214),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_147),
.B(n_113),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_211),
.B(n_215),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_139),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_212),
.B(n_229),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_145),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_120),
.B(n_125),
.Y(n_215)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_217),
.Y(n_261)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_154),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_218),
.A2(n_222),
.B1(n_228),
.B2(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_119),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_220),
.B(n_224),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_131),
.B(n_174),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_221),
.B(n_223),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_121),
.A2(n_176),
.B1(n_165),
.B2(n_132),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_138),
.B(n_168),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_121),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_138),
.A2(n_168),
.B1(n_139),
.B2(n_162),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_225),
.B(n_231),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_117),
.B(n_135),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_227),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_133),
.B(n_162),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_148),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_230),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_132),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_233),
.Y(n_270)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_148),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_117),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_237),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_156),
.A2(n_134),
.B(n_112),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_134),
.A2(n_181),
.B(n_153),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_184),
.B1(n_235),
.B2(n_193),
.Y(n_256)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_167),
.B(n_158),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g278 ( 
.A1(n_238),
.A2(n_240),
.A3(n_184),
.B1(n_149),
.B2(n_200),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_153),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_219),
.A2(n_158),
.B1(n_183),
.B2(n_211),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_218),
.A2(n_208),
.B1(n_239),
.B2(n_201),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_215),
.A2(n_229),
.B1(n_212),
.B2(n_221),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_212),
.A2(n_223),
.B1(n_238),
.B2(n_182),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_250),
.A2(n_260),
.B1(n_262),
.B2(n_264),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_213),
.A2(n_209),
.B1(n_185),
.B2(n_190),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_199),
.A2(n_236),
.B1(n_224),
.B2(n_216),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_186),
.A2(n_194),
.B1(n_226),
.B2(n_232),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_222),
.A2(n_217),
.B1(n_193),
.B2(n_210),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_267),
.A2(n_272),
.B1(n_282),
.B2(n_242),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_188),
.A2(n_204),
.B1(n_192),
.B2(n_240),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_269),
.A2(n_244),
.B1(n_267),
.B2(n_282),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_192),
.A2(n_218),
.B1(n_219),
.B2(n_201),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_276),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_240),
.B(n_262),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_284),
.A2(n_286),
.B(n_269),
.Y(n_323)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_285),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_253),
.B(n_279),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_258),
.A2(n_253),
.B1(n_246),
.B2(n_245),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_288),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_274),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_289),
.B(n_290),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_273),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_258),
.A2(n_250),
.B1(n_276),
.B2(n_247),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_292),
.A2(n_296),
.B(n_265),
.Y(n_330)
);

AOI221xp5_ASAP7_75t_L g337 ( 
.A1(n_293),
.A2(n_305),
.B1(n_286),
.B2(n_297),
.C(n_304),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_277),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_295),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_252),
.B(n_277),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_263),
.B(n_278),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_272),
.A2(n_248),
.B1(n_275),
.B2(n_279),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_297),
.A2(n_310),
.B1(n_312),
.B2(n_271),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_263),
.A2(n_283),
.B(n_259),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_298),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_280),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_301),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_255),
.B(n_283),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_304),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_274),
.B(n_241),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_255),
.B(n_260),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_306),
.C(n_313),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_261),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_248),
.B(n_251),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_242),
.B(n_243),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_309),
.Y(n_328)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_257),
.Y(n_309)
);

INVx13_ASAP7_75t_L g311 ( 
.A(n_249),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_254),
.C(n_243),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_281),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_265),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_316),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_SL g354 ( 
.A1(n_323),
.A2(n_316),
.B(n_311),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_287),
.A2(n_249),
.B1(n_271),
.B2(n_265),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_324),
.A2(n_310),
.B1(n_291),
.B2(n_314),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_308),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_336),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_330),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_333),
.A2(n_337),
.B1(n_311),
.B2(n_323),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_296),
.A2(n_305),
.B(n_284),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_334),
.A2(n_307),
.B(n_309),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_303),
.B(n_306),
.C(n_300),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_293),
.C(n_313),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_299),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_312),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_285),
.Y(n_351)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_328),
.Y(n_340)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_334),
.A2(n_293),
.B(n_288),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_341),
.A2(n_330),
.B(n_332),
.Y(n_360)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_342),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_335),
.B(n_321),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_347),
.C(n_349),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_338),
.A2(n_287),
.B1(n_302),
.B2(n_292),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_344),
.A2(n_346),
.B1(n_354),
.B2(n_355),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_294),
.Y(n_347)
);

XOR2x2_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_295),
.Y(n_348)
);

A2O1A1O1Ixp25_ASAP7_75t_L g357 ( 
.A1(n_348),
.A2(n_322),
.B(n_331),
.C(n_326),
.D(n_330),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_302),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_352),
.C(n_319),
.Y(n_365)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_351),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_315),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_353),
.A2(n_345),
.B(n_339),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_329),
.B(n_336),
.Y(n_356)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_356),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_357),
.B(n_358),
.Y(n_372)
);

NOR3xp33_ASAP7_75t_SL g358 ( 
.A(n_339),
.B(n_317),
.C(n_320),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_360),
.A2(n_361),
.B1(n_345),
.B2(n_342),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_353),
.Y(n_362)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_333),
.Y(n_380)
);

AOI322xp5_ASAP7_75t_L g366 ( 
.A1(n_341),
.A2(n_322),
.A3(n_337),
.B1(n_318),
.B2(n_332),
.C1(n_333),
.C2(n_329),
.Y(n_366)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_366),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_319),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_370),
.A2(n_344),
.B1(n_325),
.B2(n_324),
.Y(n_375)
);

AND2x6_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_348),
.Y(n_371)
);

AOI31xp67_ASAP7_75t_L g384 ( 
.A1(n_371),
.A2(n_367),
.A3(n_359),
.B(n_357),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_369),
.B(n_318),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_364),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_374),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_370),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_343),
.C(n_365),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_378),
.C(n_379),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_363),
.B(n_349),
.C(n_347),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_350),
.C(n_352),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_380),
.B(n_368),
.Y(n_387)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_382),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_386),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_SL g394 ( 
.A(n_384),
.B(n_387),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_372),
.A2(n_361),
.B(n_360),
.Y(n_386)
);

XOR2x1_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_368),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_362),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_385),
.B(n_378),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_392),
.B(n_396),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_324),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_376),
.C(n_385),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_377),
.C(n_346),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_385),
.B(n_381),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_395),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_397),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_399),
.B(n_400),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_371),
.C(n_325),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_401),
.B(n_390),
.C(n_394),
.Y(n_403)
);

NOR3xp33_ASAP7_75t_L g406 ( 
.A(n_403),
.B(n_398),
.C(n_327),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_404),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_405),
.B(n_406),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_402),
.Y(n_408)
);


endmodule