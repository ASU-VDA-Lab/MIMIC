module fake_jpeg_1543_n_164 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_0),
.B(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_30),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_35),
.Y(n_68)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_7),
.C(n_3),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_15),
.C(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_12),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g78 ( 
.A(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_4),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_46),
.Y(n_54)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_5),
.Y(n_48)
);

OR2x4_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_7),
.Y(n_49)
);

HAxp5_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_0),
.CON(n_55),
.SN(n_55)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_21),
.B1(n_27),
.B2(n_20),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_56),
.B1(n_60),
.B2(n_43),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_14),
.B1(n_13),
.B2(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_23),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_34),
.A2(n_23),
.B(n_11),
.C(n_12),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_8),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_10),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_36),
.A2(n_14),
.B(n_18),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_29),
.B(n_18),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_8),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_81),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_71),
.B1(n_73),
.B2(n_76),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_9),
.Y(n_81)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_10),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_71),
.B(n_66),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_14),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_87),
.B(n_94),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_10),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_99),
.Y(n_110)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_0),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_55),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_14),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_93),
.B(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_18),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_32),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_12),
.B1(n_40),
.B2(n_68),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_98),
.B1(n_77),
.B2(n_73),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_68),
.A2(n_70),
.B1(n_62),
.B2(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_101),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_77),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_71),
.B1(n_96),
.B2(n_52),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_85),
.C(n_87),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_97),
.C(n_86),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_112),
.B(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_74),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_74),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_123),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_107),
.A2(n_88),
.B1(n_82),
.B2(n_91),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_103),
.B1(n_102),
.B2(n_101),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_128),
.B(n_130),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_139),
.B1(n_130),
.B2(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_135),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_100),
.B1(n_114),
.B2(n_116),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_138),
.B1(n_127),
.B2(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_106),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_140),
.C(n_134),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_116),
.B1(n_109),
.B2(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_111),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_126),
.B1(n_120),
.B2(n_119),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_142),
.B1(n_146),
.B2(n_147),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_123),
.B(n_129),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_143),
.B(n_145),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_129),
.B1(n_127),
.B2(n_108),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_140),
.C(n_131),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_152),
.C(n_108),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_136),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_102),
.C(n_108),
.Y(n_154)
);

AOI321xp33_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_112),
.A3(n_142),
.B1(n_137),
.B2(n_131),
.C(n_147),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_150),
.A2(n_144),
.B1(n_135),
.B2(n_81),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_156),
.C(n_149),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_155),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_118),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_149),
.B(n_118),
.Y(n_157)
);

AOI21x1_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_158),
.B(n_67),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_53),
.A3(n_52),
.B1(n_66),
.B2(n_67),
.C1(n_104),
.C2(n_64),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_161),
.C(n_53),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_64),
.Y(n_164)
);


endmodule